magic
tech sky130A
magscale 1 2
timestamp 1702073639
<< pwell >>
rect -403 -1479 403 1479
<< nmos >>
rect -207 -1331 -147 1269
rect -89 -1331 -29 1269
rect 29 -1331 89 1269
rect 147 -1331 207 1269
<< ndiff >>
rect -265 1257 -207 1269
rect -265 -1319 -253 1257
rect -219 -1319 -207 1257
rect -265 -1331 -207 -1319
rect -147 1257 -89 1269
rect -147 -1319 -135 1257
rect -101 -1319 -89 1257
rect -147 -1331 -89 -1319
rect -29 1257 29 1269
rect -29 -1319 -17 1257
rect 17 -1319 29 1257
rect -29 -1331 29 -1319
rect 89 1257 147 1269
rect 89 -1319 101 1257
rect 135 -1319 147 1257
rect 89 -1331 147 -1319
rect 207 1257 265 1269
rect 207 -1319 219 1257
rect 253 -1319 265 1257
rect 207 -1331 265 -1319
<< ndiffc >>
rect -253 -1319 -219 1257
rect -135 -1319 -101 1257
rect -17 -1319 17 1257
rect 101 -1319 135 1257
rect 219 -1319 253 1257
<< psubdiff >>
rect -367 1409 367 1443
rect -367 -1409 -333 1409
rect 333 -1409 367 1409
rect -367 -1443 -271 -1409
rect 271 -1443 367 -1409
<< psubdiffcont >>
rect -271 -1443 271 -1409
<< poly >>
rect -210 1341 -144 1357
rect -210 1307 -194 1341
rect -160 1307 -144 1341
rect -210 1291 -144 1307
rect -92 1341 -26 1357
rect -92 1307 -76 1341
rect -42 1307 -26 1341
rect -92 1291 -26 1307
rect 26 1341 92 1357
rect 26 1307 42 1341
rect 76 1307 92 1341
rect 26 1291 92 1307
rect 144 1341 210 1357
rect 144 1307 160 1341
rect 194 1307 210 1341
rect 144 1291 210 1307
rect -207 1269 -147 1291
rect -89 1269 -29 1291
rect 29 1269 89 1291
rect 147 1269 207 1291
rect -207 -1357 -147 -1331
rect -89 -1357 -29 -1331
rect 29 -1357 89 -1331
rect 147 -1357 207 -1331
<< polycont >>
rect -194 1307 -160 1341
rect -76 1307 -42 1341
rect 42 1307 76 1341
rect 160 1307 194 1341
<< locali >>
rect -210 1307 -194 1341
rect -160 1307 -144 1341
rect -92 1307 -76 1341
rect -42 1307 -26 1341
rect 26 1307 42 1341
rect 76 1307 92 1341
rect 144 1307 160 1341
rect 194 1307 210 1341
rect -253 1257 -219 1273
rect -253 -1335 -219 -1319
rect -135 1257 -101 1273
rect -135 -1335 -101 -1319
rect -17 1257 17 1273
rect -17 -1335 17 -1319
rect 101 1257 135 1273
rect 101 -1335 135 -1319
rect 219 1257 253 1273
rect 219 -1335 253 -1319
rect -287 -1443 -271 -1409
rect 271 -1443 287 -1409
<< viali >>
rect -194 1307 -160 1341
rect -76 1307 -42 1341
rect 42 1307 76 1341
rect 160 1307 194 1341
rect -253 -1319 -219 1257
rect -135 -933 -101 871
rect -17 -1319 17 1257
rect 101 -933 135 871
rect 219 -1319 253 1257
<< metal1 >>
rect -206 1341 206 1347
rect -206 1307 -194 1341
rect -160 1307 -76 1341
rect -42 1307 42 1341
rect 76 1307 160 1341
rect 194 1307 206 1341
rect -206 1301 206 1307
rect -259 1257 -213 1269
rect -259 -1319 -253 1257
rect -219 1154 -213 1257
rect -23 1257 23 1269
rect -23 1154 -17 1257
rect -219 1118 -17 1154
rect -219 -1319 -213 1118
rect -141 871 -95 883
rect -141 -828 -135 871
rect -143 -834 -135 -828
rect -101 -828 -95 871
rect -101 -834 -91 -828
rect -143 -892 -135 -886
rect -141 -933 -135 -892
rect -101 -892 -91 -886
rect -101 -933 -95 -892
rect -141 -945 -95 -933
rect -259 -1331 -213 -1319
rect -23 -1319 -17 1118
rect 17 1154 23 1257
rect 213 1257 259 1269
rect 213 1154 219 1257
rect 17 1118 219 1154
rect 17 -1319 23 1118
rect 95 871 141 883
rect 95 -829 101 871
rect 91 -835 101 -829
rect 135 -829 141 871
rect 135 -835 143 -829
rect 91 -893 101 -887
rect 95 -933 101 -893
rect 135 -893 143 -887
rect 135 -933 141 -893
rect 95 -945 141 -933
rect -23 -1331 23 -1319
rect 213 -1319 219 1118
rect 253 -1319 259 1257
rect 213 -1331 259 -1319
<< via1 >>
rect -143 -886 -135 -834
rect -135 -886 -101 -834
rect -101 -886 -91 -834
rect 91 -887 101 -835
rect 101 -887 135 -835
rect 135 -887 143 -835
<< metal2 >>
rect -149 -886 -143 -834
rect -91 -846 -85 -834
rect 85 -846 91 -835
rect -91 -876 91 -846
rect -91 -886 -85 -876
rect 85 -887 91 -876
rect 143 -887 149 -835
<< labels >>
rlabel metal1 -160 1301 -76 1347 1 G
rlabel metal1 -219 1118 -17 1154 1 D
rlabel metal2 -91 -876 91 -846 1 S
rlabel psubdiffcont 1 -1426 1 -1426 1 B
rlabel psubdiffcont -271 -1443 271 -1409 1 B
<< properties >>
string FIXED_BBOX -350 -1426 350 1426
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 13 l 0.3 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 70 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

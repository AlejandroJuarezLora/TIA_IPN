* SPICE3 file created from opamp_flatten.ext - technology: sky130A

.subckt opamp_flatten vdd iref vin_n vin_p vout vss
X0 vss.t267 voe1.t236 vout.t101 vss.t145 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X1 vout.t117 voe1.t237 vss.t266 vss.t206 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X2 w_4660_n6791.t388 vin_n.t0 vbn.t120 w_4660_n6791.t148 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X3 voe1.t232 vin_p.t0 w_4660_n6791.t476 w_4660_n6791.t41 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X4 w_4660_n6791.t387 vin_n.t1 vbn.t119 w_4660_n6791.t37 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X5 w_4660_n6791.t386 vin_n.t2 vbn.t217 w_4660_n6791.t64 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X6 vout.t148 voe1.t238 vss.t265 vss.t203 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X7 w_4660_n6791.t385 vin_n.t3 vbn.t216 w_4660_n6791.t37 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X8 vdd.t314 iref.t30 vout.t52 vdd.t239 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X9 vss.t264 voe1.t239 vout.t159 vss.t139 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X10 vout.t158 voe1.t240 vss.t263 vss.t200 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X11 vbn.t215 vin_n.t4 w_4660_n6791.t384 w_4660_n6791.t7 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X12 vout.t147 voe1.t241 vss.t262 vss.t135 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X13 vout.t72 voe1.t242 vss.t261 vss.t197 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X14 vout.t211 iref.t31 vdd.t313 vdd.t108 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X15 vbn.t253 vin_n.t5 w_4660_n6791.t383 w_4660_n6791.t7 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X16 w_4660_n6791.t404 vin_p.t1 voe1.t165 w_4660_n6791.t291 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X17 vout.t160 voe1.t243 vss.t260 vss.t194 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=1.305 ps=9.58 w=4.5 l=0.45
X18 w_4660_n6791.t406 vin_p.t2 voe1.t167 w_4660_n6791.t141 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X19 w_4660_n6791.t405 vin_p.t3 voe1.t166 w_4660_n6791.t291 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X20 w_4660_n6791.t454 vin_p.t4 voe1.t212 w_4660_n6791.t141 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X21 vdd.t312 iref.t32 vout.t265 vdd.t100 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X22 vbn.t252 vin_n.t6 w_4660_n6791.t382 w_4660_n6791.t86 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X23 voe1.t34 vin_p.t5 w_4660_n6791.t55 w_4660_n6791.t15 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X24 vout.t90 voe1.t244 vss.t259 vss.t127 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X25 vbn.t251 vin_n.t7 w_4660_n6791.t381 w_4660_n6791.t86 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X26 voe1.t8 vin_p.t6 w_4660_n6791.t16 w_4660_n6791.t15 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X27 vdd.t311 iref.t33 vout.t0 vdd.t237 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X28 vout.t236 iref.t34 vdd.t310 vdd.t96 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X29 vout.t293 iref.t35 vdd.t309 vdd.t235 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X30 voe1.t62 vin_p.t7 w_4660_n6791.t96 w_4660_n6791.t17 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X31 vdd.t289 iref.t36 w_4660_n6791.t56 vdd.t288 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X32 w_4660_n6791.t380 vin_n.t8 vbn.t123 w_4660_n6791.t39 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X33 vdd.t308 iref.t37 vout.t245 vdd.t232 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X34 voe1.t177 vin_p.t8 w_4660_n6791.t417 w_4660_n6791.t17 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X35 vdd.t307 iref.t38 vout.t11 vdd.t90 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X36 vout.t276 iref.t39 vdd.t306 vdd.t92 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X37 vbn.t122 vin_n.t9 w_4660_n6791.t379 w_4660_n6791.t25 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X38 w_4660_n6791.t411 vin_p.t9 voe1.t172 w_4660_n6791.t98 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X39 w_4660_n6791.t104 vin_p.t10 voe1.t67 w_4660_n6791.t64 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X40 w_4660_n6791.t378 vin_n.t10 vbn.t121 w_4660_n6791.t98 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X41 w_4660_n6791.t389 vin_p.t11 voe1.t150 w_4660_n6791.t64 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X42 voe1.t105 vbn.t260 vss.t280 vss.t269 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X43 w_4660_n6791.t391 vin_p.t12 voe1.t152 w_4660_n6791.t98 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X44 vdd.t305 iref.t40 vout.t212 vdd.t84 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X45 w_4660_n6791.t377 vin_n.t11 vbn.t174 w_4660_n6791.t60 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X46 vss.t258 voe1.t245 vout.t153 vss.t125 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X47 w_4660_n6791.t376 vin_n.t12 vbn.t173 w_4660_n6791.t64 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X48 vdd.t304 iref.t41 vout.t266 vdd.t230 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X49 vss.t277 vbn.t261 voe1.t101 vss.t275 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X50 vdd.t303 iref.t42 vout.t15 vdd.t78 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X51 vout.t278 iref.t43 vdd.t302 vdd.t80 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X52 vbn.t172 vin_n.t13 w_4660_n6791.t375 w_4660_n6791.t240 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X53 vss.t257 voe1.t246 vout.t154 vss.t123 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X54 voe1.t173 vin_p.t13 w_4660_n6791.t412 w_4660_n6791.t72 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X55 vbn.t238 vin_n.t14 w_4660_n6791.t374 w_4660_n6791.t23 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X56 vdd.t301 iref.t44 vout.t286 vdd.t228 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X57 vbn.t237 vin_n.t15 w_4660_n6791.t373 w_4660_n6791.t240 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X58 vss.t313 vbn.t262 voe1.t224 vss.t285 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X59 voe1.t168 vin_p.t14 w_4660_n6791.t407 w_4660_n6791.t72 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X60 voe1.t226 vbn.t263 vss.t315 vss.t278 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X61 vdd.t300 iref.t45 vout.t1 vdd.t72 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X62 vss.t256 voe1.t247 vout.t157 vss.t121 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X63 w_4660_n6791.t390 vin_p.t15 voe1.t151 w_4660_n6791.t92 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X64 w_4660_n6791.t186 vin_p.t16 voe1.t149 w_4660_n6791.t92 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X65 w_4660_n6791.t372 vin_n.t16 vbn.t236 w_4660_n6791.t141 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X66 vbn.t112 vin_n.t17 w_4660_n6791.t371 w_4660_n6791.t168 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X67 vout.t237 iref.t46 vdd.t299 vdd.t66 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X68 vout.t277 iref.t47 vdd.t298 vdd.t225 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X69 vss.t255 voe1.t248 vout.t129 vss.t119 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X70 w_4660_n6791.t370 vin_n.t18 vbn.t111 w_4660_n6791.t141 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X71 vbn.t110 vin_n.t19 w_4660_n6791.t369 w_4660_n6791.t168 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X72 vout.t116 voe1.t249 vss.t254 vss.t190 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X73 voe1.t135 vbn.t264 vss.t290 vss.t27 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X74 w_4660_n6791.t368 vin_n.t20 vbn.t157 w_4660_n6791.t166 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X75 vout.t115 voe1.t250 vss.t253 vss.t188 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X76 w_4660_n6791.t367 vin_n.t21 vbn.t156 w_4660_n6791.t112 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X77 vout.t118 voe1.t251 vss.t252 vss.t186 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X78 w_4660_n6791.t448 vin_p.t17 voe1.t207 w_4660_n6791.t35 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X79 vbn.t155 vin_n.t22 w_4660_n6791.t366 w_4660_n6791.t168 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X80 vdd.t297 iref.t48 vout.t267 vdd.t221 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X81 w_4660_n6791.t365 vin_n.t23 vbn.t235 w_4660_n6791.t166 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X82 vdd.t296 iref.t49 vout.t16 vdd.t62 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X83 vout.t152 voe1.t252 vss.t251 vss.t184 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X84 voe1.t139 vbn.t265 vss.t294 vss.t19 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X85 w_4660_n6791.t36 vin_p.t18 voe1.t21 w_4660_n6791.t35 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X86 w_4660_n6791.t364 vin_n.t24 vbn.t234 w_4660_n6791.t144 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X87 vout.t279 iref.t50 vdd.t295 vdd.t218 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X88 vdd.t294 iref.t51 w_4660_n6791.t459 vdd.t293 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X89 vss.t250 voe1.t253 vout.t179 vss.t111 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X90 vout.t149 voe1.t254 vss.t249 vss.t182 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X91 vdd.t292 iref.t52 w_4660_n6791.t470 vdd.t291 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X92 vout.t2 iref.t53 vdd.t290 vdd.t215 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X93 w_4660_n6791.t363 vin_n.t25 vbn.t233 w_4660_n6791.t163 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X94 w_4660_n6791.t362 vin_n.t26 vbn.t194 w_4660_n6791.t112 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X95 vout.t69 voe1.t255 vss.t248 vss.t180 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X96 vbn.t59 vbn.t58 vss.t320 vss.t299 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X97 vout.t238 iref.t54 vdd.t287 vdd.t213 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X98 w_4660_n6791.t361 vin_n.t27 vbn.t193 w_4660_n6791.t112 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X99 vss.t247 voe1.t256 vout.t166 vss.t177 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X100 vss.t30 vbn.t266 voe1.t51 vss.t29 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X101 vbn.t192 vin_n.t28 w_4660_n6791.t360 w_4660_n6791.t25 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X102 iref.t9 iref.t8 vdd.t286 vdd.t285 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X103 vdd.t284 iref.t55 w_4660_n6791.t124 vdd.t283 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X104 w_4660_n6791.t58 iref.t56 vdd.t282 vdd.t281 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X105 voe1.t0 vin_p.t19 w_4660_n6791.t1 w_4660_n6791.t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X106 voe1.t171 vin_p.t20 w_4660_n6791.t410 w_4660_n6791.t109 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X107 vbn.t160 vin_n.t29 w_4660_n6791.t359 w_4660_n6791.t25 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X108 vss.t272 vbn.t267 voe1.t85 vss.t271 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X109 voe1.t169 vin_p.t21 w_4660_n6791.t408 w_4660_n6791.t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X110 voe1.t72 vin_p.t22 w_4660_n6791.t111 w_4660_n6791.t109 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X111 vdd.t279 iref.t6 iref.t7 vdd.t278 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X112 vout.t230 iref.t57 vdd.t280 vdd.t207 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X113 w_4660_n6791.t358 vin_n.t30 vbn.t159 w_4660_n6791.t30 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X114 vbn.t158 vin_n.t31 w_4660_n6791.t357 w_4660_n6791.t11 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X115 vss.t36 vbn.t56 vbn.t57 vss.t23 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X116 voe1.t2 vin_p.t23 w_4660_n6791.t4 w_4660_n6791.t2 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X117 vout.t226 iref.t58 vdd.t277 vdd.t205 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X118 vbn.t88 vin_n.t32 w_4660_n6791.t356 w_4660_n6791.t11 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X119 voe1.t1 vin_p.t24 w_4660_n6791.t3 w_4660_n6791.t2 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X120 voe1.t225 vbn.t268 vss.t314 vss.t291 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X121 w_4660_n6791.t355 vin_n.t33 vbn.t87 w_4660_n6791.t70 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X122 iref.t29 iref.t28 vdd.t182 vdd.t181 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X123 w_4660_n6791.t354 vin_n.t34 vbn.t86 w_4660_n6791.t88 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X124 vdd.t276 iref.t59 vout.t17 vdd.t201 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X125 vbn.t133 vin_n.t35 w_4660_n6791.t353 w_4660_n6791.t5 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X126 vbn.t132 vin_n.t36 w_4660_n6791.t352 w_4660_n6791.t17 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X127 w_4660_n6791.t351 vin_n.t37 vbn.t131 w_4660_n6791.t144 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X128 w_4660_n6791.t350 vin_n.t38 vbn.t250 w_4660_n6791.t163 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X129 vbn.t55 vbn.t54 vss.t9 vss.t8 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X130 w_4660_n6791.t34 vin_p.t25 voe1.t20 w_4660_n6791.t33 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X131 w_4660_n6791.t349 vin_n.t39 vbn.t249 w_4660_n6791.t122 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X132 w_4660_n6791.t348 vin_n.t40 vbn.t248 w_4660_n6791.t163 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X133 w_4660_n6791.t423 vin_p.t26 voe1.t183 w_4660_n6791.t33 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X134 vout.t292 iref.t60 vdd.t275 vdd.t187 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X135 vdd.t274 iref.t61 vout.t45 vdd.t54 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X136 vout.t300 a_10611_n7515.t11 sky130_fd_pr__cap_mim_m3_1 l=15 w=17.55
X137 w_4660_n6791.t38 vin_p.t27 voe1.t22 w_4660_n6791.t37 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X138 vss.t246 voe1.t257 vout.t199 vss.t105 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X139 w_4660_n6791.t59 vin_p.t28 voe1.t35 w_4660_n6791.t37 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X140 w_4660_n6791.t347 vin_n.t41 vbn.t214 w_4660_n6791.t50 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X141 vbn.t213 vin_n.t42 w_4660_n6791.t346 w_4660_n6791.t77 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X142 voe1.t3 vin_p.t29 w_4660_n6791.t6 w_4660_n6791.t5 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X143 voe1.t4 vin_p.t30 w_4660_n6791.t8 w_4660_n6791.t7 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X144 vout.t34 iref.t62 vdd.t273 vdd.t179 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X145 vout.t301 a_10611_n7515.t10 sky130_fd_pr__cap_mim_m3_1 l=15 w=17.55
X146 w_4660_n6791.t345 vin_n.t43 vbn.t212 w_4660_n6791.t60 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X147 vout.t111 voe1.t258 vss.t245 vss.t101 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X148 voe1.t5 vin_p.t31 w_4660_n6791.t9 w_4660_n6791.t5 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X149 voe1.t19 vin_p.t32 w_4660_n6791.t32 w_4660_n6791.t7 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X150 vout.t18 iref.t63 vdd.t272 vdd.t177 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X151 vout.t283 iref.t64 vdd.t271 vdd.t175 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X152 vss.t244 voe1.t259 vout.t94 vss.t99 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X153 vout.t95 voe1.t260 vss.t243 vss.t97 sky130_fd_pr__nfet_01v8 ad=1.305 pd=9.58 as=0.6525 ps=4.79 w=4.5 l=0.45
X154 vout.t79 voe1.t261 vss.t242 vss.t172 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X155 voe1.t79 vin_p.t33 w_4660_n6791.t117 w_4660_n6791.t86 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X156 voe1.t185 vin_p.t34 w_4660_n6791.t425 w_4660_n6791.t77 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X157 vdd.t270 iref.t65 w_4660_n6791.t440 vdd.t269 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X158 vout.t43 iref.t66 vdd.t268 vdd.t44 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X159 voe1.t203 vin_p.t35 w_4660_n6791.t444 w_4660_n6791.t86 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X160 vout.t186 voe1.t262 vss.t241 vss.t95 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X161 vss.t240 voe1.t263 vout.t146 vss.t169 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X162 vout.t151 voe1.t264 vss.t239 vss.t93 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X163 voe1.t193 vin_p.t36 w_4660_n6791.t434 w_4660_n6791.t77 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X164 vout.t207 voe1.t265 vss.t238 vss.t167 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X165 w_4660_n6791.t146 iref.t67 vdd.t186 vdd.t185 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X166 vout.t53 iref.t68 vdd.t267 vdd.t172 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X167 vout.t200 voe1.t266 vss.t237 vss.t91 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X168 vout.t121 voe1.t267 vss.t236 vss.t87 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X169 voe1.t59 vbn.t269 vss.t35 vss.t31 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X170 vdd.t266 iref.t69 vout.t221 vdd.t38 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X171 vbn.t118 vin_n.t44 w_4660_n6791.t344 w_4660_n6791.t13 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X172 vout.t184 voe1.t268 vss.t235 vss.t165 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X173 vss.t234 voe1.t269 vout.t156 vss.t163 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X174 vbn.t117 vin_n.t45 w_4660_n6791.t343 w_4660_n6791.t13 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X175 vss.t233 voe1.t270 vout.t71 vss.t161 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X176 vss.t232 voe1.t271 vout.t192 vss.t159 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X177 w_4660_n6791.t435 vin_p.t37 voe1.t194 w_4660_n6791.t148 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X178 w_4660_n6791.t342 vin_n.t46 vbn.t116 w_4660_n6791.t70 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X179 vss.t231 voe1.t272 vout.t102 vss.t157 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X180 w_4660_n6791.t436 vin_p.t38 voe1.t195 w_4660_n6791.t148 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X181 vbn.t115 vin_n.t47 w_4660_n6791.t341 w_4660_n6791.t45 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X182 vss.t230 voe1.t273 vout.t198 vss.t155 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X183 vout.t297 iref.t70 vdd.t265 vdd.t167 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X184 vbn.t114 vin_n.t48 w_4660_n6791.t340 w_4660_n6791.t15 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X185 vdd.t264 iref.t71 vout.t255 vdd.t30 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X186 w_4660_n6791.t339 vin_n.t49 vbn.t113 w_4660_n6791.t130 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X187 vbn.t151 vin_n.t50 w_4660_n6791.t338 w_4660_n6791.t13 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X188 w_4660_n6791.t337 vin_n.t51 vbn.t150 w_4660_n6791.t130 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X189 voe1.t182 vin_p.t39 w_4660_n6791.t422 w_4660_n6791.t240 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X190 vout.t36 iref.t72 vdd.t263 vdd.t162 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X191 vdd.t262 iref.t73 vout.t54 vdd.t26 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X192 vss.t18 vbn.t52 vbn.t53 vss.t17 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X193 voe1.t196 vin_p.t40 w_4660_n6791.t437 w_4660_n6791.t240 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X194 vdd.t261 iref.t74 vout.t222 vdd.t24 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X195 w_4660_n6791.t336 vin_n.t52 vbn.t149 w_4660_n6791.t39 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X196 vss.t281 vbn.t50 vbn.t51 vss.t10 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X197 voe1.t128 vin_p.t41 w_4660_n6791.t169 w_4660_n6791.t168 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X198 vbn.t171 vin_n.t53 w_4660_n6791.t335 w_4660_n6791.t45 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X199 voe1.t189 vin_p.t42 w_4660_n6791.t429 w_4660_n6791.t118 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X200 vbn.t170 vin_n.t54 w_4660_n6791.t334 w_4660_n6791.t15 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X201 voe1.t205 vin_p.t43 w_4660_n6791.t446 w_4660_n6791.t168 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X202 vbn.t169 vin_n.t55 w_4660_n6791.t333 w_4660_n6791.t45 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X203 voe1.t80 vin_p.t44 w_4660_n6791.t119 w_4660_n6791.t118 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X204 w_4660_n6791.t167 vin_p.t45 voe1.t127 w_4660_n6791.t166 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X205 vout.t57 iref.t75 vdd.t260 vdd.t158 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X206 vdd.t259 iref.t76 vout.t30 vdd.t16 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X207 vbn.t49 vbn.t48 vss.t303 vss.t302 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X208 w_4660_n6791.t424 vin_p.t46 voe1.t184 w_4660_n6791.t166 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X209 vout.t284 iref.t77 vdd.t258 vdd.t155 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X210 voe1.t204 vin_p.t47 w_4660_n6791.t445 w_4660_n6791.t47 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X211 vbn.t247 vin_n.t56 w_4660_n6791.t332 w_4660_n6791.t41 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X212 w_4660_n6791.t331 vin_n.t57 vbn.t246 w_4660_n6791.t35 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X213 vbn.t47 vbn.t46 vss.t282 vss.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X214 vout.t51 iref.t78 vdd.t257 vdd.t153 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X215 voe1.t81 vin_p.t48 w_4660_n6791.t120 w_4660_n6791.t47 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X216 vout.t66 voe1.t274 vss.t229 vss.t81 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X217 vbn.t245 vin_n.t58 w_4660_n6791.t330 w_4660_n6791.t168 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X218 vout.t285 iref.t79 vdd.t256 vdd.t12 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X219 w_4660_n6791.t157 vin_p.t49 voe1.t119 w_4660_n6791.t112 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X220 w_4660_n6791.t433 iref.t80 vdd.t255 vdd.t254 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X221 w_4660_n6791.t329 vin_n.t59 vbn.t211 w_4660_n6791.t39 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X222 vss.t274 vbn.t44 vbn.t45 vss.t273 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X223 w_4660_n6791.t432 vin_p.t50 voe1.t192 w_4660_n6791.t144 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X224 w_4660_n6791.t89 vin_p.t51 voe1.t54 w_4660_n6791.t88 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X225 w_4660_n6791.t170 vin_p.t52 voe1.t129 w_4660_n6791.t112 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X226 vss.t228 voe1.t275 vout.t67 vss.t150 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X227 vout.t80 voe1.t276 vss.t227 vss.t77 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X228 vbn.t210 vin_n.t60 w_4660_n6791.t328 w_4660_n6791.t118 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X229 w_4660_n6791.t327 vin_n.t61 vbn.t209 w_4660_n6791.t39 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X230 w_4660_n6791.t155 vin_p.t53 voe1.t117 w_4660_n6791.t144 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X231 w_4660_n6791.t156 vin_p.t54 voe1.t118 w_4660_n6791.t88 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X232 voe1.t14 vin_p.t55 w_4660_n6791.t26 w_4660_n6791.t25 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X233 vss.t226 voe1.t277 vout.t204 vss.t75 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X234 vout.t123 voe1.t278 vss.t225 vss.t73 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X235 voe1.t15 vin_p.t56 w_4660_n6791.t27 w_4660_n6791.t25 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X236 vout.t59 voe1.t279 vss.t224 vss.t69 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X237 vdd.t253 iref.t14 iref.t15 vdd.t252 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X238 vout.t12 iref.t81 vdd.t251 vdd.t149 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X239 w_4660_n6791.t431 vin_p.t57 voe1.t191 w_4660_n6791.t70 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X240 w_4660_n6791.t165 vin_p.t58 voe1.t126 w_4660_n6791.t50 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X241 vout.t60 voe1.t280 vss.t223 vss.t67 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X242 vss.t222 voe1.t281 vout.t61 vss.t147 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X243 vss.t37 vbn.t42 vbn.t43 vss.t14 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X244 vout.t213 iref.t82 vdd.t250 vdd.t146 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X245 vss.t221 voe1.t282 vout.t181 vss.t143 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X246 vout.t180 voe1.t283 vss.t220 vss.t65 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X247 w_4660_n6791.t127 vin_p.t59 voe1.t87 w_4660_n6791.t70 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X248 w_4660_n6791.t90 vin_p.t60 voe1.t55 w_4660_n6791.t50 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X249 iref.t19 iref.t18 vdd.t249 vdd.t248 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X250 vbn.t256 vin_n.t62 w_4660_n6791.t326 w_4660_n6791.t17 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X251 vout.t178 voe1.t284 vss.t219 vss.t63 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X252 voe1.t56 vin_p.t61 w_4660_n6791.t91 w_4660_n6791.t67 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X253 voe1.t52 vin_p.t62 w_4660_n6791.t85 w_4660_n6791.t11 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X254 vdd.t247 iref.t83 w_4660_n6791.t472 vdd.t246 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X255 vout.t183 voe1.t285 vss.t218 vss.t61 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X256 vbn.t255 vin_n.t63 w_4660_n6791.t325 w_4660_n6791.t67 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X257 voe1.t120 vin_p.t63 w_4660_n6791.t158 w_4660_n6791.t11 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X258 vss.t217 voe1.t286 vout.t70 vss.t141 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X259 vdd.t245 iref.t84 vout.t231 vdd.t141 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X260 w_4660_n6791.t324 vin_n.t64 vbn.t254 w_4660_n6791.t94 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X261 voe1.t190 vin_p.t64 w_4660_n6791.t430 w_4660_n6791.t67 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X262 vout.t62 voe1.t287 vss.t216 vss.t59 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X263 vss.t215 voe1.t288 vout.t100 vss.t137 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X264 w_4660_n6791.t323 vin_n.t65 vbn.t65 w_4660_n6791.t94 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X265 w_4660_n6791.t19 iref.t85 vdd.t224 vdd.t223 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X266 a_10611_n7515.t5 vdd.t315 voe1.t77 vss.t41 sky130_fd_pr__nfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=0.15
X267 vss.t214 voe1.t289 vout.t91 vss.t133 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X268 vdd.t244 iref.t86 vout.t254 vdd.t6 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X269 vbn.t64 vin_n.t66 w_4660_n6791.t322 w_4660_n6791.t47 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X270 vss.t213 voe1.t290 vout.t150 vss.t131 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X271 vdd.t243 iref.t87 vout.t294 vdd.t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X272 iref.t13 iref.t12 vdd.t242 vdd.t241 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X273 vss.t212 voe1.t291 vout.t196 vss.t129 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X274 w_4660_n6791.t164 vin_p.t65 voe1.t125 w_4660_n6791.t163 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X275 vbn.t63 vin_n.t67 w_4660_n6791.t321 w_4660_n6791.t7 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X276 w_4660_n6791.t178 vin_p.t66 voe1.t142 w_4660_n6791.t163 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X277 vbn.t62 vin_n.t68 w_4660_n6791.t320 w_4660_n6791.t107 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X278 vbn.t61 vin_n.t69 w_4660_n6791.t319 w_4660_n6791.t107 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X279 vdd.t240 iref.t88 vout.t39 vdd.t239 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X280 w_4660_n6791.t136 vin_p.t67 voe1.t94 w_4660_n6791.t122 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X281 w_4660_n6791.t159 vin_p.t68 voe1.t121 w_4660_n6791.t122 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X282 w_4660_n6791.t318 vin_n.t70 vbn.t60 w_4660_n6791.t60 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X283 w_4660_n6791.t160 vin_p.t69 voe1.t122 w_4660_n6791.t79 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X284 w_4660_n6791.t317 vin_n.t71 vbn.t106 w_4660_n6791.t60 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X285 w_4660_n6791.t161 vin_p.t70 voe1.t123 w_4660_n6791.t79 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X286 vdd.t238 iref.t89 vout.t256 vdd.t237 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X287 vout.t19 iref.t90 vdd.t236 vdd.t235 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X288 vbn.t105 vin_n.t72 w_4660_n6791.t316 w_4660_n6791.t107 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X289 vout.t223 iref.t91 vdd.t234 vdd.t120 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X290 vdd.t233 iref.t92 vout.t268 vdd.t232 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X291 vout.t195 voe1.t292 vss.t211 vss.t53 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X292 vss.t312 vbn.t270 voe1.t223 vss.t287 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X293 voe1.t124 vin_p.t71 w_4660_n6791.t162 w_4660_n6791.t83 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X294 voe1.t102 vin_p.t72 w_4660_n6791.t143 w_4660_n6791.t23 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X295 voe1.t97 vin_p.t73 w_4660_n6791.t139 w_4660_n6791.t13 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X296 vout.t99 voe1.t293 vss.t210 vss.t49 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X297 vbn.t41 vbn.t40 vss.t319 vss.t39 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X298 vbn.t104 vin_n.t73 w_4660_n6791.t315 w_4660_n6791.t25 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X299 voe1.t228 vin_p.t74 w_4660_n6791.t471 w_4660_n6791.t13 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X300 vss.t276 vbn.t271 voe1.t100 vss.t275 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X301 voe1.t98 vin_p.t75 w_4660_n6791.t140 w_4660_n6791.t83 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X302 voe1.t140 vin_p.t76 w_4660_n6791.t176 w_4660_n6791.t23 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X303 vout.t145 voe1.t294 vss.t209 vss.t45 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X304 vout.t143 voe1.t295 vss.t208 vss.t43 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X305 vbn.t259 vin_n.t74 w_4660_n6791.t314 w_4660_n6791.t86 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X306 vout.t76 voe1.t296 vss.t207 vss.t206 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X307 vss.t205 voe1.t297 vout.t163 vss.t117 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X308 voe1.t104 vbn.t272 vss.t279 vss.t278 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X309 vdd.t231 iref.t93 vout.t3 vdd.t230 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X310 vout.t122 voe1.t298 vss.t204 vss.t203 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X311 vss.t202 voe1.t299 vout.t164 vss.t115 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X312 voe1.t230 vbn.t273 vss.t318 vss.t309 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X313 vdd.t229 iref.t94 vout.t239 vdd.t228 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X314 w_4660_n6791.t137 vin_p.t77 voe1.t95 w_4660_n6791.t52 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X315 w_4660_n6791.t177 vin_p.t78 voe1.t141 w_4660_n6791.t130 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X316 vout.t44 iref.t95 vdd.t227 vdd.t118 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X317 vout.t110 voe1.t300 vss.t201 vss.t200 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X318 vss.t199 voe1.t301 vout.t97 vss.t113 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X319 w_4660_n6791.t138 vin_p.t79 voe1.t96 w_4660_n6791.t130 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X320 voe1.t48 vbn.t274 vss.t28 vss.t27 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X321 w_4660_n6791.t74 vin_p.t80 voe1.t43 w_4660_n6791.t52 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X322 w_4660_n6791.t313 vin_n.t75 vbn.t258 w_4660_n6791.t166 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X323 vout.t173 voe1.t302 vss.t198 vss.t197 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X324 vss.t196 voe1.t303 vout.t127 vss.t109 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X325 w_4660_n6791.t312 vin_n.t76 vbn.t257 w_4660_n6791.t130 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X326 w_4660_n6791.t311 vin_n.t77 vbn.t224 w_4660_n6791.t148 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X327 vout.t98 voe1.t304 vss.t195 vss.t194 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=1.305 ps=9.58 w=4.5 l=0.45
X328 vbn.t223 vin_n.t78 w_4660_n6791.t310 w_4660_n6791.t107 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X329 vout.t240 iref.t96 vdd.t226 vdd.t225 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X330 w_4660_n6791.t309 vin_n.t79 vbn.t222 w_4660_n6791.t102 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X331 vbn.t109 vin_n.t80 w_4660_n6791.t308 w_4660_n6791.t109 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X332 w_4660_n6791.t307 vin_n.t81 vbn.t108 w_4660_n6791.t102 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X333 vss.t6 vbn.t275 voe1.t11 vss.t5 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X334 vdd.t222 iref.t97 vout.t257 vdd.t221 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X335 vss.t193 voe1.t305 vout.t82 vss.t107 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X336 voe1.t24 vin_p.t81 w_4660_n6791.t42 w_4660_n6791.t41 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X337 voe1.t26 vin_p.t82 w_4660_n6791.t46 w_4660_n6791.t45 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X338 vout.t298 iref.t98 vdd.t220 vdd.t114 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X339 vout.t20 iref.t99 vdd.t219 vdd.t218 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X340 voe1.t145 vin_p.t83 w_4660_n6791.t181 w_4660_n6791.t45 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X341 vss.t293 vbn.t276 voe1.t138 vss.t29 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X342 voe1.t143 vin_p.t84 w_4660_n6791.t179 w_4660_n6791.t41 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X343 vout.t40 iref.t100 vdd.t217 vdd.t110 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X344 vout.t229 iref.t101 vdd.t216 vdd.t215 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X345 vout.t41 iref.t102 vdd.t214 vdd.t213 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X346 vbn.t107 vin_n.t82 w_4660_n6791.t306 w_4660_n6791.t62 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X347 vbn.t130 vin_n.t83 w_4660_n6791.t305 w_4660_n6791.t41 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X348 vbn.t129 vin_n.t84 w_4660_n6791.t304 w_4660_n6791.t62 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X349 voe1.t29 vbn.t277 vss.t22 vss.t21 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X350 vdd.t212 iref.t103 vout.t4 vdd.t106 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X351 w_4660_n6791.t142 vin_p.t85 voe1.t99 w_4660_n6791.t141 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X352 w_4660_n6791.t75 vin_p.t86 voe1.t44 w_4660_n6791.t39 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X353 vout.t55 iref.t104 vdd.t211 vdd.t104 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X354 w_4660_n6791.t40 vin_p.t87 voe1.t23 w_4660_n6791.t39 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X355 a_10611_n7515.t4 vdd.t316 voe1.t12 vss.t7 sky130_fd_pr__nfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=0.15
X356 voe1.t137 vbn.t278 vss.t292 vss.t291 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X357 w_4660_n6791.t441 vin_p.t88 voe1.t200 w_4660_n6791.t141 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X358 w_4660_n6791.t303 vin_n.t85 vbn.t128 w_4660_n6791.t52 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X359 vbn.t191 vin_n.t86 w_4660_n6791.t302 w_4660_n6791.t43 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X360 vout.t252 iref.t105 vdd.t210 vdd.t102 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X361 vdd.t209 iref.t106 vout.t227 vdd.t98 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X362 vout.t42 iref.t107 vdd.t208 vdd.t207 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X363 vbn.t190 vin_n.t87 w_4660_n6791.t301 w_4660_n6791.t43 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X364 w_4660_n6791.t300 vin_n.t88 vbn.t189 w_4660_n6791.t30 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X365 vout.t214 iref.t108 vdd.t206 vdd.t205 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X366 w_4660_n6791.t299 vin_n.t89 vbn.t205 w_4660_n6791.t30 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X367 w_4660_n6791.t452 iref.t109 vdd.t204 vdd.t203 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X368 vbn.t204 vin_n.t90 w_4660_n6791.t298 w_4660_n6791.t11 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X369 w_4660_n6791.t297 vin_n.t91 vbn.t203 w_4660_n6791.t30 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X370 vdd.t202 iref.t110 vout.t21 vdd.t201 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X371 vdd.t200 iref.t111 vout.t258 vdd.t94 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X372 vout.t302 a_10611_n7515.t9 sky130_fd_pr__cap_mim_m3_1 l=15 w=17.55
X373 w_4660_n6791.t457 iref.t112 vdd.t199 vdd.t198 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X374 vss.t192 voe1.t306 vout.t203 vss.t103 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X375 w_4660_n6791.t95 vin_p.t89 voe1.t61 w_4660_n6791.t94 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X376 vdd.t197 iref.t113 w_4660_n6791.t69 vdd.t196 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X377 w_4660_n6791.t65 vin_p.t90 voe1.t38 w_4660_n6791.t64 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X378 w_4660_n6791.t419 vin_p.t91 voe1.t179 w_4660_n6791.t94 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X379 w_4660_n6791.t296 vin_n.t92 vbn.t208 w_4660_n6791.t291 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X380 vout.t56 iref.t114 vdd.t195 vdd.t88 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X381 w_4660_n6791.t76 vin_p.t92 voe1.t45 w_4660_n6791.t64 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X382 vout.t132 voe1.t307 vss.t191 vss.t190 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X383 iref.t5 iref.t4 vdd.t194 vdd.t193 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X384 vdd.t192 iref.t115 w_4660_n6791.t467 vdd.t191 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X385 vdd.t190 iref.t116 vout.t31 vdd.t86 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X386 vout.t193 voe1.t308 vss.t189 vss.t188 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X387 vbn.t207 vin_n.t93 w_4660_n6791.t295 w_4660_n6791.t62 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X388 vout.t109 voe1.t309 vss.t187 vss.t186 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X389 vdd.t189 iref.t117 vout.t46 vdd.t82 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X390 vout.t253 iref.t118 vdd.t188 vdd.t187 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X391 vout.t206 voe1.t310 vss.t185 vss.t184 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X392 w_4660_n6791.t460 iref.t119 vdd.t184 vdd.t183 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X393 voe1.t186 vin_p.t93 w_4660_n6791.t426 w_4660_n6791.t107 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X394 vout.t106 voe1.t311 vss.t183 vss.t182 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X395 voe1.t146 vin_p.t94 w_4660_n6791.t182 w_4660_n6791.t107 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X396 w_4660_n6791.t294 vin_n.t94 vbn.t206 w_4660_n6791.t291 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X397 vout.t114 voe1.t312 vss.t181 vss.t180 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X398 vss.t179 voe1.t313 vout.t93 vss.t89 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X399 w_4660_n6791.t293 vin_n.t95 vbn.t188 w_4660_n6791.t291 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X400 vout.t296 iref.t120 vdd.t180 vdd.t179 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X401 vss.t178 voe1.t314 vout.t85 vss.t177 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X402 w_4660_n6791.t93 vin_p.t95 voe1.t60 w_4660_n6791.t92 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X403 w_4660_n6791.t292 vin_n.t96 vbn.t187 w_4660_n6791.t291 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X404 vbn.t154 vin_n.t97 w_4660_n6791.t290 w_4660_n6791.t118 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X405 vout.t234 iref.t121 vdd.t178 vdd.t177 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X406 w_4660_n6791.t183 vin_p.t96 voe1.t147 w_4660_n6791.t92 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X407 vbn.t153 vin_n.t98 w_4660_n6791.t289 w_4660_n6791.t15 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X408 vout.t201 voe1.t315 vss.t176 vss.t85 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X409 vout.t246 iref.t122 vdd.t176 vdd.t175 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X410 vbn.t152 vin_n.t99 w_4660_n6791.t288 w_4660_n6791.t15 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X411 w_4660_n6791.t101 vin_p.t97 voe1.t65 w_4660_n6791.t60 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X412 w_4660_n6791.t401 vin_p.t98 voe1.t162 w_4660_n6791.t60 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X413 vout.t13 iref.t123 vdd.t174 vdd.t64 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X414 vbn.t148 vin_n.t100 w_4660_n6791.t287 w_4660_n6791.t17 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X415 vss.t34 vbn.t279 voe1.t58 vss.t33 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X416 vout.t215 iref.t124 vdd.t173 vdd.t172 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X417 vbn.t147 vin_n.t101 w_4660_n6791.t286 w_4660_n6791.t17 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X418 vdd.t171 iref.t125 vout.t295 vdd.t60 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X419 w_4660_n6791.t285 vin_n.t102 vbn.t146 w_4660_n6791.t98 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X420 vout.t142 voe1.t316 vss.t175 vss.t83 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X421 w_4660_n6791.t284 vin_n.t103 vbn.t100 w_4660_n6791.t98 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X422 w_4660_n6791.t283 vin_n.t104 vbn.t99 w_4660_n6791.t94 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X423 w_4660_n6791.t20 iref.t126 vdd.t170 vdd.t169 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X424 vbn.t98 vin_n.t105 w_4660_n6791.t282 w_4660_n6791.t43 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X425 vout.t241 iref.t127 vdd.t168 vdd.t167 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X426 vdd.t166 iref.t128 vout.t22 vdd.t58 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X427 vbn.t97 vin_n.t106 w_4660_n6791.t281 w_4660_n6791.t72 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X428 vss.t11 vbn.t38 vbn.t39 vss.t10 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X429 voe1.t49 vin_p.t99 w_4660_n6791.t81 w_4660_n6791.t2 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X430 vdd.t165 iref.t129 w_4660_n6791.t461 vdd.t164 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X431 w_4660_n6791.t280 vin_n.t107 vbn.t73 w_4660_n6791.t166 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X432 vbn.t37 vbn.t36 vss.t308 vss.t307 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X433 vbn.t72 vin_n.t108 w_4660_n6791.t279 w_4660_n6791.t72 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X434 voe1.t176 vin_p.t100 w_4660_n6791.t416 w_4660_n6791.t2 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X435 vout.t6 iref.t130 vdd.t163 vdd.t162 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X436 vss.t174 voe1.t317 vout.t139 vss.t79 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X437 vbn.t35 vbn.t34 vss.t298 vss.t296 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X438 vbn.t71 vin_n.t109 w_4660_n6791.t278 w_4660_n6791.t47 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X439 w_4660_n6791.t147 vin_p.t101 voe1.t106 w_4660_n6791.t102 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X440 iref.t21 iref.t20 vdd.t161 vdd.t160 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X441 w_4660_n6791.t277 vin_n.t110 vbn.t70 w_4660_n6791.t35 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X442 vbn.t33 vbn.t32 vss.t13 vss.t12 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X443 w_4660_n6791.t442 vin_p.t102 voe1.t201 w_4660_n6791.t33 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X444 vout.t188 voe1.t318 vss.t173 vss.t172 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X445 vss.t171 voe1.t319 vout.t197 vss.t71 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X446 vss.t1 vbn.t30 vbn.t31 vss.t0 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X447 vbn.t77 vin_n.t111 w_4660_n6791.t276 w_4660_n6791.t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X448 w_4660_n6791.t275 vin_n.t112 vbn.t76 w_4660_n6791.t35 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X449 w_4660_n6791.t103 vin_p.t103 voe1.t66 w_4660_n6791.t102 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X450 w_4660_n6791.t66 vin_p.t104 voe1.t39 w_4660_n6791.t33 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X451 vbn.t75 vin_n.t113 w_4660_n6791.t274 w_4660_n6791.t13 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X452 w_4660_n6791.t273 vin_n.t114 vbn.t74 w_4660_n6791.t122 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X453 vout.t242 iref.t131 vdd.t159 vdd.t158 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X454 vss.t170 voe1.t320 vout.t185 vss.t169 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X455 vss.t295 vbn.t28 vbn.t29 vss.t273 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X456 vbn.t242 vin_n.t115 w_4660_n6791.t272 w_4660_n6791.t83 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X457 vdd.t157 iref.t132 vout.t259 vdd.t56 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X458 vout.t269 iref.t133 vdd.t156 vdd.t155 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X459 vout.t126 voe1.t321 vss.t168 vss.t167 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X460 w_4660_n6791.t402 vin_p.t105 voe1.t163 w_4660_n6791.t37 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X461 vss.t3 vbn.t26 vbn.t27 vss.t2 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X462 vout.t5 iref.t134 vdd.t154 vdd.t153 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X463 vout.t81 voe1.t322 vss.t166 vss.t165 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X464 w_4660_n6791.t393 vin_p.t106 voe1.t154 w_4660_n6791.t37 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X465 vbn.t241 vin_n.t116 w_4660_n6791.t271 w_4660_n6791.t45 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X466 vss.t164 voe1.t323 vout.t167 vss.t163 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X467 voe1.t161 vin_p.t107 w_4660_n6791.t400 w_4660_n6791.t62 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X468 vbn.t240 vin_n.t117 w_4660_n6791.t270 w_4660_n6791.t109 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X469 vbn.t239 vin_n.t118 w_4660_n6791.t269 w_4660_n6791.t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X470 vss.t162 voe1.t324 vout.t64 vss.t161 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X471 vss.t15 vbn.t24 vbn.t25 vss.t14 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X472 voe1.t68 vin_p.t108 w_4660_n6791.t105 w_4660_n6791.t7 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X473 vout.t270 iref.t135 vdd.t152 vdd.t52 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X474 voe1.t37 vin_p.t109 w_4660_n6791.t63 w_4660_n6791.t62 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X475 vbn.t202 vin_n.t119 w_4660_n6791.t268 w_4660_n6791.t109 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X476 vbn.t201 vin_n.t120 w_4660_n6791.t267 w_4660_n6791.t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X477 vss.t160 voe1.t325 vout.t107 vss.t159 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X478 vout.t303 a_10611_n7515.t8 sky130_fd_pr__cap_mim_m3_1 l=15 w=17.55
X479 voe1.t178 vin_p.t110 w_4660_n6791.t418 w_4660_n6791.t7 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X480 vss.t158 voe1.t326 vout.t63 vss.t157 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X481 vdd.t151 iref.t136 vout.t23 vdd.t48 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X482 vout.t287 iref.t137 vdd.t150 vdd.t149 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X483 vout.t288 iref.t138 vdd.t148 vdd.t50 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X484 vss.t156 voe1.t327 vout.t155 vss.t155 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X485 vout.t177 voe1.t328 vss.t154 vss.t57 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X486 voe1.t208 vin_p.t111 w_4660_n6791.t449 w_4660_n6791.t86 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X487 voe1.t164 vin_p.t112 w_4660_n6791.t403 w_4660_n6791.t43 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X488 vbn.t23 vbn.t22 vss.t301 vss.t25 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X489 vout.t7 iref.t139 vdd.t147 vdd.t146 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X490 voe1.t155 vin_p.t113 w_4660_n6791.t394 w_4660_n6791.t43 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X491 voe1.t53 vin_p.t114 w_4660_n6791.t87 w_4660_n6791.t86 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X492 vdd.t145 iref.t140 vout.t243 vdd.t46 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X493 vbn.t200 vin_n.t121 w_4660_n6791.t266 w_4660_n6791.t109 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X494 vbn.t199 vin_n.t122 w_4660_n6791.t265 w_4660_n6791.t72 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X495 w_4660_n6791.t392 vin_p.t115 voe1.t153 w_4660_n6791.t30 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X496 vdd.t144 iref.t141 vout.t260 vdd.t40 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X497 vout.t216 iref.t142 vdd.t143 vdd.t42 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X498 vdd.t142 iref.t143 vout.t271 vdd.t141 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X499 w_4660_n6791.t399 vin_p.t116 voe1.t160 w_4660_n6791.t30 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X500 vbn.t186 vin_n.t123 w_4660_n6791.t264 w_4660_n6791.t23 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X501 vbn.t185 vin_n.t124 w_4660_n6791.t263 w_4660_n6791.t62 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X502 vout.t228 iref.t144 vdd.t140 vdd.t36 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X503 iref.t25 iref.t24 vdd.t139 vdd.t138 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X504 vdd.t137 iref.t145 w_4660_n6791.t97 vdd.t136 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X505 vdd.t135 iref.t146 vout.t24 vdd.t34 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X506 w_4660_n6791.t468 iref.t147 vdd.t134 vdd.t133 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X507 vbn.t184 vin_n.t125 w_4660_n6791.t262 w_4660_n6791.t83 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X508 vdd.t132 iref.t148 vout.t49 vdd.t32 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X509 vss.t153 voe1.t329 vout.t124 vss.t55 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X510 w_4660_n6791.t57 iref.t149 vdd.t131 vdd.t130 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X511 vdd.t125 iref.t150 w_4660_n6791.t125 vdd.t124 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X512 w_4660_n6791.t261 vin_n.t126 vbn.t183 w_4660_n6791.t88 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X513 vout.t251 iref.t151 vdd.t129 vdd.t28 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X514 voe1.t159 vin_p.t117 w_4660_n6791.t398 w_4660_n6791.t240 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X515 vbn.t198 vin_n.t127 w_4660_n6791.t260 w_4660_n6791.t5 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X516 vss.t152 voe1.t330 vout.t135 vss.t51 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X517 voe1.t158 vin_p.t118 w_4660_n6791.t397 w_4660_n6791.t240 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X518 vbn.t197 vin_n.t128 w_4660_n6791.t259 w_4660_n6791.t5 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X519 w_4660_n6791.t396 vin_p.t119 voe1.t157 w_4660_n6791.t291 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X520 vdd.t128 iref.t152 vout.t8 vdd.t22 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X521 vss.t151 voe1.t331 vout.t119 vss.t150 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X522 vbn.t196 vin_n.t129 w_4660_n6791.t258 w_4660_n6791.t43 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X523 a_10611_n7515.t3 vdd.t317 voe1.t78 vss.t42 sky130_fd_pr__nfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=0.15
X524 w_4660_n6791.t395 vin_p.t120 voe1.t156 w_4660_n6791.t291 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X525 vss.t149 voe1.t332 vout.t190 vss.t47 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X526 vdd.t127 iref.t22 iref.t23 vdd.t126 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X527 w_4660_n6791.t414 iref.t153 vdd.t123 vdd.t122 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X528 voe1.t175 vin_p.t121 w_4660_n6791.t415 w_4660_n6791.t168 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X529 voe1.t211 vin_p.t122 w_4660_n6791.t453 w_4660_n6791.t15 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X530 vbn.t195 vin_n.t130 w_4660_n6791.t257 w_4660_n6791.t77 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X531 vbn.t232 vin_n.t131 w_4660_n6791.t256 w_4660_n6791.t7 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X532 w_4660_n6791.t255 vin_n.t132 vbn.t231 w_4660_n6791.t33 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X533 voe1.t17 vin_p.t123 w_4660_n6791.t29 w_4660_n6791.t15 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X534 vss.t288 vbn.t280 voe1.t114 vss.t287 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X535 voe1.t202 vin_p.t124 w_4660_n6791.t443 w_4660_n6791.t168 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X536 vbn.t230 vin_n.t133 w_4660_n6791.t254 w_4660_n6791.t77 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X537 vss.t148 voe1.t333 vout.t75 vss.t147 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X538 vss.t146 voe1.t334 vout.t137 vss.t145 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X539 w_4660_n6791.t469 vin_p.t125 voe1.t227 w_4660_n6791.t166 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X540 vss.t144 voe1.t335 vout.t77 vss.t143 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X541 vbn.t21 vbn.t20 vss.t40 vss.t39 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X542 w_4660_n6791.t413 vin_p.t126 voe1.t174 w_4660_n6791.t166 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X543 vout.t48 iref.t154 vdd.t121 vdd.t120 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X544 vss.t142 voe1.t336 vout.t104 vss.t141 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X545 voe1.t9 vin_p.t127 w_4660_n6791.t18 w_4660_n6791.t17 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X546 vss.t140 voe1.t337 vout.t112 vss.t139 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X547 voe1.t76 vin_p.t128 w_4660_n6791.t116 w_4660_n6791.t17 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X548 vbn.t229 vin_n.t134 w_4660_n6791.t253 w_4660_n6791.t5 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X549 vss.t138 voe1.t338 vout.t130 vss.t137 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X550 vout.t168 voe1.t339 vss.t136 vss.t135 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X551 w_4660_n6791.t113 vin_p.t129 voe1.t73 w_4660_n6791.t112 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X552 w_4660_n6791.t99 vin_p.t130 voe1.t63 w_4660_n6791.t98 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X553 w_4660_n6791.t252 vin_n.t135 vbn.t137 w_4660_n6791.t148 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X554 w_4660_n6791.t172 vin_p.t131 voe1.t131 w_4660_n6791.t98 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X555 vss.t134 voe1.t340 vout.t141 vss.t133 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X556 voe1.t220 vbn.t281 vss.t310 vss.t309 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X557 w_4660_n6791.t451 vin_p.t132 voe1.t210 w_4660_n6791.t112 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X558 w_4660_n6791.t251 vin_n.t136 vbn.t136 w_4660_n6791.t148 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X559 voe1.t214 vin_p.t133 w_4660_n6791.t456 w_4660_n6791.t25 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X560 vss.t132 voe1.t341 vout.t140 vss.t131 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X561 voe1.t219 vin_p.t134 w_4660_n6791.t465 w_4660_n6791.t25 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X562 vss.t130 voe1.t342 vout.t182 vss.t129 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X563 vout.t78 voe1.t343 vss.t128 vss.t127 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X564 vbn.t135 vin_n.t137 w_4660_n6791.t250 w_4660_n6791.t86 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X565 w_4660_n6791.t249 vin_n.t138 vbn.t134 w_4660_n6791.t50 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X566 w_4660_n6791.t248 vin_n.t139 vbn.t92 w_4660_n6791.t92 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X567 vout.t261 iref.t155 vdd.t119 vdd.t118 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X568 voe1.t6 vin_p.t135 w_4660_n6791.t12 w_4660_n6791.t11 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X569 voe1.t42 vin_p.t136 w_4660_n6791.t73 w_4660_n6791.t72 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X570 voe1.t136 vin_p.t137 w_4660_n6791.t175 w_4660_n6791.t72 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X571 vss.t311 vbn.t282 voe1.t222 vss.t5 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X572 voe1.t30 vin_p.t138 w_4660_n6791.t49 w_4660_n6791.t11 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X573 w_4660_n6791.t184 iref.t156 vdd.t117 vdd.t116 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X574 vbn.t91 vin_n.t140 w_4660_n6791.t247 w_4660_n6791.t240 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X575 vbn.t90 vin_n.t141 w_4660_n6791.t246 w_4660_n6791.t118 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X576 w_4660_n6791.t245 vin_n.t142 vbn.t89 w_4660_n6791.t37 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X577 vbn.t81 vin_n.t143 w_4660_n6791.t244 w_4660_n6791.t118 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X578 vout.t299 iref.t157 vdd.t115 vdd.t114 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X579 vss.t126 voe1.t344 vout.t172 vss.t125 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X580 w_4660_n6791.t409 vin_p.t139 voe1.t170 w_4660_n6791.t163 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X581 w_4660_n6791.t150 vin_p.t140 voe1.t108 w_4660_n6791.t35 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X582 vdd.t113 iref.t0 iref.t1 vdd.t112 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X583 w_4660_n6791.t185 vin_p.t141 voe1.t148 w_4660_n6791.t35 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X584 voe1.t199 vbn.t283 vss.t305 vss.t21 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X585 w_4660_n6791.t174 vin_p.t142 voe1.t134 w_4660_n6791.t163 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X586 vout.t25 iref.t158 vdd.t111 vdd.t110 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X587 vbn.t80 vin_n.t144 w_4660_n6791.t243 w_4660_n6791.t47 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X588 vbn.t79 vin_n.t145 w_4660_n6791.t242 w_4660_n6791.t47 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X589 vss.t124 voe1.t345 vout.t165 vss.t123 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X590 vbn.t78 vin_n.t146 w_4660_n6791.t241 w_4660_n6791.t240 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X591 vbn.t103 vin_n.t147 w_4660_n6791.t239 w_4660_n6791.t77 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X592 w_4660_n6791.t238 vin_n.t148 vbn.t102 w_4660_n6791.t88 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X593 w_4660_n6791.t237 vin_n.t149 vbn.t101 w_4660_n6791.t144 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X594 w_4660_n6791.t236 vin_n.t150 vbn.t164 w_4660_n6791.t35 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X595 vout.t26 iref.t159 vdd.t109 vdd.t108 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X596 w_4660_n6791.t235 vin_n.t151 vbn.t163 w_4660_n6791.t88 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X597 vss.t122 voe1.t346 vout.t189 vss.t121 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X598 w_4660_n6791.t234 vin_n.t152 vbn.t162 w_4660_n6791.t94 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X599 vdd.t107 iref.t160 vout.t233 vdd.t106 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X600 w_4660_n6791.t233 vin_n.t153 vbn.t161 w_4660_n6791.t144 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X601 vout.t262 iref.t161 vdd.t105 vdd.t104 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X602 voe1.t86 vin_p.t143 w_4660_n6791.t126 w_4660_n6791.t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X603 voe1.t130 vin_p.t144 w_4660_n6791.t171 w_4660_n6791.t109 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X604 w_4660_n6791.t232 vin_n.t154 vbn.t127 w_4660_n6791.t79 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X605 voe1.t71 vin_p.t145 w_4660_n6791.t110 w_4660_n6791.t109 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X606 voe1.t115 vin_p.t146 w_4660_n6791.t153 w_4660_n6791.t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X607 vout.t224 iref.t162 vdd.t103 vdd.t102 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X608 w_4660_n6791.t231 vin_n.t155 vbn.t126 w_4660_n6791.t50 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X609 w_4660_n6791.t230 vin_n.t156 vbn.t125 w_4660_n6791.t70 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X610 vss.t120 voe1.t347 vout.t120 vss.t119 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X611 vdd.t101 iref.t163 vout.t210 vdd.t100 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X612 vdd.t99 iref.t164 vout.t232 vdd.t98 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X613 w_4660_n6791.t229 vin_n.t157 vbn.t124 w_4660_n6791.t50 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X614 w_4660_n6791.t228 vin_n.t158 vbn.t69 w_4660_n6791.t70 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X615 vss.t118 voe1.t348 vout.t138 vss.t117 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X616 vbn.t68 vin_n.t159 w_4660_n6791.t227 w_4660_n6791.t67 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X617 vss.t116 voe1.t349 vout.t96 vss.t115 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X618 vout.t217 iref.t165 vdd.t97 vdd.t96 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X619 vbn.t67 vin_n.t160 w_4660_n6791.t226 w_4660_n6791.t67 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X620 vdd.t95 iref.t166 vout.t272 vdd.t94 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X621 vss.t114 voe1.t350 vout.t191 vss.t113 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X622 vss.t112 voe1.t351 vout.t83 vss.t111 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X623 w_4660_n6791.t225 vin_n.t161 vbn.t66 w_4660_n6791.t52 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X624 vss.t110 voe1.t352 vout.t205 vss.t109 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X625 vout.t47 iref.t167 vdd.t93 vdd.t92 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X626 vdd.t91 iref.t168 vout.t27 vdd.t90 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X627 a_10611_n7515.t2 vdd.t318 voe1.t111 vss.t284 sky130_fd_pr__nfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=0.15
X628 voe1.t7 vin_p.t147 w_4660_n6791.t14 w_4660_n6791.t13 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X629 vout.t280 iref.t169 vdd.t89 vdd.t88 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X630 voe1.t16 vin_p.t148 w_4660_n6791.t28 w_4660_n6791.t13 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X631 vdd.t87 iref.t170 vout.t244 vdd.t86 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X632 vdd.t85 iref.t171 vout.t37 vdd.t84 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X633 vss.t108 voe1.t353 vout.t170 vss.t107 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X634 w_4660_n6791.t224 vin_n.t162 vbn.t145 w_4660_n6791.t163 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X635 vdd.t83 iref.t172 vout.t225 vdd.t82 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X636 w_4660_n6791.t223 vin_n.t163 vbn.t144 w_4660_n6791.t102 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X637 w_4660_n6791.t222 vin_n.t164 vbn.t143 w_4660_n6791.t112 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X638 vout.t304 a_10611_n7515.t7 sky130_fd_pr__cap_mim_m3_1 l=15 w=17.55
X639 voe1.t84 vbn.t284 vss.t270 vss.t269 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X640 vout.t289 iref.t173 vdd.t81 vdd.t80 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X641 w_4660_n6791.t221 vin_n.t165 vbn.t142 w_4660_n6791.t122 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X642 vdd.t79 iref.t174 vout.t32 vdd.t78 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X643 w_4660_n6791.t131 vin_p.t149 voe1.t89 w_4660_n6791.t130 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X644 w_4660_n6791.t220 vin_n.t166 vbn.t141 w_4660_n6791.t122 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X645 vdd.t77 iref.t175 w_4660_n6791.t473 vdd.t76 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X646 w_4660_n6791.t10 iref.t176 vdd.t75 vdd.t74 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X647 w_4660_n6791.t466 vin_p.t150 voe1.t221 w_4660_n6791.t130 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X648 voe1.t197 vin_p.t151 w_4660_n6791.t438 w_4660_n6791.t5 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X649 vdd.t73 iref.t177 vout.t248 vdd.t72 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X650 voe1.t180 vin_p.t152 w_4660_n6791.t420 w_4660_n6791.t5 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X651 w_4660_n6791.t219 vin_n.t167 vbn.t140 w_4660_n6791.t79 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X652 vss.t317 vbn.t285 voe1.t229 vss.t33 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X653 vdd.t71 iref.t16 iref.t17 vdd.t70 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X654 w_4660_n6791.t474 iref.t178 vdd.t69 vdd.t68 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X655 vout.t235 iref.t179 vdd.t67 vdd.t66 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X656 w_4660_n6791.t218 vin_n.t168 vbn.t139 w_4660_n6791.t102 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X657 w_4660_n6791.t217 vin_n.t169 vbn.t138 w_4660_n6791.t79 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X658 vss.t286 vbn.t286 voe1.t113 vss.t285 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X659 voe1.t92 vin_p.t153 w_4660_n6791.t134 w_4660_n6791.t45 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X660 voe1.t46 vin_p.t154 w_4660_n6791.t78 w_4660_n6791.t77 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X661 vout.t247 iref.t180 vdd.t65 vdd.t64 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X662 voe1.t206 vin_p.t155 w_4660_n6791.t447 w_4660_n6791.t77 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X663 voe1.t93 vin_p.t156 w_4660_n6791.t135 w_4660_n6791.t45 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X664 vdd.t63 iref.t181 vout.t14 vdd.t62 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X665 vss.t106 voe1.t354 vout.t103 vss.t105 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X666 vdd.t61 iref.t182 vout.t218 vdd.t60 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X667 vbn.t96 vin_n.t170 w_4660_n6791.t216 w_4660_n6791.t23 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X668 vbn.t95 vin_n.t171 w_4660_n6791.t215 w_4660_n6791.t83 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X669 w_4660_n6791.t214 vin_n.t172 vbn.t94 w_4660_n6791.t33 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X670 vss.t104 voe1.t355 vout.t68 vss.t103 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X671 vbn.t93 vin_n.t173 w_4660_n6791.t213 w_4660_n6791.t23 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X672 vbn.t178 vin_n.t174 w_4660_n6791.t212 w_4660_n6791.t83 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X673 voe1.t28 vbn.t287 vss.t20 vss.t19 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X674 w_4660_n6791.t211 vin_n.t175 vbn.t177 w_4660_n6791.t92 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X675 vout.t74 voe1.t356 vss.t102 vss.t101 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X676 w_4660_n6791.t455 vin_p.t157 voe1.t213 w_4660_n6791.t39 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X677 w_4660_n6791.t151 vin_p.t158 voe1.t109 w_4660_n6791.t148 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X678 vbn.t19 vbn.t18 vss.t316 vss.t307 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X679 w_4660_n6791.t149 vin_p.t159 voe1.t107 w_4660_n6791.t148 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X680 vss.t100 voe1.t357 vout.t92 vss.t99 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X681 w_4660_n6791.t428 vin_p.t160 voe1.t188 w_4660_n6791.t39 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X682 vbn.t17 vbn.t16 vss.t300 vss.t299 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X683 vout.t73 voe1.t358 vss.t98 vss.t97 sky130_fd_pr__nfet_01v8 ad=1.305 pd=9.58 as=0.6525 ps=4.79 w=4.5 l=0.45
X684 vout.t65 voe1.t359 vss.t96 vss.t95 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X685 vdd.t59 iref.t183 vout.t273 vdd.t58 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X686 w_4660_n6791.t210 vin_n.t176 vbn.t176 w_4660_n6791.t52 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X687 vout.t202 voe1.t360 vss.t94 vss.t93 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X688 vbn.t15 vbn.t14 vss.t297 vss.t296 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X689 w_4660_n6791.t209 vin_n.t177 vbn.t175 w_4660_n6791.t52 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X690 vss.t289 vbn.t288 voe1.t132 vss.t271 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X691 vout.t87 voe1.t361 vss.t92 vss.t91 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X692 vss.t90 voe1.t362 vout.t208 vss.t89 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X693 vout.t105 voe1.t363 vss.t88 vss.t87 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X694 vss.t38 vbn.t12 vbn.t13 vss.t0 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X695 w_4660_n6791.t427 vin_p.t161 voe1.t187 w_4660_n6791.t94 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X696 vss.t24 vbn.t10 vbn.t11 vss.t23 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X697 w_4660_n6791.t208 vin_n.t178 vbn.t182 w_4660_n6791.t37 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X698 w_4660_n6791.t479 vin_p.t162 voe1.t235 w_4660_n6791.t94 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X699 vout.t194 voe1.t364 vss.t86 vss.t85 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X700 vbn.t181 vin_n.t179 w_4660_n6791.t207 w_4660_n6791.t41 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X701 vss.t16 vbn.t8 vbn.t9 vss.t2 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X702 voe1.t133 vin_p.t163 w_4660_n6791.t173 w_4660_n6791.t118 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X703 vout.t305 a_10611_n7515.t6 sky130_fd_pr__cap_mim_m3_1 l=15 w=17.55
X704 vbn.t180 vin_n.t180 w_4660_n6791.t206 w_4660_n6791.t41 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X705 voe1.t90 vin_p.t164 w_4660_n6791.t132 w_4660_n6791.t118 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X706 vdd.t57 iref.t184 vout.t219 vdd.t56 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X707 voe1.t70 vin_p.t165 w_4660_n6791.t108 w_4660_n6791.t107 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X708 voe1.t27 vin_p.t166 w_4660_n6791.t48 w_4660_n6791.t47 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X709 vdd.t55 iref.t185 vout.t274 vdd.t54 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X710 vbn.t7 vbn.t6 vss.t304 vss.t8 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X711 voe1.t69 vin_p.t167 w_4660_n6791.t106 w_4660_n6791.t47 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X712 voe1.t233 vin_p.t168 w_4660_n6791.t477 w_4660_n6791.t107 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X713 vout.t169 voe1.t365 vss.t84 vss.t83 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X714 w_4660_n6791.t21 iref.t186 vdd.t5 vdd.t4 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X715 w_4660_n6791.t478 vin_p.t169 voe1.t234 w_4660_n6791.t88 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X716 vout.t281 iref.t187 vdd.t53 vdd.t52 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X717 w_4660_n6791.t205 vin_n.t181 vbn.t179 w_4660_n6791.t141 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X718 vbn.t5 vbn.t4 vss.t26 vss.t25 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X719 w_4660_n6791.t154 vin_p.t170 voe1.t116 w_4660_n6791.t144 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X720 w_4660_n6791.t204 vin_n.t182 vbn.t228 w_4660_n6791.t141 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X721 w_4660_n6791.t421 vin_p.t171 voe1.t181 w_4660_n6791.t88 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X722 w_4660_n6791.t145 vin_p.t172 voe1.t103 w_4660_n6791.t144 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X723 vout.t9 iref.t188 vdd.t51 vdd.t50 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X724 vdd.t49 iref.t189 vout.t249 vdd.t48 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X725 w_4660_n6791.t180 vin_p.t173 voe1.t144 w_4660_n6791.t60 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X726 w_4660_n6791.t71 vin_p.t174 voe1.t41 w_4660_n6791.t70 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X727 w_4660_n6791.t114 vin_p.t175 voe1.t74 w_4660_n6791.t50 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X728 vbn.t227 vin_n.t183 w_4660_n6791.t203 w_4660_n6791.t72 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X729 vdd.t47 iref.t190 vout.t263 vdd.t46 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X730 w_4660_n6791.t51 vin_p.t176 voe1.t31 w_4660_n6791.t50 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X731 w_4660_n6791.t439 vin_p.t177 voe1.t198 w_4660_n6791.t70 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X732 w_4660_n6791.t61 vin_p.t178 voe1.t36 w_4660_n6791.t60 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X733 vout.t264 iref.t191 vdd.t45 vdd.t44 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X734 voe1.t40 vin_p.t179 w_4660_n6791.t68 w_4660_n6791.t67 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X735 vout.t220 iref.t192 vdd.t43 vdd.t42 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X736 vdd.t41 iref.t193 vout.t275 vdd.t40 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X737 w_4660_n6791.t202 vin_n.t184 vbn.t226 w_4660_n6791.t130 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X738 voe1.t75 vin_p.t180 w_4660_n6791.t115 w_4660_n6791.t67 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X739 vdd.t39 iref.t194 vout.t28 vdd.t38 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X740 w_4660_n6791.t201 vin_n.t185 vbn.t225 w_4660_n6791.t64 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X741 vout.t133 voe1.t366 vss.t82 vss.t81 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X742 vss.t80 voe1.t367 vout.t89 vss.t79 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X743 vout.t282 iref.t195 vdd.t37 vdd.t36 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X744 w_4660_n6791.t200 vin_n.t186 vbn.t168 w_4660_n6791.t64 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X745 vout.t136 voe1.t368 vss.t78 vss.t77 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X746 vdd.t35 iref.t196 vout.t290 vdd.t34 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X747 vss.t76 voe1.t369 vout.t187 vss.t75 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X748 vout.t162 voe1.t370 vss.t74 vss.t73 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X749 vdd.t33 iref.t197 vout.t10 vdd.t32 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X750 vss.t72 voe1.t371 vout.t84 vss.t71 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X751 voe1.t57 vbn.t289 vss.t32 vss.t31 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X752 vout.t131 voe1.t372 vss.t70 vss.t69 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X753 vout.t86 voe1.t373 vss.t68 vss.t67 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X754 w_4660_n6791.t199 vin_n.t187 vbn.t167 w_4660_n6791.t98 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X755 vout.t144 voe1.t374 vss.t66 vss.t65 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X756 vdd.t31 iref.t198 vout.t250 vdd.t30 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X757 vout.t35 iref.t199 vdd.t29 vdd.t28 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X758 vout.t171 voe1.t375 vss.t64 vss.t63 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X759 w_4660_n6791.t123 vin_p.t181 voe1.t83 w_4660_n6791.t122 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X760 vdd.t27 iref.t200 vout.t209 vdd.t26 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X761 vout.t176 voe1.t376 vss.t62 vss.t61 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X762 vbn.t166 vin_n.t188 w_4660_n6791.t198 w_4660_n6791.t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X763 w_4660_n6791.t197 vin_n.t189 vbn.t165 w_4660_n6791.t92 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X764 w_4660_n6791.t463 vin_p.t182 voe1.t217 w_4660_n6791.t122 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X765 vbn.t221 vin_n.t190 w_4660_n6791.t196 w_4660_n6791.t11 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X766 vdd.t25 iref.t201 vout.t29 vdd.t24 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X767 vout.t161 voe1.t377 vss.t60 vss.t59 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X768 w_4660_n6791.t195 vin_n.t191 vbn.t220 w_4660_n6791.t92 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X769 vdd.t23 iref.t202 vout.t38 vdd.t22 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X770 w_4660_n6791.t22 iref.t203 vdd.t21 vdd.t20 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X771 vdd.t19 iref.t204 w_4660_n6791.t82 vdd.t18 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X772 w_4660_n6791.t194 vin_n.t192 vbn.t219 w_4660_n6791.t79 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X773 w_4660_n6791.t464 vin_p.t183 voe1.t218 w_4660_n6791.t79 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X774 vss.t268 vbn.t2 vbn.t3 vss.t17 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X775 w_4660_n6791.t462 vin_p.t184 voe1.t216 w_4660_n6791.t102 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X776 w_4660_n6791.t80 vin_p.t185 voe1.t47 w_4660_n6791.t79 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X777 vout.t128 voe1.t378 vss.t58 vss.t57 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X778 a_10611_n7515.t1 vdd.t319 voe1.t10 vss.t4 sky130_fd_pr__nfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=0.15
X779 w_4660_n6791.t128 vin_p.t186 voe1.t88 w_4660_n6791.t102 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X780 vdd.t17 iref.t205 vout.t291 vdd.t16 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X781 vdd.t15 iref.t26 iref.t27 vdd.t14 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X782 vout.t50 iref.t206 vdd.t13 vdd.t12 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X783 voe1.t112 vin_p.t187 w_4660_n6791.t152 w_4660_n6791.t62 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X784 voe1.t64 vin_p.t188 w_4660_n6791.t100 w_4660_n6791.t83 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X785 voe1.t13 vin_p.t189 w_4660_n6791.t24 w_4660_n6791.t23 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X786 vbn.t1 vbn.t0 vss.t306 vss.t302 sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X787 voe1.t215 vin_p.t190 w_4660_n6791.t458 w_4660_n6791.t23 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X788 voe1.t50 vin_p.t191 w_4660_n6791.t84 w_4660_n6791.t83 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X789 iref.t11 iref.t10 vdd.t11 vdd.t10 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X790 vdd.t9 iref.t207 w_4660_n6791.t129 vdd.t8 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X791 voe1.t231 vin_p.t192 w_4660_n6791.t475 w_4660_n6791.t62 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X792 vbn.t218 vin_n.t193 w_4660_n6791.t193 w_4660_n6791.t2 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X793 vbn.t85 vin_n.t194 w_4660_n6791.t192 w_4660_n6791.t67 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X794 vss.t56 voe1.t379 vout.t88 vss.t55 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X795 voe1.t209 vin_p.t193 w_4660_n6791.t450 w_4660_n6791.t43 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X796 vbn.t84 vin_n.t195 w_4660_n6791.t191 w_4660_n6791.t2 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X797 vbn.t83 vin_n.t196 w_4660_n6791.t190 w_4660_n6791.t2 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X798 vdd.t3 iref.t2 iref.t3 vdd.t2 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X799 voe1.t25 vin_p.t194 w_4660_n6791.t44 w_4660_n6791.t43 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X800 vbn.t82 vin_n.t197 w_4660_n6791.t189 w_4660_n6791.t2 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X801 w_4660_n6791.t121 vin_p.t195 voe1.t82 w_4660_n6791.t30 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X802 w_4660_n6791.t54 vin_p.t196 voe1.t33 w_4660_n6791.t52 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X803 w_4660_n6791.t53 vin_p.t197 voe1.t32 w_4660_n6791.t52 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X804 a_10611_n7515.t0 vdd.t320 voe1.t110 vss.t283 sky130_fd_pr__nfet_01v8 ad=0.2175 pd=2.08 as=0.2175 ps=2.08 w=0.75 l=0.15
X805 vout.t175 voe1.t380 vss.t54 vss.t53 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X806 vss.t52 voe1.t381 vout.t125 vss.t51 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X807 w_4660_n6791.t31 vin_p.t198 voe1.t18 w_4660_n6791.t30 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X808 vout.t134 voe1.t382 vss.t50 vss.t49 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X809 vdd.t7 iref.t208 vout.t58 vdd.t6 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X810 w_4660_n6791.t188 vin_n.t198 vbn.t244 w_4660_n6791.t33 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X811 vss.t48 voe1.t383 vout.t174 vss.t47 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X812 vdd.t1 iref.t209 vout.t33 vdd.t0 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X813 w_4660_n6791.t187 vin_n.t199 vbn.t243 w_4660_n6791.t33 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X814 vout.t108 voe1.t384 vss.t46 vss.t45 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X815 vout.t113 voe1.t385 vss.t44 vss.t43 sky130_fd_pr__nfet_01v8 ad=0.6525 pd=4.79 as=0.6525 ps=4.79 w=4.5 l=0.45
X816 voe1.t91 vin_p.t199 w_4660_n6791.t133 w_4660_n6791.t41 sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
R0 voe1.n81 voe1.t243 294.981
R1 voe1.n81 voe1.t304 294.981
R2 voe1.n80 voe1.t369 294.981
R3 voe1.n80 voe1.t277 294.981
R4 voe1.n79 voe1.t268 294.981
R5 voe1.n79 voe1.t322 294.981
R6 voe1.n78 voe1.t346 294.981
R7 voe1.n78 voe1.t247 294.981
R8 voe1.n77 voe1.t238 294.981
R9 voe1.n77 voe1.t298 294.981
R10 voe1.n76 voe1.t334 294.981
R11 voe1.n76 voe1.t236 294.981
R12 voe1.n75 voe1.t261 294.981
R13 voe1.n75 voe1.t318 294.981
R14 voe1.n74 voe1.t357 294.981
R15 voe1.n74 voe1.t259 294.981
R16 voe1.n73 voe1.t255 294.981
R17 voe1.n73 voe1.t312 294.981
R18 voe1.n72 voe1.t351 294.981
R19 voe1.n72 voe1.t253 294.981
R20 voe1.n71 voe1.t375 294.981
R21 voe1.n71 voe1.t284 294.981
R22 voe1.n70 voe1.t354 294.981
R23 voe1.n70 voe1.t257 294.981
R24 voe1.n69 voe1.t251 294.981
R25 voe1.n69 voe1.t309 294.981
R26 voe1.n68 voe1.t347 294.981
R27 voe1.n68 voe1.t248 294.981
R28 voe1.n67 voe1.t242 294.981
R29 voe1.n67 voe1.t302 294.981
R30 voe1.n66 voe1.t337 294.981
R31 voe1.n66 voe1.t239 294.981
R32 voe1.n65 voe1.t265 294.981
R33 voe1.n65 voe1.t321 294.981
R34 voe1.n64 voe1.t299 294.981
R35 voe1.n64 voe1.t349 294.981
R36 voe1.n63 voe1.t237 294.981
R37 voe1.n63 voe1.t296 294.981
R38 voe1.n62 voe1.t289 294.981
R39 voe1.n62 voe1.t340 294.981
R40 voe1.n61 voe1.t377 294.981
R41 voe1.n61 voe1.t287 294.981
R42 voe1.n60 voe1.t313 294.981
R43 voe1.n60 voe1.t362 294.981
R44 voe1.n59 voe1.t254 294.981
R45 voe1.n59 voe1.t311 294.981
R46 voe1.n58 voe1.t305 294.981
R47 voe1.n58 voe1.t353 294.981
R48 voe1.n57 voe1.t373 294.981
R49 voe1.n57 voe1.t280 294.981
R50 voe1.n56 voe1.t271 294.981
R51 voe1.n56 voe1.t325 294.981
R52 voe1.n55 voe1.t249 294.981
R53 voe1.n55 voe1.t307 294.981
R54 voe1.n54 voe1.t303 294.981
R55 voe1.n54 voe1.t352 294.981
R56 voe1.n53 voe1.t240 294.981
R57 voe1.n53 voe1.t300 294.981
R58 voe1.n52 voe1.t291 294.981
R59 voe1.n52 voe1.t342 294.981
R60 voe1.n51 voe1.t359 294.981
R61 voe1.n51 voe1.t262 294.981
R62 voe1.n50 voe1.t297 294.981
R63 voe1.n50 voe1.t348 294.981
R64 voe1.n49 voe1.t384 294.981
R65 voe1.n49 voe1.t294 294.981
R66 voe1.n48 voe1.t288 294.981
R67 voe1.n48 voe1.t338 294.981
R68 voe1.n47 voe1.t376 294.981
R69 voe1.n47 voe1.t285 294.981
R70 voe1.n46 voe1.t273 294.981
R71 voe1.n46 voe1.t327 294.981
R72 voe1.n45 voe1.t252 294.981
R73 voe1.n45 voe1.t310 294.981
R74 voe1.n44 voe1.t281 294.981
R75 voe1.n44 voe1.t333 294.981
R76 voe1.n43 voe1.t370 294.981
R77 voe1.n43 voe1.t278 294.981
R78 voe1.n42 voe1.t269 294.981
R79 voe1.n42 voe1.t323 294.981
R80 voe1.n41 voe1.t361 294.981
R81 voe1.n41 voe1.t266 294.981
R82 voe1.n40 voe1.t301 294.981
R83 voe1.n40 voe1.t350 294.981
R84 voe1.n39 voe1.t343 294.981
R85 voe1.n39 voe1.t244 294.981
R86 voe1.n38 voe1.t290 294.981
R87 voe1.n38 voe1.t341 294.981
R88 voe1.n37 voe1.t315 294.981
R89 voe1.n37 voe1.t364 294.981
R90 voe1.n36 voe1.t256 294.981
R91 voe1.n36 voe1.t314 294.981
R92 voe1.n35 voe1.t339 294.981
R93 voe1.n35 voe1.t241 294.981
R94 voe1.n34 voe1.t286 294.981
R95 voe1.n34 voe1.t336 294.981
R96 voe1.n33 voe1.t328 294.981
R97 voe1.n33 voe1.t378 294.981
R98 voe1.n32 voe1.t272 294.981
R99 voe1.n32 voe1.t326 294.981
R100 voe1.n31 voe1.t316 294.981
R101 voe1.n31 voe1.t365 294.981
R102 voe1.n30 voe1.t344 294.981
R103 voe1.n30 voe1.t245 294.981
R104 voe1.n29 voe1.t382 294.981
R105 voe1.n29 voe1.t293 294.981
R106 voe1.n28 voe1.t330 294.981
R107 voe1.n28 voe1.t381 294.981
R108 voe1.n27 voe1.t374 294.981
R109 voe1.n27 voe1.t283 294.981
R110 voe1.n26 voe1.t319 294.981
R111 voe1.n26 voe1.t371 294.981
R112 voe1.n25 voe1.t250 294.981
R113 voe1.n25 voe1.t308 294.981
R114 voe1.n24 voe1.t329 294.981
R115 voe1.n24 voe1.t379 294.981
R116 voe1.n23 voe1.t368 294.981
R117 voe1.n23 voe1.t276 294.981
R118 voe1.n22 voe1.t317 294.981
R119 voe1.n22 voe1.t367 294.981
R120 voe1.n21 voe1.t360 294.981
R121 voe1.n21 voe1.t264 294.981
R122 voe1.n20 voe1.t345 294.981
R123 voe1.n20 voe1.t246 294.981
R124 voe1.n19 voe1.t385 294.981
R125 voe1.n19 voe1.t295 294.981
R126 voe1.n18 voe1.t332 294.981
R127 voe1.n18 voe1.t383 294.981
R128 voe1.n17 voe1.t356 294.981
R129 voe1.n17 voe1.t258 294.981
R130 voe1.n16 voe1.t306 294.981
R131 voe1.n16 voe1.t355 294.981
R132 voe1.n15 voe1.t380 294.981
R133 voe1.n15 voe1.t292 294.981
R134 voe1.n14 voe1.t282 294.981
R135 voe1.n14 voe1.t335 294.981
R136 voe1.n13 voe1.t372 294.981
R137 voe1.n13 voe1.t279 294.981
R138 voe1.n12 voe1.t270 294.981
R139 voe1.n12 voe1.t324 294.981
R140 voe1.n11 voe1.t363 294.981
R141 voe1.n11 voe1.t267 294.981
R142 voe1.n10 voe1.t275 294.981
R143 voe1.n10 voe1.t331 294.981
R144 voe1.n9 voe1.t366 294.981
R145 voe1.n9 voe1.t274 294.981
R146 voe1.n8 voe1.t263 294.981
R147 voe1.n8 voe1.t320 294.981
R148 voe1.n7 voe1.t358 294.981
R149 voe1.n7 voe1.t260 294.981
R150 voe1.n5 voe1.t10 129.55
R151 voe1.n1 voe1.t111 124.24
R152 voe1.n5 voe1.t12 123.966
R153 voe1.n5 voe1.t110 123.966
R154 voe1.n5 voe1.t77 123.966
R155 voe1.n5 voe1.t78 123.966
R156 voe1.n5 voe1.n159 75.3571
R157 voe1.n6 voe1.n85 75.3571
R158 voe1.n5 voe1.n110 75.3571
R159 voe1.n5 voe1.n135 75.3571
R160 voe1.n6 voe1.n108 75.3477
R161 voe1.n5 voe1.n133 75.3477
R162 voe1.n5 voe1.n158 75.3477
R163 voe1.n5 voe1.n183 75.3477
R164 voe1.n5 voe1.n160 75.3376
R165 voe1.n5 voe1.n161 75.3376
R166 voe1.n5 voe1.n162 75.3376
R167 voe1.n5 voe1.n163 75.3376
R168 voe1.n5 voe1.n164 75.3376
R169 voe1.n5 voe1.n165 75.3376
R170 voe1.n5 voe1.n166 75.3376
R171 voe1.n5 voe1.n167 75.3376
R172 voe1.n5 voe1.n169 75.3376
R173 voe1.n5 voe1.n170 75.3376
R174 voe1.n5 voe1.n171 75.3376
R175 voe1.n5 voe1.n172 75.3376
R176 voe1.n6 voe1.n86 75.3376
R177 voe1.n6 voe1.n87 75.3376
R178 voe1.n6 voe1.n88 75.3376
R179 voe1.n6 voe1.n89 75.3376
R180 voe1.n6 voe1.n90 75.3376
R181 voe1.n6 voe1.n91 75.3376
R182 voe1.n6 voe1.n92 75.3376
R183 voe1.n6 voe1.n93 75.3376
R184 voe1.n6 voe1.n94 75.3376
R185 voe1.n6 voe1.n95 75.3376
R186 voe1.n6 voe1.n96 75.3376
R187 voe1.n6 voe1.n97 75.3376
R188 voe1.n6 voe1.n84 75.3376
R189 voe1.n6 voe1.n99 75.3376
R190 voe1.n6 voe1.n98 75.3376
R191 voe1.n6 voe1.n101 75.3376
R192 voe1.n6 voe1.n100 75.3376
R193 voe1.n6 voe1.n103 75.3376
R194 voe1.n6 voe1.n102 75.3376
R195 voe1.n6 voe1.n105 75.3376
R196 voe1.n6 voe1.n104 75.3376
R197 voe1.n6 voe1.n107 75.3376
R198 voe1.n6 voe1.n106 75.3376
R199 voe1.n5 voe1.n111 75.3376
R200 voe1.n5 voe1.n112 75.3376
R201 voe1.n5 voe1.n113 75.3376
R202 voe1.n5 voe1.n114 75.3376
R203 voe1.n5 voe1.n115 75.3376
R204 voe1.n5 voe1.n116 75.3376
R205 voe1.n5 voe1.n117 75.3376
R206 voe1.n5 voe1.n118 75.3376
R207 voe1.n5 voe1.n119 75.3376
R208 voe1.n5 voe1.n120 75.3376
R209 voe1.n5 voe1.n121 75.3376
R210 voe1.n5 voe1.n122 75.3376
R211 voe1.n5 voe1.n109 75.3376
R212 voe1.n5 voe1.n124 75.3376
R213 voe1.n5 voe1.n123 75.3376
R214 voe1.n5 voe1.n126 75.3376
R215 voe1.n5 voe1.n125 75.3376
R216 voe1.n5 voe1.n128 75.3376
R217 voe1.n5 voe1.n127 75.3376
R218 voe1.n5 voe1.n130 75.3376
R219 voe1.n5 voe1.n129 75.3376
R220 voe1.n5 voe1.n132 75.3376
R221 voe1.n5 voe1.n131 75.3376
R222 voe1.n5 voe1.n136 75.3376
R223 voe1.n5 voe1.n137 75.3376
R224 voe1.n5 voe1.n138 75.3376
R225 voe1.n5 voe1.n139 75.3376
R226 voe1.n5 voe1.n140 75.3376
R227 voe1.n5 voe1.n141 75.3376
R228 voe1.n5 voe1.n142 75.3376
R229 voe1.n5 voe1.n143 75.3376
R230 voe1.n5 voe1.n144 75.3376
R231 voe1.n5 voe1.n145 75.3376
R232 voe1.n5 voe1.n146 75.3376
R233 voe1.n5 voe1.n147 75.3376
R234 voe1.n5 voe1.n134 75.3376
R235 voe1.n5 voe1.n149 75.3376
R236 voe1.n5 voe1.n148 75.3376
R237 voe1.n5 voe1.n151 75.3376
R238 voe1.n5 voe1.n150 75.3376
R239 voe1.n5 voe1.n153 75.3376
R240 voe1.n5 voe1.n152 75.3376
R241 voe1.n5 voe1.n155 75.3376
R242 voe1.n5 voe1.n154 75.3376
R243 voe1.n5 voe1.n157 75.3376
R244 voe1.n5 voe1.n156 75.3376
R245 voe1.n5 voe1.n174 75.3376
R246 voe1.n5 voe1.n173 75.3376
R247 voe1.n5 voe1.n176 75.3376
R248 voe1.n5 voe1.n175 75.3376
R249 voe1.n5 voe1.n178 75.3376
R250 voe1.n5 voe1.n177 75.3376
R251 voe1.n5 voe1.n180 75.3376
R252 voe1.n5 voe1.n179 75.3376
R253 voe1.n5 voe1.n182 75.3376
R254 voe1.n5 voe1.n181 75.3376
R255 voe1.n5 voe1.n168 75.3376
R256 voe1.n4 voe1.n7 70.7757
R257 voe1.n1 voe1.n81 70.6694
R258 voe1.n1 voe1.n80 70.6694
R259 voe1.n1 voe1.n79 70.6694
R260 voe1.n1 voe1.n78 70.6694
R261 voe1.n1 voe1.n77 70.6694
R262 voe1.n1 voe1.n76 70.6694
R263 voe1.n1 voe1.n75 70.6694
R264 voe1.n1 voe1.n74 70.6694
R265 voe1.n1 voe1.n73 70.6694
R266 voe1.n1 voe1.n72 70.6694
R267 voe1.n1 voe1.n71 70.6694
R268 voe1.n1 voe1.n70 70.6694
R269 voe1.n1 voe1.n69 70.6694
R270 voe1.n1 voe1.n68 70.6694
R271 voe1.n1 voe1.n67 70.6694
R272 voe1.n1 voe1.n66 70.6694
R273 voe1.n0 voe1.n65 70.6694
R274 voe1.n0 voe1.n64 70.6694
R275 voe1.n0 voe1.n63 70.6694
R276 voe1.n0 voe1.n62 70.6694
R277 voe1.n0 voe1.n61 70.6694
R278 voe1.n0 voe1.n60 70.6694
R279 voe1.n0 voe1.n59 70.6694
R280 voe1.n0 voe1.n58 70.6694
R281 voe1.n0 voe1.n57 70.6694
R282 voe1.n0 voe1.n56 70.6694
R283 voe1.n0 voe1.n55 70.6694
R284 voe1.n0 voe1.n54 70.6694
R285 voe1.n0 voe1.n53 70.6694
R286 voe1.n0 voe1.n52 70.6694
R287 voe1.n0 voe1.n51 70.6694
R288 voe1.n0 voe1.n50 70.6694
R289 voe1.n2 voe1.n49 70.6694
R290 voe1.n2 voe1.n48 70.6694
R291 voe1.n2 voe1.n47 70.6694
R292 voe1.n2 voe1.n46 70.6694
R293 voe1.n2 voe1.n45 70.6694
R294 voe1.n2 voe1.n44 70.6694
R295 voe1.n2 voe1.n43 70.6694
R296 voe1.n2 voe1.n42 70.6694
R297 voe1.n2 voe1.n41 70.6694
R298 voe1.n2 voe1.n40 70.6694
R299 voe1.n2 voe1.n39 70.6694
R300 voe1.n2 voe1.n38 70.6694
R301 voe1.n2 voe1.n37 70.6694
R302 voe1.n2 voe1.n36 70.6694
R303 voe1.n2 voe1.n35 70.6694
R304 voe1.n2 voe1.n34 70.6694
R305 voe1.n3 voe1.n33 70.6694
R306 voe1.n3 voe1.n32 70.6694
R307 voe1.n3 voe1.n31 70.6694
R308 voe1.n3 voe1.n30 70.6694
R309 voe1.n3 voe1.n29 70.6694
R310 voe1.n3 voe1.n28 70.6694
R311 voe1.n3 voe1.n27 70.6694
R312 voe1.n3 voe1.n26 70.6694
R313 voe1.n3 voe1.n25 70.6694
R314 voe1.n3 voe1.n24 70.6694
R315 voe1.n3 voe1.n23 70.6694
R316 voe1.n3 voe1.n22 70.6694
R317 voe1.n3 voe1.n21 70.6694
R318 voe1.n3 voe1.n20 70.6694
R319 voe1.n3 voe1.n19 70.6694
R320 voe1.n3 voe1.n18 70.6694
R321 voe1.n4 voe1.n17 70.6694
R322 voe1.n4 voe1.n16 70.6694
R323 voe1.n4 voe1.n15 70.6694
R324 voe1.n4 voe1.n14 70.6694
R325 voe1.n4 voe1.n13 70.6694
R326 voe1.n4 voe1.n12 70.6694
R327 voe1.n4 voe1.n11 70.6694
R328 voe1.n4 voe1.n10 70.6694
R329 voe1.n4 voe1.n9 70.6694
R330 voe1.n4 voe1.n8 70.6694
R331 voe1.n5 voe1.t29 31.9205
R332 voe1.n5 voe1.t199 31.1376
R333 voe1.n5 voe1.n83 26.1251
R334 voe1.n5 voe1.n189 25.8248
R335 voe1.n5 voe1.n184 25.8248
R336 voe1.n5 voe1.n188 25.8248
R337 voe1.n5 voe1.n185 25.8248
R338 voe1.n5 voe1.n187 25.8248
R339 voe1.n5 voe1.n186 25.8248
R340 voe1.n5 voe1.n191 25.3811
R341 voe1.n5 voe1.n190 25.3376
R342 voe1.n5 voe1.n193 25.3376
R343 voe1.n5 voe1.n192 25.3376
R344 voe1.n5 voe1.n195 25.3376
R345 voe1.n5 voe1.n194 25.3376
R346 voe1.n5 voe1.n82 25.3376
R347 voe1.n159 voe1.t194 9.52217
R348 voe1.n159 voe1.t185 9.52217
R349 voe1.n160 voe1.t60 9.52217
R350 voe1.n160 voe1.t171 9.52217
R351 voe1.n161 voe1.t89 9.52217
R352 voe1.n161 voe1.t7 9.52217
R353 voe1.n162 voe1.t213 9.52217
R354 voe1.n162 voe1.t92 9.52217
R355 voe1.n163 voe1.t38 9.52217
R356 voe1.n163 voe1.t3 9.52217
R357 voe1.n164 voe1.t95 9.52217
R358 voe1.n164 voe1.t102 9.52217
R359 voe1.n165 voe1.t99 9.52217
R360 voe1.n165 voe1.t24 9.52217
R361 voe1.n166 voe1.t172 9.52217
R362 voe1.n166 voe1.t34 9.52217
R363 voe1.n167 voe1.t207 9.52217
R364 voe1.n167 voe1.t173 9.52217
R365 voe1.n169 voe1.t73 9.52217
R366 voe1.n169 voe1.t175 9.52217
R367 voe1.n170 voe1.t170 9.52217
R368 voe1.n170 voe1.t6 9.52217
R369 voe1.n171 voe1.t122 9.52217
R370 voe1.n171 voe1.t209 9.52217
R371 voe1.n172 voe1.t54 9.52217
R372 voe1.n172 voe1.t124 9.52217
R373 voe1.n85 voe1.t107 9.52217
R374 voe1.n85 voe1.t206 9.52217
R375 voe1.n86 voe1.t149 9.52217
R376 voe1.n86 voe1.t71 9.52217
R377 voe1.n87 voe1.t96 9.52217
R378 voe1.n87 voe1.t228 9.52217
R379 voe1.n88 voe1.t23 9.52217
R380 voe1.n88 voe1.t145 9.52217
R381 voe1.n89 voe1.t150 9.52217
R382 voe1.n89 voe1.t180 9.52217
R383 voe1.n90 voe1.t32 9.52217
R384 voe1.n90 voe1.t215 9.52217
R385 voe1.n91 voe1.t212 9.52217
R386 voe1.n91 voe1.t232 9.52217
R387 voe1.n92 voe1.t131 9.52217
R388 voe1.n92 voe1.t17 9.52217
R389 voe1.n93 voe1.t148 9.52217
R390 voe1.n93 voe1.t136 9.52217
R391 voe1.n94 voe1.t31 9.52217
R392 voe1.n94 voe1.t115 9.52217
R393 voe1.n95 voe1.t129 9.52217
R394 voe1.n95 voe1.t205 9.52217
R395 voe1.n96 voe1.t142 9.52217
R396 voe1.n96 voe1.t120 9.52217
R397 voe1.n97 voe1.t47 9.52217
R398 voe1.n97 voe1.t155 9.52217
R399 voe1.n84 voe1.t181 9.52217
R400 voe1.n84 voe1.t50 9.52217
R401 voe1.n99 voe1.t35 9.52217
R402 voe1.n99 voe1.t75 9.52217
R403 voe1.n98 voe1.t66 9.52217
R404 voe1.n98 voe1.t203 9.52217
R405 voe1.n101 voe1.t160 9.52217
R406 voe1.n101 voe1.t37 9.52217
R407 voe1.n100 voe1.t198 9.52217
R408 voe1.n100 voe1.t69 9.52217
R409 voe1.n103 voe1.t183 9.52217
R410 voe1.n103 voe1.t1 9.52217
R411 voe1.n102 voe1.t179 9.52217
R412 voe1.n102 voe1.t19 9.52217
R413 voe1.n105 voe1.t162 9.52217
R414 voe1.n105 voe1.t146 9.52217
R415 voe1.n104 voe1.t103 9.52217
R416 voe1.n104 voe1.t90 9.52217
R417 voe1.n107 voe1.t184 9.52217
R418 voe1.n107 voe1.t196 9.52217
R419 voe1.n106 voe1.t156 9.52217
R420 voe1.n106 voe1.t15 9.52217
R421 voe1.n108 voe1.t217 9.52217
R422 voe1.n108 voe1.t76 9.52217
R423 voe1.n110 voe1.t109 9.52217
R424 voe1.n110 voe1.t46 9.52217
R425 voe1.n111 voe1.t151 9.52217
R426 voe1.n111 voe1.t130 9.52217
R427 voe1.n112 voe1.t141 9.52217
R428 voe1.n112 voe1.t97 9.52217
R429 voe1.n113 voe1.t44 9.52217
R430 voe1.n113 voe1.t26 9.52217
R431 voe1.n114 voe1.t67 9.52217
R432 voe1.n114 voe1.t197 9.52217
R433 voe1.n115 voe1.t33 9.52217
R434 voe1.n115 voe1.t13 9.52217
R435 voe1.n116 voe1.t167 9.52217
R436 voe1.n116 voe1.t91 9.52217
R437 voe1.n117 voe1.t63 9.52217
R438 voe1.n117 voe1.t211 9.52217
R439 voe1.n118 voe1.t108 9.52217
R440 voe1.n118 voe1.t42 9.52217
R441 voe1.n119 voe1.t74 9.52217
R442 voe1.n119 voe1.t86 9.52217
R443 voe1.n120 voe1.t119 9.52217
R444 voe1.n120 voe1.t128 9.52217
R445 voe1.n121 voe1.t125 9.52217
R446 voe1.n121 voe1.t52 9.52217
R447 voe1.n122 voe1.t218 9.52217
R448 voe1.n122 voe1.t164 9.52217
R449 voe1.n109 voe1.t234 9.52217
R450 voe1.n109 voe1.t64 9.52217
R451 voe1.n124 voe1.t22 9.52217
R452 voe1.n124 voe1.t40 9.52217
R453 voe1.n123 voe1.t106 9.52217
R454 voe1.n123 voe1.t79 9.52217
R455 voe1.n126 voe1.t153 9.52217
R456 voe1.n126 voe1.t161 9.52217
R457 voe1.n125 voe1.t41 9.52217
R458 voe1.n125 voe1.t27 9.52217
R459 voe1.n128 voe1.t20 9.52217
R460 voe1.n128 voe1.t2 9.52217
R461 voe1.n127 voe1.t61 9.52217
R462 voe1.n127 voe1.t4 9.52217
R463 voe1.n130 voe1.t65 9.52217
R464 voe1.n130 voe1.t186 9.52217
R465 voe1.n129 voe1.t116 9.52217
R466 voe1.n129 voe1.t133 9.52217
R467 voe1.n132 voe1.t127 9.52217
R468 voe1.n132 voe1.t182 9.52217
R469 voe1.n131 voe1.t157 9.52217
R470 voe1.n131 voe1.t14 9.52217
R471 voe1.n133 voe1.t83 9.52217
R472 voe1.n133 voe1.t9 9.52217
R473 voe1.n135 voe1.t195 9.52217
R474 voe1.n135 voe1.t193 9.52217
R475 voe1.n136 voe1.t147 9.52217
R476 voe1.n136 voe1.t72 9.52217
R477 voe1.n137 voe1.t221 9.52217
R478 voe1.n137 voe1.t16 9.52217
R479 voe1.n138 voe1.t188 9.52217
R480 voe1.n138 voe1.t93 9.52217
R481 voe1.n139 voe1.t45 9.52217
R482 voe1.n139 voe1.t5 9.52217
R483 voe1.n140 voe1.t43 9.52217
R484 voe1.n140 voe1.t140 9.52217
R485 voe1.n141 voe1.t200 9.52217
R486 voe1.n141 voe1.t143 9.52217
R487 voe1.n142 voe1.t152 9.52217
R488 voe1.n142 voe1.t8 9.52217
R489 voe1.n143 voe1.t21 9.52217
R490 voe1.n143 voe1.t168 9.52217
R491 voe1.n144 voe1.t55 9.52217
R492 voe1.n144 voe1.t169 9.52217
R493 voe1.n145 voe1.t210 9.52217
R494 voe1.n145 voe1.t202 9.52217
R495 voe1.n146 voe1.t134 9.52217
R496 voe1.n146 voe1.t30 9.52217
R497 voe1.n147 voe1.t123 9.52217
R498 voe1.n147 voe1.t25 9.52217
R499 voe1.n134 voe1.t118 9.52217
R500 voe1.n134 voe1.t98 9.52217
R501 voe1.n149 voe1.t154 9.52217
R502 voe1.n149 voe1.t190 9.52217
R503 voe1.n148 voe1.t88 9.52217
R504 voe1.n148 voe1.t53 9.52217
R505 voe1.n151 voe1.t18 9.52217
R506 voe1.n151 voe1.t231 9.52217
R507 voe1.n150 voe1.t87 9.52217
R508 voe1.n150 voe1.t81 9.52217
R509 voe1.n153 voe1.t39 9.52217
R510 voe1.n153 voe1.t176 9.52217
R511 voe1.n152 voe1.t235 9.52217
R512 voe1.n152 voe1.t178 9.52217
R513 voe1.n155 voe1.t36 9.52217
R514 voe1.n155 voe1.t233 9.52217
R515 voe1.n154 voe1.t117 9.52217
R516 voe1.n154 voe1.t80 9.52217
R517 voe1.n157 voe1.t174 9.52217
R518 voe1.n157 voe1.t158 9.52217
R519 voe1.n156 voe1.t166 9.52217
R520 voe1.n156 voe1.t219 9.52217
R521 voe1.n158 voe1.t121 9.52217
R522 voe1.n158 voe1.t177 9.52217
R523 voe1.n174 voe1.t163 9.52217
R524 voe1.n174 voe1.t56 9.52217
R525 voe1.n173 voe1.t216 9.52217
R526 voe1.n173 voe1.t208 9.52217
R527 voe1.n176 voe1.t82 9.52217
R528 voe1.n176 voe1.t112 9.52217
R529 voe1.n175 voe1.t191 9.52217
R530 voe1.n175 voe1.t204 9.52217
R531 voe1.n178 voe1.t201 9.52217
R532 voe1.n178 voe1.t49 9.52217
R533 voe1.n177 voe1.t187 9.52217
R534 voe1.n177 voe1.t68 9.52217
R535 voe1.n180 voe1.t144 9.52217
R536 voe1.n180 voe1.t70 9.52217
R537 voe1.n179 voe1.t192 9.52217
R538 voe1.n179 voe1.t189 9.52217
R539 voe1.n182 voe1.t227 9.52217
R540 voe1.n182 voe1.t159 9.52217
R541 voe1.n181 voe1.t165 9.52217
R542 voe1.n181 voe1.t214 9.52217
R543 voe1.n183 voe1.t94 9.52217
R544 voe1.n183 voe1.t62 9.52217
R545 voe1.n168 voe1.t126 9.52217
R546 voe1.n168 voe1.t0 9.52217
R547 voe1.n189 voe1.t51 5.8005
R548 voe1.n189 voe1.t135 5.8005
R549 voe1.n184 voe1.t58 5.8005
R550 voe1.n184 voe1.t225 5.8005
R551 voe1.n188 voe1.t113 5.8005
R552 voe1.n188 voe1.t84 5.8005
R553 voe1.n185 voe1.t132 5.8005
R554 voe1.n185 voe1.t28 5.8005
R555 voe1.n187 voe1.t223 5.8005
R556 voe1.n187 voe1.t226 5.8005
R557 voe1.n186 voe1.t11 5.8005
R558 voe1.n186 voe1.t230 5.8005
R559 voe1.n83 voe1.t101 5.8005
R560 voe1.n83 voe1.t57 5.8005
R561 voe1.n191 voe1.t100 5.8005
R562 voe1.n191 voe1.t59 5.8005
R563 voe1.n190 voe1.t138 5.8005
R564 voe1.n190 voe1.t48 5.8005
R565 voe1.n193 voe1.t229 5.8005
R566 voe1.n193 voe1.t137 5.8005
R567 voe1.n192 voe1.t224 5.8005
R568 voe1.n192 voe1.t105 5.8005
R569 voe1.n195 voe1.t85 5.8005
R570 voe1.n195 voe1.t139 5.8005
R571 voe1.n194 voe1.t114 5.8005
R572 voe1.n194 voe1.t104 5.8005
R573 voe1.n82 voe1.t222 5.8005
R574 voe1.n82 voe1.t220 5.8005
R575 voe1.n5 voe1.n1 2.15113
R576 voe1.n5 voe1.n6 1.70285
R577 voe1.n2 voe1.n3 1.70165
R578 voe1.n0 voe1.n2 1.70165
R579 voe1.n1 voe1.n0 1.70165
R580 voe1.n3 voe1.n4 1.59533
R581 vout.n270 vout.t226 85.9418
R582 vout.n230 vout.t297 85.9418
R583 vout.n183 vout.t283 85.9418
R584 vout.n270 vout.t214 85.3464
R585 vout.n230 vout.t241 85.3464
R586 vout.n183 vout.t246 85.3464
R587 vout.n274 vout.n272 76.4201
R588 vout.n268 vout.n266 76.4201
R589 vout.n285 vout.n283 76.4201
R590 vout.n263 vout.n261 76.4201
R591 vout.n258 vout.n256 76.4201
R592 vout.n302 vout.n300 76.4201
R593 vout.n252 vout.n250 76.4201
R594 vout.n247 vout.n245 76.4201
R595 vout.n318 vout.n316 76.4201
R596 vout.n242 vout.n240 76.4201
R597 vout.n237 vout.n235 76.4201
R598 vout.n234 vout.n232 76.4201
R599 vout.n227 vout.n225 76.4201
R600 vout.n344 vout.n342 76.4201
R601 vout.n222 vout.n220 76.4201
R602 vout.n217 vout.n215 76.4201
R603 vout.n209 vout.n207 76.4201
R604 vout.n366 vout.n364 76.4201
R605 vout.n206 vout.n204 76.4201
R606 vout.n201 vout.n199 76.4201
R607 vout.n383 vout.n381 76.4201
R608 vout.n196 vout.n194 76.4201
R609 vout.n191 vout.n189 76.4201
R610 vout.n188 vout.n186 76.4201
R611 vout.n405 vout.n403 76.4201
R612 vout.n180 vout.n178 76.4201
R613 vout.n175 vout.n173 76.4201
R614 vout.n421 vout.n419 76.4201
R615 vout.n170 vout.n168 76.4201
R616 vout.n432 vout.n430 76.4201
R617 vout.n165 vout.n163 76.4201
R618 vout.n440 vout.n438 76.4201
R619 vout.n445 vout.n443 76.4201
R620 vout.n450 vout.n448 76.4201
R621 vout.n454 vout.n452 76.4201
R622 vout.n457 vout.n455 76.4201
R623 vout.n274 vout.n273 75.8248
R624 vout.n268 vout.n267 75.8248
R625 vout.n285 vout.n284 75.8248
R626 vout.n263 vout.n262 75.8248
R627 vout.n258 vout.n257 75.8248
R628 vout.n302 vout.n301 75.8248
R629 vout.n252 vout.n251 75.8248
R630 vout.n247 vout.n246 75.8248
R631 vout.n318 vout.n317 75.8248
R632 vout.n242 vout.n241 75.8248
R633 vout.n237 vout.n236 75.8248
R634 vout.n234 vout.n233 75.8248
R635 vout.n227 vout.n226 75.8248
R636 vout.n344 vout.n343 75.8248
R637 vout.n222 vout.n221 75.8248
R638 vout.n217 vout.n216 75.8248
R639 vout.n209 vout.n208 75.8248
R640 vout.n366 vout.n365 75.8248
R641 vout.n206 vout.n205 75.8248
R642 vout.n201 vout.n200 75.8248
R643 vout.n383 vout.n382 75.8248
R644 vout.n196 vout.n195 75.8248
R645 vout.n191 vout.n190 75.8248
R646 vout.n188 vout.n187 75.8248
R647 vout.n405 vout.n404 75.8248
R648 vout.n180 vout.n179 75.8248
R649 vout.n175 vout.n174 75.8248
R650 vout.n421 vout.n420 75.8248
R651 vout.n170 vout.n169 75.8248
R652 vout.n432 vout.n431 75.8248
R653 vout.n165 vout.n164 75.8248
R654 vout.n440 vout.n439 75.8248
R655 vout.n445 vout.n444 75.8248
R656 vout.n450 vout.n449 75.8248
R657 vout.n454 vout.n453 75.8248
R658 vout.n457 vout.n456 75.8248
R659 vout.n80 vout.n79 57.8105
R660 vout.n18 vout.t95 20.6431
R661 vout.n18 vout.t73 19.9282
R662 vout.n66 vout.n64 16.7764
R663 vout.n61 vout.n59 16.7764
R664 vout.n56 vout.n54 16.7764
R665 vout.n51 vout.n49 16.7764
R666 vout.n46 vout.n44 16.7764
R667 vout.n136 vout.n134 16.7764
R668 vout.n552 vout.n550 16.7764
R669 vout.n549 vout.n547 16.7764
R670 vout.n128 vout.n126 16.7764
R671 vout.n123 vout.n121 16.7764
R672 vout.n118 vout.n116 16.7764
R673 vout.n114 vout.n112 16.7764
R674 vout.n109 vout.n107 16.7764
R675 vout.n103 vout.n101 16.7764
R676 vout.n98 vout.n96 16.7764
R677 vout.n94 vout.n92 16.7764
R678 vout.n89 vout.n87 16.7764
R679 vout.n84 vout.n82 16.7764
R680 vout.n77 vout.n75 16.7764
R681 vout.n482 vout.n480 16.7764
R682 vout.n159 vout.n157 16.7764
R683 vout.n154 vout.n152 16.7764
R684 vout.n150 vout.n148 16.7764
R685 vout.n145 vout.n143 16.7764
R686 vout.n140 vout.n138 16.7764
R687 vout.n133 vout.n131 16.7764
R688 vout.n496 vout.n494 16.7764
R689 vout.n500 vout.n498 16.7764
R690 vout.n492 vout.n490 16.7764
R691 vout.n487 vout.n485 16.7764
R692 vout.n7 vout.n5 16.7764
R693 vout.n12 vout.n10 16.7764
R694 vout.n17 vout.n15 16.7764
R695 vout.n42 vout.n40 16.7764
R696 vout.n34 vout.n32 16.7764
R697 vout.n63 vout.n62 16.6901
R698 vout.n79 vout.n78 16.5309
R699 vout.n68 vout.n67 16.0615
R700 vout.n66 vout.n65 16.0615
R701 vout.n61 vout.n60 16.0615
R702 vout.n56 vout.n55 16.0615
R703 vout.n51 vout.n50 16.0615
R704 vout.n46 vout.n45 16.0615
R705 vout.n136 vout.n135 16.0615
R706 vout.n552 vout.n551 16.0615
R707 vout.n549 vout.n548 16.0615
R708 vout.n128 vout.n127 16.0615
R709 vout.n123 vout.n122 16.0615
R710 vout.n118 vout.n117 16.0615
R711 vout.n114 vout.n113 16.0615
R712 vout.n109 vout.n108 16.0615
R713 vout.n103 vout.n102 16.0615
R714 vout.n98 vout.n97 16.0615
R715 vout.n94 vout.n93 16.0615
R716 vout.n89 vout.n88 16.0615
R717 vout.n84 vout.n83 16.0615
R718 vout.n74 vout.n73 16.0615
R719 vout.n77 vout.n76 16.0615
R720 vout.n482 vout.n481 16.0615
R721 vout.n159 vout.n158 16.0615
R722 vout.n154 vout.n153 16.0615
R723 vout.n150 vout.n149 16.0615
R724 vout.n145 vout.n144 16.0615
R725 vout.n140 vout.n139 16.0615
R726 vout.n133 vout.n132 16.0615
R727 vout.n496 vout.n495 16.0615
R728 vout.n500 vout.n499 16.0615
R729 vout.n492 vout.n491 16.0615
R730 vout.n487 vout.n486 16.0615
R731 vout.n7 vout.n6 16.0615
R732 vout.n12 vout.n11 16.0615
R733 vout.n17 vout.n16 16.0615
R734 vout.n42 vout.n41 16.0615
R735 vout.n34 vout.n33 16.0615
R736 vout.n272 vout.t46 9.52217
R737 vout.n272 vout.t293 9.52217
R738 vout.n273 vout.t225 9.52217
R739 vout.n273 vout.t19 9.52217
R740 vout.n266 vout.t8 9.52217
R741 vout.n266 vout.t50 9.52217
R742 vout.n267 vout.t38 9.52217
R743 vout.n267 vout.t285 9.52217
R744 vout.n283 vout.t231 9.52217
R745 vout.n283 vout.t213 9.52217
R746 vout.n284 vout.t271 9.52217
R747 vout.n284 vout.t7 9.52217
R748 vout.n261 vout.t274 9.52217
R749 vout.n261 vout.t56 9.52217
R750 vout.n262 vout.t45 9.52217
R751 vout.n262 vout.t280 9.52217
R752 vout.n256 vout.t248 9.52217
R753 vout.n256 vout.t238 9.52217
R754 vout.n257 vout.t1 9.52217
R755 vout.n257 vout.t41 9.52217
R756 vout.n300 vout.t258 9.52217
R757 vout.n300 vout.t289 9.52217
R758 vout.n301 vout.t272 9.52217
R759 vout.n301 vout.t278 9.52217
R760 vout.n250 vout.t49 9.52217
R761 vout.n250 vout.t228 9.52217
R762 vout.n251 vout.t10 9.52217
R763 vout.n251 vout.t282 9.52217
R764 vout.n245 vout.t29 9.52217
R765 vout.n245 vout.t51 9.52217
R766 vout.n246 vout.t222 9.52217
R767 vout.n246 vout.t5 9.52217
R768 vout.n316 vout.t260 9.52217
R769 vout.n316 vout.t18 9.52217
R770 vout.n317 vout.t275 9.52217
R771 vout.n317 vout.t234 9.52217
R772 vout.n240 vout.t37 9.52217
R773 vout.n240 vout.t277 9.52217
R774 vout.n241 vout.t212 9.52217
R775 vout.n241 vout.t240 9.52217
R776 vout.n235 vout.t4 9.52217
R777 vout.n235 vout.t47 9.52217
R778 vout.n236 vout.t233 9.52217
R779 vout.n236 vout.t276 9.52217
R780 vout.n232 vout.t58 9.52217
R781 vout.n232 vout.t288 9.52217
R782 vout.n233 vout.t254 9.52217
R783 vout.n233 vout.t9 9.52217
R784 vout.n225 vout.t14 9.52217
R785 vout.n225 vout.t230 9.52217
R786 vout.n226 vout.t16 9.52217
R787 vout.n226 vout.t42 9.52217
R788 vout.n342 vout.t31 9.52217
R789 vout.n342 vout.t235 9.52217
R790 vout.n343 vout.t244 9.52217
R791 vout.n343 vout.t237 9.52217
R792 vout.n220 vout.t0 9.52217
R793 vout.n220 vout.t251 9.52217
R794 vout.n221 vout.t256 9.52217
R795 vout.n221 vout.t35 9.52217
R796 vout.n215 vout.t291 9.52217
R797 vout.n215 vout.t12 9.52217
R798 vout.n216 vout.t30 9.52217
R799 vout.n216 vout.t287 9.52217
R800 vout.n207 vout.t24 9.52217
R801 vout.n207 vout.t53 9.52217
R802 vout.n208 vout.t290 9.52217
R803 vout.n208 vout.t215 9.52217
R804 vout.n364 vout.t22 9.52217
R805 vout.n364 vout.t2 9.52217
R806 vout.n365 vout.t273 9.52217
R807 vout.n365 vout.t229 9.52217
R808 vout.n204 vout.t267 9.52217
R809 vout.n204 vout.t252 9.52217
R810 vout.n205 vout.t257 9.52217
R811 vout.n205 vout.t224 9.52217
R812 vout.n199 vout.t52 9.52217
R813 vout.n199 vout.t223 9.52217
R814 vout.n200 vout.t39 9.52217
R815 vout.n200 vout.t48 9.52217
R816 vout.n381 vout.t209 9.52217
R817 vout.n381 vout.t284 9.52217
R818 vout.n382 vout.t54 9.52217
R819 vout.n382 vout.t269 9.52217
R820 vout.n194 vout.t243 9.52217
R821 vout.n194 vout.t34 9.52217
R822 vout.n195 vout.t263 9.52217
R823 vout.n195 vout.t296 9.52217
R824 vout.n189 vout.t295 9.52217
R825 vout.n189 vout.t13 9.52217
R826 vout.n190 vout.t218 9.52217
R827 vout.n190 vout.t247 9.52217
R828 vout.n186 vout.t286 9.52217
R829 vout.n186 vout.t40 9.52217
R830 vout.n187 vout.t239 9.52217
R831 vout.n187 vout.t25 9.52217
R832 vout.n403 vout.t32 9.52217
R833 vout.n403 vout.t279 9.52217
R834 vout.n404 vout.t15 9.52217
R835 vout.n404 vout.t20 9.52217
R836 vout.n178 vout.t227 9.52217
R837 vout.n178 vout.t55 9.52217
R838 vout.n179 vout.t232 9.52217
R839 vout.n179 vout.t262 9.52217
R840 vout.n173 vout.t33 9.52217
R841 vout.n173 vout.t216 9.52217
R842 vout.n174 vout.t294 9.52217
R843 vout.n174 vout.t220 9.52217
R844 vout.n419 vout.t250 9.52217
R845 vout.n419 vout.t57 9.52217
R846 vout.n420 vout.t255 9.52217
R847 vout.n420 vout.t242 9.52217
R848 vout.n168 vout.t23 9.52217
R849 vout.n168 vout.t292 9.52217
R850 vout.n169 vout.t249 9.52217
R851 vout.n169 vout.t253 9.52217
R852 vout.n430 vout.t27 9.52217
R853 vout.n430 vout.t217 9.52217
R854 vout.n431 vout.t11 9.52217
R855 vout.n431 vout.t236 9.52217
R856 vout.n163 vout.t266 9.52217
R857 vout.n163 vout.t298 9.52217
R858 vout.n164 vout.t3 9.52217
R859 vout.n164 vout.t299 9.52217
R860 vout.n438 vout.t210 9.52217
R861 vout.n438 vout.t270 9.52217
R862 vout.n439 vout.t265 9.52217
R863 vout.n439 vout.t281 9.52217
R864 vout.n443 vout.t28 9.52217
R865 vout.n443 vout.t36 9.52217
R866 vout.n444 vout.t221 9.52217
R867 vout.n444 vout.t6 9.52217
R868 vout.n448 vout.t259 9.52217
R869 vout.n448 vout.t264 9.52217
R870 vout.n449 vout.t219 9.52217
R871 vout.n449 vout.t43 9.52217
R872 vout.n452 vout.t17 9.52217
R873 vout.n452 vout.t26 9.52217
R874 vout.n453 vout.t21 9.52217
R875 vout.n453 vout.t211 9.52217
R876 vout.n455 vout.t245 9.52217
R877 vout.n455 vout.t44 9.52217
R878 vout.n456 vout.t268 9.52217
R879 vout.n456 vout.t261 9.52217
R880 vout.n62 vout.t84 3.86717
R881 vout.n62 vout.t180 3.86717
R882 vout.n67 vout.t197 3.86717
R883 vout.n67 vout.t144 3.86717
R884 vout.n64 vout.t125 3.86717
R885 vout.n64 vout.t99 3.86717
R886 vout.n65 vout.t135 3.86717
R887 vout.n65 vout.t134 3.86717
R888 vout.n59 vout.t88 3.86717
R889 vout.n59 vout.t193 3.86717
R890 vout.n60 vout.t124 3.86717
R891 vout.n60 vout.t115 3.86717
R892 vout.n54 vout.t89 3.86717
R893 vout.n54 vout.t80 3.86717
R894 vout.n55 vout.t139 3.86717
R895 vout.n55 vout.t136 3.86717
R896 vout.n49 vout.t154 3.86717
R897 vout.n49 vout.t151 3.86717
R898 vout.n50 vout.t165 3.86717
R899 vout.n50 vout.t202 3.86717
R900 vout.n44 vout.t174 3.86717
R901 vout.n44 vout.t143 3.86717
R902 vout.n45 vout.t190 3.86717
R903 vout.n45 vout.t113 3.86717
R904 vout.n134 vout.t170 3.86717
R905 vout.n134 vout.t106 3.86717
R906 vout.n135 vout.t82 3.86717
R907 vout.n135 vout.t149 3.86717
R908 vout.n550 vout.t107 3.86717
R909 vout.n550 vout.t60 3.86717
R910 vout.n551 vout.t192 3.86717
R911 vout.n551 vout.t86 3.86717
R912 vout.n547 vout.t205 3.86717
R913 vout.n547 vout.t132 3.86717
R914 vout.n548 vout.t127 3.86717
R915 vout.n548 vout.t116 3.86717
R916 vout.n126 vout.t182 3.86717
R917 vout.n126 vout.t110 3.86717
R918 vout.n127 vout.t196 3.86717
R919 vout.n127 vout.t158 3.86717
R920 vout.n121 vout.t138 3.86717
R921 vout.n121 vout.t186 3.86717
R922 vout.n122 vout.t163 3.86717
R923 vout.n122 vout.t65 3.86717
R924 vout.n116 vout.t130 3.86717
R925 vout.n116 vout.t145 3.86717
R926 vout.n117 vout.t100 3.86717
R927 vout.n117 vout.t108 3.86717
R928 vout.n112 vout.t155 3.86717
R929 vout.n112 vout.t183 3.86717
R930 vout.n113 vout.t198 3.86717
R931 vout.n113 vout.t176 3.86717
R932 vout.n107 vout.t75 3.86717
R933 vout.n107 vout.t206 3.86717
R934 vout.n108 vout.t61 3.86717
R935 vout.n108 vout.t152 3.86717
R936 vout.n101 vout.t167 3.86717
R937 vout.n101 vout.t123 3.86717
R938 vout.n102 vout.t156 3.86717
R939 vout.n102 vout.t162 3.86717
R940 vout.n96 vout.t191 3.86717
R941 vout.n96 vout.t200 3.86717
R942 vout.n97 vout.t97 3.86717
R943 vout.n97 vout.t87 3.86717
R944 vout.n92 vout.t140 3.86717
R945 vout.n92 vout.t90 3.86717
R946 vout.n93 vout.t150 3.86717
R947 vout.n93 vout.t78 3.86717
R948 vout.n87 vout.t85 3.86717
R949 vout.n87 vout.t194 3.86717
R950 vout.n88 vout.t166 3.86717
R951 vout.n88 vout.t201 3.86717
R952 vout.n82 vout.t104 3.86717
R953 vout.n82 vout.t147 3.86717
R954 vout.n83 vout.t70 3.86717
R955 vout.n83 vout.t168 3.86717
R956 vout.n78 vout.t63 3.86717
R957 vout.n78 vout.t128 3.86717
R958 vout.n73 vout.t102 3.86717
R959 vout.n73 vout.t177 3.86717
R960 vout.n75 vout.t153 3.86717
R961 vout.n75 vout.t169 3.86717
R962 vout.n76 vout.t172 3.86717
R963 vout.n76 vout.t142 3.86717
R964 vout.n480 vout.t179 3.86717
R965 vout.n480 vout.t114 3.86717
R966 vout.n481 vout.t83 3.86717
R967 vout.n481 vout.t69 3.86717
R968 vout.n157 vout.t199 3.86717
R969 vout.n157 vout.t178 3.86717
R970 vout.n158 vout.t103 3.86717
R971 vout.n158 vout.t171 3.86717
R972 vout.n152 vout.t129 3.86717
R973 vout.n152 vout.t109 3.86717
R974 vout.n153 vout.t120 3.86717
R975 vout.n153 vout.t118 3.86717
R976 vout.n148 vout.t159 3.86717
R977 vout.n148 vout.t173 3.86717
R978 vout.n149 vout.t112 3.86717
R979 vout.n149 vout.t72 3.86717
R980 vout.n143 vout.t96 3.86717
R981 vout.n143 vout.t126 3.86717
R982 vout.n144 vout.t164 3.86717
R983 vout.n144 vout.t207 3.86717
R984 vout.n138 vout.t141 3.86717
R985 vout.n138 vout.t76 3.86717
R986 vout.n139 vout.t91 3.86717
R987 vout.n139 vout.t117 3.86717
R988 vout.n131 vout.t208 3.86717
R989 vout.n131 vout.t62 3.86717
R990 vout.n132 vout.t93 3.86717
R991 vout.n132 vout.t161 3.86717
R992 vout.n494 vout.t204 3.86717
R993 vout.n494 vout.t98 3.86717
R994 vout.n495 vout.t187 3.86717
R995 vout.n495 vout.t160 3.86717
R996 vout.n498 vout.t157 3.86717
R997 vout.n498 vout.t81 3.86717
R998 vout.n499 vout.t189 3.86717
R999 vout.n499 vout.t184 3.86717
R1000 vout.n490 vout.t101 3.86717
R1001 vout.n490 vout.t122 3.86717
R1002 vout.n491 vout.t137 3.86717
R1003 vout.n491 vout.t148 3.86717
R1004 vout.n485 vout.t94 3.86717
R1005 vout.n485 vout.t188 3.86717
R1006 vout.n486 vout.t92 3.86717
R1007 vout.n486 vout.t79 3.86717
R1008 vout.n5 vout.t64 3.86717
R1009 vout.n5 vout.t59 3.86717
R1010 vout.n6 vout.t71 3.86717
R1011 vout.n6 vout.t131 3.86717
R1012 vout.n10 vout.t119 3.86717
R1013 vout.n10 vout.t121 3.86717
R1014 vout.n11 vout.t67 3.86717
R1015 vout.n11 vout.t105 3.86717
R1016 vout.n15 vout.t185 3.86717
R1017 vout.n15 vout.t66 3.86717
R1018 vout.n16 vout.t146 3.86717
R1019 vout.n16 vout.t133 3.86717
R1020 vout.n40 vout.t68 3.86717
R1021 vout.n40 vout.t111 3.86717
R1022 vout.n41 vout.t203 3.86717
R1023 vout.n41 vout.t74 3.86717
R1024 vout.n32 vout.t77 3.86717
R1025 vout.n32 vout.t195 3.86717
R1026 vout.n33 vout.t181 3.86717
R1027 vout.n33 vout.t175 3.86717
R1028 vout.n368 vout.n367 3.4105
R1029 vout.n371 vout.n370 3.4105
R1030 vout.n70 vout.n63 2.75235
R1031 vout.n369 vout.n368 1.70282
R1032 vout.n373 vout.n212 1.70282
R1033 vout.n360 vout.n211 1.70282
R1034 vout.n372 vout.n213 1.70282
R1035 vout.n371 vout.n361 1.70282
R1036 vout.n80 vout.n77 1.69312
R1037 vout.n399 vout.n184 1.15193
R1038 vout.n335 vout.n334 1.14771
R1039 vout.n396 vout.n185 1.13717
R1040 vout.n395 vout.n394 1.13717
R1041 vout.n393 vout.n392 1.13717
R1042 vout.n391 vout.n193 1.13717
R1043 vout.n389 vout.n388 1.13717
R1044 vout.n387 vout.n197 1.13717
R1045 vout.n386 vout.n385 1.13717
R1046 vout.n380 vout.n198 1.13717
R1047 vout.n379 vout.n378 1.13717
R1048 vout.n377 vout.n376 1.13717
R1049 vout.n375 vout.n203 1.13717
R1050 vout.n359 vout.n358 1.13717
R1051 vout.n357 vout.n214 1.13717
R1052 vout.n356 vout.n355 1.13717
R1053 vout.n354 vout.n353 1.13717
R1054 vout.n352 vout.n219 1.13717
R1055 vout.n350 vout.n349 1.13717
R1056 vout.n348 vout.n223 1.13717
R1057 vout.n347 vout.n346 1.13717
R1058 vout.n341 vout.n224 1.13717
R1059 vout.n340 vout.n339 1.13717
R1060 vout.n338 vout.n337 1.13717
R1061 vout.n336 vout.n229 1.13717
R1062 vout.n331 vout.n231 1.13717
R1063 vout.n330 vout.n329 1.13717
R1064 vout.n328 vout.n327 1.13717
R1065 vout.n326 vout.n239 1.13717
R1066 vout.n324 vout.n323 1.13717
R1067 vout.n322 vout.n243 1.13717
R1068 vout.n321 vout.n320 1.13717
R1069 vout.n315 vout.n244 1.13717
R1070 vout.n314 vout.n313 1.13717
R1071 vout.n312 vout.n311 1.13717
R1072 vout.n310 vout.n249 1.13717
R1073 vout.n308 vout.n307 1.13717
R1074 vout.n306 vout.n253 1.13717
R1075 vout.n305 vout.n304 1.13717
R1076 vout.n298 vout.n254 1.13717
R1077 vout.n297 vout.n296 1.13717
R1078 vout.n295 vout.n294 1.13717
R1079 vout.n293 vout.n260 1.13717
R1080 vout.n291 vout.n290 1.13717
R1081 vout.n289 vout.n264 1.13717
R1082 vout.n288 vout.n287 1.13717
R1083 vout.n282 vout.n265 1.13717
R1084 vout.n280 vout.n279 1.13717
R1085 vout.n278 vout.n269 1.13717
R1086 vout.n277 vout.n276 1.13717
R1087 vout.n429 vout.n167 1.13717
R1088 vout.n427 vout.n426 1.13717
R1089 vout.n425 vout.n171 1.13717
R1090 vout.n424 vout.n423 1.13717
R1091 vout.n418 vout.n172 1.13717
R1092 vout.n417 vout.n416 1.13717
R1093 vout.n415 vout.n414 1.13717
R1094 vout.n413 vout.n177 1.13717
R1095 vout.n411 vout.n410 1.13717
R1096 vout.n409 vout.n181 1.13717
R1097 vout.n408 vout.n407 1.13717
R1098 vout.n402 vout.n182 1.13717
R1099 vout.n401 vout.n400 1.13717
R1100 vout.n460 vout.n447 1.13717
R1101 vout.n462 vout.n461 1.13717
R1102 vout.n463 vout.n446 1.13717
R1103 vout.n465 vout.n464 1.13717
R1104 vout.n467 vout.n442 1.13717
R1105 vout.n469 vout.n468 1.13717
R1106 vout.n471 vout.n470 1.13717
R1107 vout.n472 vout.n437 1.13717
R1108 vout.n474 vout.n473 1.13717
R1109 vout.n476 vout.n475 1.13717
R1110 vout.n436 vout.n162 1.13717
R1111 vout.n435 vout.n434 1.13717
R1112 vout.n605 vout.n71 1.13717
R1113 vout.n503 vout.n502 1.13717
R1114 vout.n504 vout.n493 1.13717
R1115 vout.n506 vout.n505 1.13717
R1116 vout.n508 vout.n489 1.13717
R1117 vout.n510 vout.n509 1.13717
R1118 vout.n512 vout.n511 1.13717
R1119 vout.n513 vout.n484 1.13717
R1120 vout.n515 vout.n514 1.13717
R1121 vout.n517 vout.n516 1.13717
R1122 vout.n519 vout.n161 1.13717
R1123 vout.n521 vout.n520 1.13717
R1124 vout.n523 vout.n522 1.13717
R1125 vout.n524 vout.n156 1.13717
R1126 vout.n526 vout.n525 1.13717
R1127 vout.n528 vout.n527 1.13717
R1128 vout.n529 vout.n147 1.13717
R1129 vout.n531 vout.n530 1.13717
R1130 vout.n532 vout.n146 1.13717
R1131 vout.n534 vout.n533 1.13717
R1132 vout.n535 vout.n142 1.13717
R1133 vout.n538 vout.n537 1.13717
R1134 vout.n539 vout.n141 1.13717
R1135 vout.n541 vout.n540 1.13717
R1136 vout.n543 vout.n130 1.13717
R1137 vout.n545 vout.n544 1.13717
R1138 vout.n554 vout.n546 1.13717
R1139 vout.n556 vout.n555 1.13717
R1140 vout.n558 vout.n557 1.13717
R1141 vout.n559 vout.n125 1.13717
R1142 vout.n561 vout.n560 1.13717
R1143 vout.n563 vout.n562 1.13717
R1144 vout.n564 vout.n120 1.13717
R1145 vout.n566 vout.n565 1.13717
R1146 vout.n568 vout.n567 1.13717
R1147 vout.n569 vout.n111 1.13717
R1148 vout.n571 vout.n570 1.13717
R1149 vout.n572 vout.n110 1.13717
R1150 vout.n574 vout.n573 1.13717
R1151 vout.n575 vout.n105 1.13717
R1152 vout.n578 vout.n577 1.13717
R1153 vout.n579 vout.n104 1.13717
R1154 vout.n581 vout.n580 1.13717
R1155 vout.n583 vout.n100 1.13717
R1156 vout.n585 vout.n584 1.13717
R1157 vout.n587 vout.n586 1.13717
R1158 vout.n588 vout.n91 1.13717
R1159 vout.n590 vout.n589 1.13717
R1160 vout.n591 vout.n90 1.13717
R1161 vout.n593 vout.n592 1.13717
R1162 vout.n594 vout.n86 1.13717
R1163 vout.n597 vout.n596 1.13717
R1164 vout.n598 vout.n85 1.13717
R1165 vout.n600 vout.n599 1.13717
R1166 vout.n602 vout.n72 1.13717
R1167 vout.n604 vout.n603 1.13717
R1168 vout.n607 vout.n606 1.13717
R1169 vout.n608 vout.n58 1.13717
R1170 vout.n611 vout.n610 1.13717
R1171 vout.n612 vout.n57 1.13717
R1172 vout.n614 vout.n613 1.13717
R1173 vout.n616 vout.n53 1.13717
R1174 vout.n618 vout.n617 1.13717
R1175 vout.n620 vout.n619 1.13717
R1176 vout.n621 vout.n48 1.13717
R1177 vout.n623 vout.n622 1.13717
R1178 vout.n625 vout.n624 1.13717
R1179 vout.n626 vout.n39 1.13717
R1180 vout.n628 vout.n627 1.13717
R1181 vout.n37 vout.n36 1.13717
R1182 vout.n31 vout.n4 1.13717
R1183 vout.n30 vout.n29 1.13717
R1184 vout.n28 vout.n27 1.13717
R1185 vout.n26 vout.n9 1.13717
R1186 vout.n25 vout.n24 1.13717
R1187 vout.n23 vout.n22 1.13717
R1188 vout.n21 vout.n14 1.13717
R1189 vout.n629 vout.n3 1.13717
R1190 vout.n631 vout.n630 1.13717
R1191 vout.n38 vout.n2 1.13717
R1192 vout.n69 vout.n66 0.709343
R1193 vout.n69 vout.n68 0.704661
R1194 vout.n137 vout.n136 0.66979
R1195 vout.n553 vout.n552 0.66979
R1196 vout.n333 vout.n332 0.572856
R1197 vout.n398 vout.n397 0.571952
R1198 vout.n19 vout.n18 0.491863
R1199 vout.n497 vout.n496 0.489753
R1200 vout.n81 vout.n74 0.479273
R1201 vout.n609 vout.n61 0.472974
R1202 vout.n615 vout.n56 0.472974
R1203 vout.n52 vout.n51 0.472974
R1204 vout.n47 vout.n46 0.472974
R1205 vout.n553 vout.n549 0.472974
R1206 vout.n129 vout.n128 0.472974
R1207 vout.n124 vout.n123 0.472974
R1208 vout.n119 vout.n118 0.472974
R1209 vout.n115 vout.n114 0.472974
R1210 vout.n576 vout.n109 0.472974
R1211 vout.n582 vout.n103 0.472974
R1212 vout.n99 vout.n98 0.472974
R1213 vout.n95 vout.n94 0.472974
R1214 vout.n595 vout.n89 0.472974
R1215 vout.n601 vout.n84 0.472974
R1216 vout.n483 vout.n482 0.472974
R1217 vout.n160 vout.n159 0.472974
R1218 vout.n155 vout.n154 0.472974
R1219 vout.n151 vout.n150 0.472974
R1220 vout.n536 vout.n145 0.472974
R1221 vout.n542 vout.n140 0.472974
R1222 vout.n137 vout.n133 0.472974
R1223 vout.n501 vout.n500 0.472974
R1224 vout.n507 vout.n492 0.472974
R1225 vout.n488 vout.n487 0.472974
R1226 vout.n8 vout.n7 0.472974
R1227 vout.n13 vout.n12 0.472974
R1228 vout.n20 vout.n17 0.472974
R1229 vout.n43 vout.n42 0.472974
R1230 vout.n35 vout.n34 0.472974
R1231 vout.n458 vout.n457 0.45495
R1232 vout.n271 vout.n270 0.449638
R1233 vout.n368 vout.n366 0.445531
R1234 vout.n275 vout.n274 0.439167
R1235 vout.n281 vout.n268 0.439167
R1236 vout.n286 vout.n285 0.439167
R1237 vout.n292 vout.n263 0.439167
R1238 vout.n259 vout.n258 0.439167
R1239 vout.n303 vout.n302 0.439167
R1240 vout.n309 vout.n252 0.439167
R1241 vout.n248 vout.n247 0.439167
R1242 vout.n319 vout.n318 0.439167
R1243 vout.n325 vout.n242 0.439167
R1244 vout.n238 vout.n237 0.439167
R1245 vout.n332 vout.n234 0.439167
R1246 vout.n335 vout.n230 0.439167
R1247 vout.n228 vout.n227 0.439167
R1248 vout.n345 vout.n344 0.439167
R1249 vout.n351 vout.n222 0.439167
R1250 vout.n218 vout.n217 0.439167
R1251 vout.n210 vout.n209 0.439167
R1252 vout.n374 vout.n206 0.439167
R1253 vout.n202 vout.n201 0.439167
R1254 vout.n384 vout.n383 0.439167
R1255 vout.n390 vout.n196 0.439167
R1256 vout.n192 vout.n191 0.439167
R1257 vout.n397 vout.n188 0.439167
R1258 vout.n184 vout.n183 0.439167
R1259 vout.n406 vout.n405 0.439167
R1260 vout.n412 vout.n180 0.439167
R1261 vout.n176 vout.n175 0.439167
R1262 vout.n422 vout.n421 0.439167
R1263 vout.n428 vout.n170 0.439167
R1264 vout.n433 vout.n432 0.439167
R1265 vout.n166 vout.n165 0.439167
R1266 vout.n441 vout.n440 0.439167
R1267 vout.n466 vout.n445 0.439167
R1268 vout.n451 vout.n450 0.439167
R1269 vout.n459 vout.n454 0.439167
R1270 vout.n635 vout.n0 0.40423
R1271 vout.n277 vout.n271 0.395966
R1272 vout.n68 vout.n63 0.342089
R1273 vout.n458 vout.n447 0.30251
R1274 vout vout.n634 0.296012
R1275 vout.n79 vout.n74 0.255553
R1276 vout.n503 vout.n497 0.249543
R1277 vout.n19 vout.n14 0.248362
R1278 vout.n334 vout.n333 0.143382
R1279 vout.n363 vout.n362 0.141125
R1280 vout.n479 vout.n478 0.141125
R1281 vout.n399 vout.n398 0.140689
R1282 vout.n634 vout.n1 0.139783
R1283 vout.n605 vout.n604 0.135258
R1284 vout.n546 vout.n545 0.132565
R1285 vout.n0 vout 0.0623497
R1286 vout.n371 vout.n363 0.0580834
R1287 vout.n362 vout.n106 0.0522084
R1288 vout.n518 vout.n479 0.0522084
R1289 vout.n478 vout.n477 0.0517188
R1290 vout.n633 vout.n632 0.051474
R1291 vout.n299 vout.n255 0.0491168
R1292 vout vout.n635 0.0475
R1293 vout.n501 vout.n497 0.0302612
R1294 vout.n20 vout.n19 0.0279613
R1295 vout.n275 vout.n271 0.0273537
R1296 vout.n635 vout 0.024
R1297 vout.n459 vout.n458 0.0226014
R1298 vout.n603 vout.n81 0.021891
R1299 vout.n333 vout.n231 0.0207578
R1300 vout.n398 vout.n185 0.0207578
R1301 vout.n627 vout.n626 0.0161667
R1302 vout.n626 vout.n625 0.0161667
R1303 vout.n622 vout.n621 0.0161667
R1304 vout.n621 vout.n620 0.0161667
R1305 vout.n617 vout.n616 0.0161667
R1306 vout.n614 vout.n57 0.0161667
R1307 vout.n610 vout.n57 0.0161667
R1308 vout.n608 vout.n607 0.0161667
R1309 vout.n607 vout.n71 0.0161667
R1310 vout.n276 vout.n269 0.0161667
R1311 vout.n280 vout.n269 0.0161667
R1312 vout.n287 vout.n282 0.0161667
R1313 vout.n291 vout.n264 0.0161667
R1314 vout.n294 vout.n293 0.0161667
R1315 vout.n298 vout.n297 0.0161667
R1316 vout.n308 vout.n253 0.0161667
R1317 vout.n311 vout.n310 0.0161667
R1318 vout.n315 vout.n314 0.0161667
R1319 vout.n320 vout.n315 0.0161667
R1320 vout.n324 vout.n243 0.0161667
R1321 vout.n327 vout.n326 0.0161667
R1322 vout.n331 vout.n330 0.0161667
R1323 vout.n337 vout.n336 0.0161667
R1324 vout.n341 vout.n340 0.0161667
R1325 vout.n346 vout.n341 0.0161667
R1326 vout.n350 vout.n223 0.0161667
R1327 vout.n353 vout.n352 0.0161667
R1328 vout.n357 vout.n356 0.0161667
R1329 vout.n358 vout.n357 0.0161667
R1330 vout.n574 vout.n110 0.0161667
R1331 vout.n570 vout.n569 0.0161667
R1332 vout.n569 vout.n568 0.0161667
R1333 vout.n565 vout.n564 0.0161667
R1334 vout.n564 vout.n563 0.0161667
R1335 vout.n560 vout.n559 0.0161667
R1336 vout.n559 vout.n558 0.0161667
R1337 vout.n555 vout.n554 0.0161667
R1338 vout.n603 vout.n602 0.0161667
R1339 vout.n600 vout.n85 0.0161667
R1340 vout.n596 vout.n85 0.0161667
R1341 vout.n594 vout.n593 0.0161667
R1342 vout.n593 vout.n90 0.0161667
R1343 vout.n589 vout.n588 0.0161667
R1344 vout.n588 vout.n587 0.0161667
R1345 vout.n584 vout.n583 0.0161667
R1346 vout.n581 vout.n104 0.0161667
R1347 vout.n376 vout.n375 0.0161667
R1348 vout.n380 vout.n379 0.0161667
R1349 vout.n385 vout.n380 0.0161667
R1350 vout.n389 vout.n197 0.0161667
R1351 vout.n392 vout.n391 0.0161667
R1352 vout.n396 vout.n395 0.0161667
R1353 vout.n402 vout.n401 0.0161667
R1354 vout.n407 vout.n402 0.0161667
R1355 vout.n411 vout.n181 0.0161667
R1356 vout.n414 vout.n413 0.0161667
R1357 vout.n418 vout.n417 0.0161667
R1358 vout.n423 vout.n418 0.0161667
R1359 vout.n427 vout.n171 0.0161667
R1360 vout.n434 vout.n429 0.0161667
R1361 vout.n473 vout.n472 0.0161667
R1362 vout.n472 vout.n471 0.0161667
R1363 vout.n468 vout.n467 0.0161667
R1364 vout.n465 vout.n446 0.0161667
R1365 vout.n461 vout.n460 0.0161667
R1366 vout.n544 vout.n543 0.0161667
R1367 vout.n541 vout.n141 0.0161667
R1368 vout.n537 vout.n141 0.0161667
R1369 vout.n535 vout.n534 0.0161667
R1370 vout.n534 vout.n146 0.0161667
R1371 vout.n530 vout.n529 0.0161667
R1372 vout.n529 vout.n528 0.0161667
R1373 vout.n525 vout.n524 0.0161667
R1374 vout.n524 vout.n523 0.0161667
R1375 vout.n520 vout.n519 0.0161667
R1376 vout.n514 vout.n513 0.0161667
R1377 vout.n513 vout.n512 0.0161667
R1378 vout.n509 vout.n508 0.0161667
R1379 vout.n506 vout.n493 0.0161667
R1380 vout.n502 vout.n493 0.0161667
R1381 vout.n22 vout.n21 0.0161667
R1382 vout.n26 vout.n25 0.0161667
R1383 vout.n27 vout.n26 0.0161667
R1384 vout.n31 vout.n30 0.0161667
R1385 vout.n36 vout.n31 0.0161667
R1386 vout.n575 vout.n574 0.0161667
R1387 vout.n584 vout.n99 0.016016
R1388 vout.n631 vout.n3 0.0158711
R1389 vout.n616 vout.n615 0.0158654
R1390 vout.n422 vout.n171 0.0158654
R1391 vout.n509 vout.n488 0.0158654
R1392 vout.n294 vout.n259 0.0155641
R1393 vout.n319 vout.n243 0.0155641
R1394 vout.n337 vout.n228 0.0152628
R1395 vout.n543 vout.n542 0.0152628
R1396 vout.n21 vout.n20 0.0152628
R1397 vout.n554 vout.n553 0.0151122
R1398 vout.n477 vout.n476 0.0151122
R1399 vout.n518 vout.n517 0.0151122
R1400 vout.n299 vout.n298 0.0148109
R1401 vout.n555 vout.n129 0.0148109
R1402 vout.n384 vout.n197 0.0146603
R1403 vout.n397 vout.n396 0.0146603
R1404 vout.n468 vout.n441 0.0146603
R1405 vout.n460 vout.n459 0.0146603
R1406 vout.n544 vout.n137 0.0146603
R1407 vout.n22 vout.n13 0.0146603
R1408 vout.n632 vout.n2 0.0145409
R1409 vout.n617 vout.n52 0.0140577
R1410 vout.n508 vout.n507 0.0140577
R1411 vout.n583 vout.n582 0.0139071
R1412 vout.n282 vout.n281 0.0137564
R1413 vout.n332 vout.n331 0.0137564
R1414 vout.n589 vout.n95 0.0136058
R1415 vout.n610 vout.n609 0.0134551
R1416 vout.n376 vout.n202 0.0134551
R1417 vout.n476 vout.n166 0.0134551
R1418 vout.n514 vout.n483 0.0134551
R1419 vout.n278 vout.n277 0.0132292
R1420 vout.n279 vout.n278 0.0132292
R1421 vout.n279 vout.n265 0.0132292
R1422 vout.n288 vout.n265 0.0132292
R1423 vout.n289 vout.n288 0.0132292
R1424 vout.n290 vout.n289 0.0132292
R1425 vout.n290 vout.n260 0.0132292
R1426 vout.n295 vout.n260 0.0132292
R1427 vout.n296 vout.n295 0.0132292
R1428 vout.n296 vout.n254 0.0132292
R1429 vout.n305 vout.n254 0.0132292
R1430 vout.n306 vout.n305 0.0132292
R1431 vout.n307 vout.n306 0.0132292
R1432 vout.n307 vout.n249 0.0132292
R1433 vout.n312 vout.n249 0.0132292
R1434 vout.n313 vout.n312 0.0132292
R1435 vout.n313 vout.n244 0.0132292
R1436 vout.n321 vout.n244 0.0132292
R1437 vout.n322 vout.n321 0.0132292
R1438 vout.n323 vout.n322 0.0132292
R1439 vout.n323 vout.n239 0.0132292
R1440 vout.n328 vout.n239 0.0132292
R1441 vout.n329 vout.n328 0.0132292
R1442 vout.n329 vout.n231 0.0132292
R1443 vout.n334 vout.n229 0.0132292
R1444 vout.n338 vout.n229 0.0132292
R1445 vout.n339 vout.n338 0.0132292
R1446 vout.n339 vout.n224 0.0132292
R1447 vout.n347 vout.n224 0.0132292
R1448 vout.n348 vout.n347 0.0132292
R1449 vout.n349 vout.n348 0.0132292
R1450 vout.n349 vout.n219 0.0132292
R1451 vout.n354 vout.n219 0.0132292
R1452 vout.n355 vout.n354 0.0132292
R1453 vout.n355 vout.n214 0.0132292
R1454 vout.n359 vout.n214 0.0132292
R1455 vout.n360 vout.n359 0.0132292
R1456 vout.n213 vout.n203 0.0132292
R1457 vout.n377 vout.n203 0.0132292
R1458 vout.n378 vout.n377 0.0132292
R1459 vout.n378 vout.n198 0.0132292
R1460 vout.n386 vout.n198 0.0132292
R1461 vout.n387 vout.n386 0.0132292
R1462 vout.n388 vout.n387 0.0132292
R1463 vout.n388 vout.n193 0.0132292
R1464 vout.n393 vout.n193 0.0132292
R1465 vout.n394 vout.n393 0.0132292
R1466 vout.n394 vout.n185 0.0132292
R1467 vout.n400 vout.n399 0.0132292
R1468 vout.n400 vout.n182 0.0132292
R1469 vout.n408 vout.n182 0.0132292
R1470 vout.n409 vout.n408 0.0132292
R1471 vout.n410 vout.n409 0.0132292
R1472 vout.n410 vout.n177 0.0132292
R1473 vout.n415 vout.n177 0.0132292
R1474 vout.n416 vout.n415 0.0132292
R1475 vout.n416 vout.n172 0.0132292
R1476 vout.n424 vout.n172 0.0132292
R1477 vout.n425 vout.n424 0.0132292
R1478 vout.n426 vout.n425 0.0132292
R1479 vout.n426 vout.n167 0.0132292
R1480 vout.n435 vout.n167 0.0132292
R1481 vout.n436 vout.n435 0.0132292
R1482 vout.n475 vout.n436 0.0132292
R1483 vout.n475 vout.n474 0.0132292
R1484 vout.n474 vout.n437 0.0132292
R1485 vout.n470 vout.n437 0.0132292
R1486 vout.n470 vout.n469 0.0132292
R1487 vout.n469 vout.n442 0.0132292
R1488 vout.n464 vout.n442 0.0132292
R1489 vout.n464 vout.n463 0.0132292
R1490 vout.n463 vout.n462 0.0132292
R1491 vout.n462 vout.n447 0.0132292
R1492 vout.n23 vout.n14 0.0132292
R1493 vout.n24 vout.n23 0.0132292
R1494 vout.n24 vout.n9 0.0132292
R1495 vout.n28 vout.n9 0.0132292
R1496 vout.n29 vout.n28 0.0132292
R1497 vout.n29 vout.n4 0.0132292
R1498 vout.n37 vout.n4 0.0132292
R1499 vout.n38 vout.n37 0.0132292
R1500 vout.n630 vout.n38 0.0132292
R1501 vout.n630 vout.n629 0.0132292
R1502 vout.n629 vout.n628 0.0132292
R1503 vout.n628 vout.n39 0.0132292
R1504 vout.n624 vout.n39 0.0132292
R1505 vout.n624 vout.n623 0.0132292
R1506 vout.n623 vout.n48 0.0132292
R1507 vout.n619 vout.n48 0.0132292
R1508 vout.n619 vout.n618 0.0132292
R1509 vout.n618 vout.n53 0.0132292
R1510 vout.n613 vout.n53 0.0132292
R1511 vout.n613 vout.n612 0.0132292
R1512 vout.n612 vout.n611 0.0132292
R1513 vout.n611 vout.n58 0.0132292
R1514 vout.n606 vout.n58 0.0132292
R1515 vout.n606 vout.n605 0.0132292
R1516 vout.n604 vout.n72 0.0132292
R1517 vout.n599 vout.n72 0.0132292
R1518 vout.n599 vout.n598 0.0132292
R1519 vout.n598 vout.n597 0.0132292
R1520 vout.n597 vout.n86 0.0132292
R1521 vout.n592 vout.n86 0.0132292
R1522 vout.n592 vout.n591 0.0132292
R1523 vout.n591 vout.n590 0.0132292
R1524 vout.n590 vout.n91 0.0132292
R1525 vout.n586 vout.n91 0.0132292
R1526 vout.n586 vout.n585 0.0132292
R1527 vout.n585 vout.n100 0.0132292
R1528 vout.n580 vout.n100 0.0132292
R1529 vout.n580 vout.n579 0.0132292
R1530 vout.n579 vout.n578 0.0132292
R1531 vout.n578 vout.n105 0.0132292
R1532 vout.n573 vout.n105 0.0132292
R1533 vout.n573 vout.n572 0.0132292
R1534 vout.n572 vout.n571 0.0132292
R1535 vout.n571 vout.n111 0.0132292
R1536 vout.n567 vout.n111 0.0132292
R1537 vout.n567 vout.n566 0.0132292
R1538 vout.n566 vout.n120 0.0132292
R1539 vout.n562 vout.n120 0.0132292
R1540 vout.n562 vout.n561 0.0132292
R1541 vout.n561 vout.n125 0.0132292
R1542 vout.n557 vout.n125 0.0132292
R1543 vout.n557 vout.n556 0.0132292
R1544 vout.n556 vout.n546 0.0132292
R1545 vout.n545 vout.n130 0.0132292
R1546 vout.n540 vout.n130 0.0132292
R1547 vout.n540 vout.n539 0.0132292
R1548 vout.n539 vout.n538 0.0132292
R1549 vout.n538 vout.n142 0.0132292
R1550 vout.n533 vout.n142 0.0132292
R1551 vout.n533 vout.n532 0.0132292
R1552 vout.n532 vout.n531 0.0132292
R1553 vout.n531 vout.n147 0.0132292
R1554 vout.n527 vout.n147 0.0132292
R1555 vout.n527 vout.n526 0.0132292
R1556 vout.n526 vout.n156 0.0132292
R1557 vout.n522 vout.n156 0.0132292
R1558 vout.n522 vout.n521 0.0132292
R1559 vout.n521 vout.n161 0.0132292
R1560 vout.n516 vout.n161 0.0132292
R1561 vout.n516 vout.n515 0.0132292
R1562 vout.n515 vout.n484 0.0132292
R1563 vout.n511 vout.n484 0.0132292
R1564 vout.n511 vout.n510 0.0132292
R1565 vout.n510 vout.n489 0.0132292
R1566 vout.n505 vout.n489 0.0132292
R1567 vout.n505 vout.n504 0.0132292
R1568 vout.n504 vout.n503 0.0132292
R1569 vout.n345 vout.n223 0.0128526
R1570 vout.n406 vout.n181 0.0128526
R1571 vout.n537 vout.n536 0.0128526
R1572 vout.n303 vout.n253 0.0125513
R1573 vout.n311 vout.n248 0.0125513
R1574 vout.n560 vout.n124 0.0124006
R1575 vout.n353 vout.n218 0.01225
R1576 vout.n414 vout.n176 0.01225
R1577 vout.n27 vout.n8 0.01225
R1578 vout.n622 vout.n47 0.0116474
R1579 vout.n429 vout.n428 0.0116474
R1580 vout.n502 vout.n501 0.0116474
R1581 vout.n577 vout.n576 0.0114968
R1582 vout.n292 vout.n291 0.0113462
R1583 vout.n326 vout.n325 0.0113462
R1584 vout.n595 vout.n594 0.0111955
R1585 vout.n520 vout.n160 0.0110449
R1586 vout.n391 vout.n390 0.0104423
R1587 vout.n392 vout.n192 0.0104423
R1588 vout.n466 vout.n465 0.0104423
R1589 vout.n451 vout.n446 0.0104423
R1590 vout.n151 vout.n146 0.0104423
R1591 vout.n577 vout.n106 0.010141
R1592 vout.n565 vout.n119 0.00999038
R1593 vout.n36 vout.n35 0.00968342
R1594 vout.n286 vout.n264 0.00953846
R1595 vout.n327 vout.n238 0.00953846
R1596 vout.n434 vout.n433 0.00923718
R1597 vout.n627 vout.n43 0.00912917
R1598 vout.n115 vout.n110 0.00908654
R1599 vout.n601 vout.n600 0.00878526
R1600 vout.n352 vout.n351 0.00863461
R1601 vout.n373 vout.n210 0.00863461
R1602 vout.n413 vout.n412 0.00863461
R1603 vout.n525 vout.n155 0.00863461
R1604 vout.n309 vout.n308 0.00833333
R1605 vout.n310 vout.n309 0.00833333
R1606 vout.n351 vout.n350 0.00803205
R1607 vout.n412 vout.n411 0.00803205
R1608 vout.n528 vout.n155 0.00803205
R1609 vout.n602 vout.n601 0.00788141
R1610 vout.n570 vout.n115 0.00758013
R1611 vout.n375 vout.n374 0.00742949
R1612 vout.n433 vout.n162 0.00742949
R1613 vout.n373 vout.n211 0.00735273
R1614 vout.n372 vout.n371 0.00735273
R1615 vout.n367 vout.n361 0.00735273
R1616 vout.n367 vout.n212 0.00735273
R1617 vout.n369 vout.n213 0.00735273
R1618 vout.n370 vout.n369 0.00735273
R1619 vout.n368 vout.n211 0.00735273
R1620 vout.n373 vout.n372 0.00735273
R1621 vout.n370 vout.n212 0.00735273
R1622 vout.n361 vout.n360 0.00735273
R1623 vout.n43 vout.n3 0.00729874
R1624 vout.n287 vout.n286 0.00712821
R1625 vout.n330 vout.n238 0.00712821
R1626 vout.n71 vout.n70 0.00682692
R1627 vout.n35 vout.n2 0.00670755
R1628 vout.n568 vout.n119 0.00667628
R1629 vout.n106 vout.n104 0.00652564
R1630 vout.n81 vout.n80 0.00622436
R1631 vout.n390 vout.n389 0.00622436
R1632 vout.n395 vout.n192 0.00622436
R1633 vout.n467 vout.n466 0.00622436
R1634 vout.n461 vout.n451 0.00622436
R1635 vout.n530 vout.n151 0.00622436
R1636 vout.n336 vout.n335 0.00562179
R1637 vout.n374 vout.n373 0.00562179
R1638 vout.n523 vout.n160 0.00562179
R1639 vout.n596 vout.n595 0.00547115
R1640 vout.n293 vout.n292 0.00532051
R1641 vout.n325 vout.n324 0.00532051
R1642 vout.n576 vout.n575 0.00516987
R1643 vout.n625 vout.n47 0.00501923
R1644 vout.n428 vout.n427 0.00501923
R1645 vout.n356 vout.n218 0.00441667
R1646 vout.n417 vout.n176 0.00441667
R1647 vout.n30 vout.n8 0.00441667
R1648 vout.n563 vout.n124 0.00426603
R1649 vout.n304 vout.n303 0.00411538
R1650 vout.n314 vout.n248 0.00411538
R1651 vout.n346 vout.n345 0.0038141
R1652 vout.n407 vout.n406 0.0038141
R1653 vout.n536 vout.n535 0.0038141
R1654 vout.n255 vout.n0 0.0037247
R1655 vout.n362 vout.t305 0.00340698
R1656 vout.n363 vout.t302 0.00340698
R1657 vout.n478 vout.t304 0.00340698
R1658 vout.n479 vout.t301 0.00340698
R1659 vout.n633 vout.t303 0.00340698
R1660 vout.n1 vout.t300 0.00340698
R1661 vout.n609 vout.n608 0.00321154
R1662 vout.n379 vout.n202 0.00321154
R1663 vout.n473 vout.n166 0.00321154
R1664 vout.n517 vout.n483 0.00321154
R1665 vout.n255 vout.n1 0.00310198
R1666 vout.n95 vout.n90 0.0030609
R1667 vout.n281 vout.n280 0.00291026
R1668 vout.n582 vout.n581 0.00275962
R1669 vout.n620 vout.n52 0.00260897
R1670 vout.n507 vout.n506 0.00260897
R1671 vout.n276 vout.n275 0.00230769
R1672 vout.n70 vout.n69 0.00200641
R1673 vout.n385 vout.n384 0.00200641
R1674 vout.n471 vout.n441 0.00200641
R1675 vout.n25 vout.n13 0.00200641
R1676 vout.n304 vout.n299 0.00185577
R1677 vout.n558 vout.n129 0.00185577
R1678 vout.n634 vout.n633 0.00184207
R1679 vout.n632 vout.n631 0.00183019
R1680 vout.n477 vout.n162 0.00155449
R1681 vout.n519 vout.n518 0.00155449
R1682 vout.n340 vout.n228 0.00140385
R1683 vout.n401 vout.n184 0.00140385
R1684 vout.n542 vout.n541 0.00140385
R1685 vout.n297 vout.n259 0.00110256
R1686 vout.n320 vout.n319 0.00110256
R1687 vout.n615 vout.n614 0.000801282
R1688 vout.n358 vout.n210 0.000801282
R1689 vout.n423 vout.n422 0.000801282
R1690 vout.n512 vout.n488 0.000801282
R1691 vout.n587 vout.n99 0.000650641
R1692 vss.n3029 vss.n3028 8.28156e+06
R1693 vss.n3028 vss.n3025 95564.8
R1694 vss.n2275 vss.n2250 39475.3
R1695 vss.n2279 vss.n2250 39475.3
R1696 vss.n2275 vss.n2261 39475.3
R1697 vss.n2279 vss.n2261 39475.3
R1698 vss.n3028 vss.n3027 17199.2
R1699 vss.n5913 vss.n221 10707.5
R1700 vss.n5914 vss.n221 10707.5
R1701 vss.n5919 vss.n216 10707.5
R1702 vss.n5919 vss.n217 10707.5
R1703 vss.n5913 vss.n225 5788.32
R1704 vss.n225 vss.n216 5788.32
R1705 vss.n5914 vss.n222 5788.32
R1706 vss.n222 vss.n217 5788.32
R1707 vss.n2640 vss.n225 4919.21
R1708 vss.n2640 vss.n222 4919.21
R1709 vss.n2276 vss.n2262 2564.89
R1710 vss.n2278 vss.n2262 2564.89
R1711 vss.n2277 vss.n2276 2564.89
R1712 vss.n2278 vss.n2277 2564.89
R1713 vss.n2300 vss.n2232 2161.21
R1714 vss.n2301 vss.n2232 2161.21
R1715 vss.n5529 vss.n304 2161.21
R1716 vss.n5529 vss.n305 2161.21
R1717 vss.n2436 vss.n2383 1245.74
R1718 vss.n2436 vss.n2384 1245.74
R1719 vss.n2402 vss.n2328 1245.74
R1720 vss.n2402 vss.n2332 1245.74
R1721 vss.n2970 vss.n2202 1245.74
R1722 vss.n2970 vss.n2331 1245.74
R1723 vss.n4224 vss.n1306 1245.74
R1724 vss.n4224 vss.n1307 1245.74
R1725 vss.n2224 vss.n2204 1245.74
R1726 vss.n2224 vss.n2206 1245.74
R1727 vss.n2300 vss.n2204 915.471
R1728 vss.n2323 vss.n2204 915.471
R1729 vss.n2323 vss.n1306 915.471
R1730 vss.n3019 vss.n1306 915.471
R1731 vss.n3019 vss.n2202 915.471
R1732 vss.n3015 vss.n2202 915.471
R1733 vss.n3015 vss.n2328 915.471
R1734 vss.n2416 vss.n2328 915.471
R1735 vss.n2416 vss.n2383 915.471
R1736 vss.n2383 vss.n304 915.471
R1737 vss.n2301 vss.n2206 915.471
R1738 vss.n2322 vss.n2206 915.471
R1739 vss.n2322 vss.n1307 915.471
R1740 vss.n2201 vss.n1307 915.471
R1741 vss.n2331 vss.n2201 915.471
R1742 vss.n3014 vss.n2331 915.471
R1743 vss.n3014 vss.n2332 915.471
R1744 vss.n2413 vss.n2332 915.471
R1745 vss.n2413 vss.n2384 915.471
R1746 vss.n2384 vss.n305 915.471
R1747 vss.n4587 vss.n4586 696.351
R1748 vss.n5918 vss.n5917 695.718
R1749 vss.n5915 vss.n220 695.718
R1750 vss.n3027 vss.n3026 686.067
R1751 vss.n5148 vss.n1115 590.609
R1752 vss.n939 vss.n880 590.609
R1753 vss.n1116 vss.n1115 590.609
R1754 vss.n907 vss.n880 590.609
R1755 vss.n5144 vss.n1115 590.609
R1756 vss.n965 vss.n880 590.609
R1757 vss.n1261 vss.n1115 590.609
R1758 vss.n5330 vss.n880 590.609
R1759 vss.n5022 vss.n1115 590.609
R1760 vss.n995 vss.n880 590.609
R1761 vss.n4743 vss.n1115 590.609
R1762 vss.n4865 vss.n880 590.609
R1763 vss.n4235 vss.n1115 590.609
R1764 vss.n4237 vss.n880 590.609
R1765 vss.n4589 vss.n1115 590.609
R1766 vss.n4711 vss.n880 590.609
R1767 vss.n4329 vss.n1115 590.609
R1768 vss.n4348 vss.n1033 585
R1769 vss.n5182 vss.n1050 585
R1770 vss.n4345 vss.n1045 585
R1771 vss.n5176 vss.n1062 585
R1772 vss.n4342 vss.n1057 585
R1773 vss.n5170 vss.n1074 585
R1774 vss.n4339 vss.n1069 585
R1775 vss.n5164 vss.n1086 585
R1776 vss.n4336 vss.n1081 585
R1777 vss.n5158 vss.n1098 585
R1778 vss.n4333 vss.n1093 585
R1779 vss.n5152 vss.n1110 585
R1780 vss.n4330 vss.n1105 585
R1781 vss.n5146 vss.n1290 585
R1782 vss.n4608 vss.n1033 585
R1783 vss.n5182 vss.n1049 585
R1784 vss.n4605 vss.n1045 585
R1785 vss.n5176 vss.n1061 585
R1786 vss.n4602 vss.n1057 585
R1787 vss.n5170 vss.n1073 585
R1788 vss.n4599 vss.n1069 585
R1789 vss.n5164 vss.n1085 585
R1790 vss.n4596 vss.n1081 585
R1791 vss.n5158 vss.n1097 585
R1792 vss.n4593 vss.n1093 585
R1793 vss.n5152 vss.n1109 585
R1794 vss.n4590 vss.n1105 585
R1795 vss.n5146 vss.n1289 585
R1796 vss.n5001 vss.n1033 585
R1797 vss.n5182 vss.n1052 585
R1798 vss.n5004 vss.n1045 585
R1799 vss.n5176 vss.n1064 585
R1800 vss.n5007 vss.n1057 585
R1801 vss.n5170 vss.n1076 585
R1802 vss.n5010 vss.n1069 585
R1803 vss.n5164 vss.n1088 585
R1804 vss.n5013 vss.n1081 585
R1805 vss.n5158 vss.n1100 585
R1806 vss.n5016 vss.n1093 585
R1807 vss.n5152 vss.n1112 585
R1808 vss.n5020 vss.n1105 585
R1809 vss.n5146 vss.n5021 585
R1810 vss.n4762 vss.n1033 585
R1811 vss.n5182 vss.n1048 585
R1812 vss.n4759 vss.n1045 585
R1813 vss.n5176 vss.n1060 585
R1814 vss.n4756 vss.n1057 585
R1815 vss.n5170 vss.n1072 585
R1816 vss.n4753 vss.n1069 585
R1817 vss.n5164 vss.n1084 585
R1818 vss.n4750 vss.n1081 585
R1819 vss.n5158 vss.n1096 585
R1820 vss.n4747 vss.n1093 585
R1821 vss.n5152 vss.n1108 585
R1822 vss.n4744 vss.n1105 585
R1823 vss.n5146 vss.n1288 585
R1824 vss.n5123 vss.n1033 585
R1825 vss.n5182 vss.n1053 585
R1826 vss.n5126 vss.n1045 585
R1827 vss.n5176 vss.n1065 585
R1828 vss.n5129 vss.n1057 585
R1829 vss.n5170 vss.n1077 585
R1830 vss.n5132 vss.n1069 585
R1831 vss.n5164 vss.n1089 585
R1832 vss.n5135 vss.n1081 585
R1833 vss.n5158 vss.n1101 585
R1834 vss.n5138 vss.n1093 585
R1835 vss.n5152 vss.n1113 585
R1836 vss.n5142 vss.n1105 585
R1837 vss.n5146 vss.n5143 585
R1838 vss.n1267 vss.n1033 585
R1839 vss.n5182 vss.n1047 585
R1840 vss.n1270 vss.n1045 585
R1841 vss.n5176 vss.n1059 585
R1842 vss.n1273 vss.n1057 585
R1843 vss.n5170 vss.n1071 585
R1844 vss.n1276 vss.n1069 585
R1845 vss.n5164 vss.n1083 585
R1846 vss.n1279 vss.n1081 585
R1847 vss.n5158 vss.n1095 585
R1848 vss.n1282 vss.n1093 585
R1849 vss.n5152 vss.n1107 585
R1850 vss.n1286 vss.n1105 585
R1851 vss.n5146 vss.n1287 585
R1852 vss.n1033 vss.n1032 585
R1853 vss.n5182 vss.n5181 585
R1854 vss.n1054 vss.n1045 585
R1855 vss.n5177 vss.n5176 585
R1856 vss.n1057 vss.n1056 585
R1857 vss.n5170 vss.n5169 585
R1858 vss.n1078 vss.n1069 585
R1859 vss.n5165 vss.n5164 585
R1860 vss.n1081 vss.n1080 585
R1861 vss.n5158 vss.n5157 585
R1862 vss.n1102 vss.n1093 585
R1863 vss.n5153 vss.n5152 585
R1864 vss.n1105 vss.n1104 585
R1865 vss.n5146 vss.n5145 585
R1866 vss.n1240 vss.n1033 585
R1867 vss.n5182 vss.n1046 585
R1868 vss.n1243 vss.n1045 585
R1869 vss.n5176 vss.n1058 585
R1870 vss.n1246 vss.n1057 585
R1871 vss.n5170 vss.n1070 585
R1872 vss.n1249 vss.n1069 585
R1873 vss.n5164 vss.n1082 585
R1874 vss.n1252 vss.n1081 585
R1875 vss.n5158 vss.n1094 585
R1876 vss.n1255 vss.n1093 585
R1877 vss.n5152 vss.n1106 585
R1878 vss.n1259 vss.n1105 585
R1879 vss.n5146 vss.n1260 585
R1880 vss.n1042 vss.n1033 585
R1881 vss.n5183 vss.n5182 585
R1882 vss.n1045 vss.n1044 585
R1883 vss.n5176 vss.n5175 585
R1884 vss.n1066 vss.n1057 585
R1885 vss.n5171 vss.n5170 585
R1886 vss.n1069 vss.n1068 585
R1887 vss.n5164 vss.n5163 585
R1888 vss.n1090 vss.n1081 585
R1889 vss.n5159 vss.n5158 585
R1890 vss.n1093 vss.n1092 585
R1891 vss.n5152 vss.n5151 585
R1892 vss.n1114 vss.n1105 585
R1893 vss.n5147 vss.n5146 585
R1894 vss.n2284 vss.n2248 585
R1895 vss.n2284 vss.n2283 585
R1896 vss.n2285 vss.n2241 585
R1897 vss.n2286 vss.n2285 585
R1898 vss.n2242 vss.n2215 585
R1899 vss.n2234 vss.n2215 585
R1900 vss.n2310 vss.n2209 585
R1901 vss.n2310 vss.n2309 585
R1902 vss.n2312 vss.n2311 585
R1903 vss.n2311 vss.n1291 585
R1904 vss.n2214 vss.n1292 585
R1905 vss.n4233 vss.n1292 585
R1906 vss.n2213 vss.n2212 585
R1907 vss.n2212 vss.n2211 585
R1908 vss.n2210 vss.n1304 585
R1909 vss.n4227 vss.n1304 585
R1910 vss.n2195 vss.n1311 585
R1911 vss.n2195 vss.n2194 585
R1912 vss.n2197 vss.n2196 585
R1913 vss.n3024 vss.n2196 585
R1914 vss.n2199 vss.n2198 585
R1915 vss.n2200 vss.n2199 585
R1916 vss.n1324 vss.n1317 585
R1917 vss.n4206 vss.n1324 585
R1918 vss.n2981 vss.n2980 585
R1919 vss.n2980 vss.n2979 585
R1920 vss.n2984 vss.n2967 585
R1921 vss.n2989 vss.n2967 585
R1922 vss.n2983 vss.n2982 585
R1923 vss.n2982 vss.n2330 585
R1924 vss.n2342 vss.n2336 585
R1925 vss.n3007 vss.n2342 585
R1926 vss.n2394 vss.n2392 585
R1927 vss.n2400 vss.n2394 585
R1928 vss.n2423 vss.n2422 585
R1929 vss.n2422 vss.n2421 585
R1930 vss.n2424 vss.n2386 585
R1931 vss.n2417 vss.n2386 585
R1932 vss.n2246 vss.n2245 585
R1933 vss.n2283 vss.n2246 585
R1934 vss.n2288 vss.n2287 585
R1935 vss.n2287 vss.n2286 585
R1936 vss.n2229 vss.n2228 585
R1937 vss.n2234 vss.n2228 585
R1938 vss.n2308 vss.n2307 585
R1939 vss.n2309 vss.n2308 585
R1940 vss.n1297 vss.n1295 585
R1941 vss.n1295 vss.n1291 585
R1942 vss.n4232 vss.n4231 585
R1943 vss.n4233 vss.n4232 585
R1944 vss.n4230 vss.n1296 585
R1945 vss.n2211 vss.n1296 585
R1946 vss.n4229 vss.n4228 585
R1947 vss.n4228 vss.n4227 585
R1948 vss.n1302 vss.n1301 585
R1949 vss.n2194 vss.n1302 585
R1950 vss.n3023 vss.n3022 585
R1951 vss.n3024 vss.n3023 585
R1952 vss.n1321 vss.n1319 585
R1953 vss.n2200 vss.n1321 585
R1954 vss.n4208 vss.n4207 585
R1955 vss.n4207 vss.n4206 585
R1956 vss.n1322 vss.n1320 585
R1957 vss.n2979 vss.n1322 585
R1958 vss.n2988 vss.n2987 585
R1959 vss.n2989 vss.n2988 585
R1960 vss.n2340 vss.n2338 585
R1961 vss.n2340 vss.n2330 585
R1962 vss.n3009 vss.n3008 585
R1963 vss.n3008 vss.n3007 585
R1964 vss.n2341 vss.n2339 585
R1965 vss.n2400 vss.n2341 585
R1966 vss.n2420 vss.n2390 585
R1967 vss.n2421 vss.n2420 585
R1968 vss.n2427 vss.n2389 585
R1969 vss.n2417 vss.n2389 585
R1970 vss.n5364 vss.n848 585
R1971 vss.n853 vss.n834 585
R1972 vss.n5370 vss.n836 585
R1973 vss.n835 vss.n815 585
R1974 vss.n5374 vss.n816 585
R1975 vss.n821 vss.n799 585
R1976 vss.n5380 vss.n801 585
R1977 vss.n800 vss.n782 585
R1978 vss.n5384 vss.n783 585
R1979 vss.n4577 vss.n766 585
R1980 vss.n5390 vss.n767 585
R1981 vss.n4581 vss.n754 585
R1982 vss.n5394 vss.n753 585
R1983 vss.n5364 vss.n846 585
R1984 vss.n854 vss.n834 585
R1985 vss.n5370 vss.n833 585
R1986 vss.n832 vss.n815 585
R1987 vss.n5374 vss.n813 585
R1988 vss.n822 vss.n799 585
R1989 vss.n5380 vss.n798 585
R1990 vss.n797 vss.n782 585
R1991 vss.n5384 vss.n781 585
R1992 vss.n4578 vss.n766 585
R1993 vss.n5390 vss.n765 585
R1994 vss.n4582 vss.n754 585
R1995 vss.n5394 vss.n755 585
R1996 vss.n4588 vss.n4266 585
R1997 vss.n5406 vss.n734 585
R1998 vss.n4571 vss.n719 585
R1999 vss.n5410 vss.n720 585
R2000 vss.n4269 vss.n705 585
R2001 vss.n5414 vss.n706 585
R2002 vss.n4563 vss.n691 585
R2003 vss.n5418 vss.n692 585
R2004 vss.n4555 vss.n677 585
R2005 vss.n5422 vss.n678 585
R2006 vss.n4274 vss.n663 585
R2007 vss.n5426 vss.n664 585
R2008 vss.n4543 vss.n649 585
R2009 vss.n5430 vss.n650 585
R2010 vss.n4535 vss.n635 585
R2011 vss.n5434 vss.n636 585
R2012 vss.n4279 vss.n621 585
R2013 vss.n5438 vss.n622 585
R2014 vss.n4523 vss.n607 585
R2015 vss.n5442 vss.n608 585
R2016 vss.n4515 vss.n593 585
R2017 vss.n5446 vss.n594 585
R2018 vss.n4284 vss.n579 585
R2019 vss.n5450 vss.n580 585
R2020 vss.n4503 vss.n565 585
R2021 vss.n5454 vss.n566 585
R2022 vss.n4497 vss.n551 585
R2023 vss.n5458 vss.n552 585
R2024 vss.n4493 vss.n537 585
R2025 vss.n5462 vss.n538 585
R2026 vss.n4486 vss.n523 585
R2027 vss.n5466 vss.n524 585
R2028 vss.n4481 vss.n509 585
R2029 vss.n5470 vss.n510 585
R2030 vss.n4473 vss.n495 585
R2031 vss.n5474 vss.n496 585
R2032 vss.n4294 vss.n481 585
R2033 vss.n5478 vss.n482 585
R2034 vss.n4461 vss.n467 585
R2035 vss.n5482 vss.n468 585
R2036 vss.n4453 vss.n453 585
R2037 vss.n5486 vss.n454 585
R2038 vss.n4299 vss.n439 585
R2039 vss.n5490 vss.n440 585
R2040 vss.n4441 vss.n425 585
R2041 vss.n5494 vss.n426 585
R2042 vss.n4433 vss.n411 585
R2043 vss.n5498 vss.n412 585
R2044 vss.n4304 vss.n397 585
R2045 vss.n5502 vss.n398 585
R2046 vss.n4308 vss.n383 585
R2047 vss.n5506 vss.n384 585
R2048 vss.n4416 vss.n369 585
R2049 vss.n5510 vss.n370 585
R2050 vss.n4410 vss.n355 585
R2051 vss.n5514 vss.n356 585
R2052 vss.n4403 vss.n341 585
R2053 vss.n5518 vss.n342 585
R2054 vss.n4316 vss.n327 585
R2055 vss.n5522 vss.n328 585
R2056 vss.n4319 vss.n313 585
R2057 vss.n5526 vss.n314 585
R2058 vss.n4387 vss.n308 585
R2059 vss.n5208 vss.n1013 585
R2060 vss.n4356 vss.n1009 585
R2061 vss.n5201 vss.n1026 585
R2062 vss.n4327 vss.n1021 585
R2063 vss.n5188 vss.n1038 585
R2064 vss.n5364 vss.n849 585
R2065 vss.n4722 vss.n834 585
R2066 vss.n5370 vss.n837 585
R2067 vss.n4725 vss.n815 585
R2068 vss.n5374 vss.n817 585
R2069 vss.n4728 vss.n799 585
R2070 vss.n5380 vss.n802 585
R2071 vss.n4731 vss.n782 585
R2072 vss.n5384 vss.n784 585
R2073 vss.n4734 vss.n766 585
R2074 vss.n5390 vss.n768 585
R2075 vss.n4737 vss.n754 585
R2076 vss.n5394 vss.n750 585
R2077 vss.n4742 vss.n4741 585
R2078 vss.n4742 vss.n215 585
R2079 vss.n5406 vss.n732 585
R2080 vss.n4707 vss.n719 585
R2081 vss.n5410 vss.n718 585
R2082 vss.n4704 vss.n705 585
R2083 vss.n5414 vss.n704 585
R2084 vss.n4701 vss.n691 585
R2085 vss.n5418 vss.n690 585
R2086 vss.n4698 vss.n677 585
R2087 vss.n5422 vss.n676 585
R2088 vss.n4695 vss.n663 585
R2089 vss.n5426 vss.n662 585
R2090 vss.n4692 vss.n649 585
R2091 vss.n5430 vss.n648 585
R2092 vss.n4689 vss.n635 585
R2093 vss.n5434 vss.n634 585
R2094 vss.n4686 vss.n621 585
R2095 vss.n5438 vss.n620 585
R2096 vss.n4683 vss.n607 585
R2097 vss.n5442 vss.n606 585
R2098 vss.n4680 vss.n593 585
R2099 vss.n5446 vss.n592 585
R2100 vss.n4677 vss.n579 585
R2101 vss.n5450 vss.n578 585
R2102 vss.n4674 vss.n565 585
R2103 vss.n5454 vss.n564 585
R2104 vss.n4671 vss.n551 585
R2105 vss.n5458 vss.n550 585
R2106 vss.n4668 vss.n537 585
R2107 vss.n5462 vss.n536 585
R2108 vss.n4665 vss.n523 585
R2109 vss.n5466 vss.n522 585
R2110 vss.n4662 vss.n509 585
R2111 vss.n5470 vss.n508 585
R2112 vss.n4659 vss.n495 585
R2113 vss.n5474 vss.n494 585
R2114 vss.n4656 vss.n481 585
R2115 vss.n5478 vss.n480 585
R2116 vss.n4653 vss.n467 585
R2117 vss.n5482 vss.n466 585
R2118 vss.n4650 vss.n453 585
R2119 vss.n5486 vss.n452 585
R2120 vss.n4647 vss.n439 585
R2121 vss.n5490 vss.n438 585
R2122 vss.n4644 vss.n425 585
R2123 vss.n5494 vss.n424 585
R2124 vss.n4641 vss.n411 585
R2125 vss.n5498 vss.n410 585
R2126 vss.n4638 vss.n397 585
R2127 vss.n5502 vss.n396 585
R2128 vss.n4635 vss.n383 585
R2129 vss.n5506 vss.n382 585
R2130 vss.n4632 vss.n369 585
R2131 vss.n5510 vss.n368 585
R2132 vss.n4629 vss.n355 585
R2133 vss.n5514 vss.n354 585
R2134 vss.n4626 vss.n341 585
R2135 vss.n5518 vss.n340 585
R2136 vss.n4623 vss.n327 585
R2137 vss.n5522 vss.n326 585
R2138 vss.n4620 vss.n313 585
R2139 vss.n5526 vss.n312 585
R2140 vss.n4617 vss.n308 585
R2141 vss.n5208 vss.n1012 585
R2142 vss.n4614 vss.n1009 585
R2143 vss.n5201 vss.n1025 585
R2144 vss.n4611 vss.n1021 585
R2145 vss.n5188 vss.n1037 585
R2146 vss.n5364 vss.n845 585
R2147 vss.n4248 vss.n834 585
R2148 vss.n5370 vss.n831 585
R2149 vss.n4251 vss.n815 585
R2150 vss.n5374 vss.n812 585
R2151 vss.n4254 vss.n799 585
R2152 vss.n5380 vss.n796 585
R2153 vss.n4257 vss.n782 585
R2154 vss.n5384 vss.n780 585
R2155 vss.n4260 vss.n766 585
R2156 vss.n5390 vss.n764 585
R2157 vss.n4263 vss.n754 585
R2158 vss.n5394 vss.n756 585
R2159 vss.n4899 vss.n4898 585
R2160 vss.n5406 vss.n735 585
R2161 vss.n4902 vss.n719 585
R2162 vss.n5410 vss.n722 585
R2163 vss.n4905 vss.n705 585
R2164 vss.n5414 vss.n708 585
R2165 vss.n4908 vss.n691 585
R2166 vss.n5418 vss.n694 585
R2167 vss.n4911 vss.n677 585
R2168 vss.n5422 vss.n680 585
R2169 vss.n4914 vss.n663 585
R2170 vss.n5426 vss.n666 585
R2171 vss.n4917 vss.n649 585
R2172 vss.n5430 vss.n652 585
R2173 vss.n4920 vss.n635 585
R2174 vss.n5434 vss.n638 585
R2175 vss.n4923 vss.n621 585
R2176 vss.n5438 vss.n624 585
R2177 vss.n4926 vss.n607 585
R2178 vss.n5442 vss.n610 585
R2179 vss.n4929 vss.n593 585
R2180 vss.n5446 vss.n596 585
R2181 vss.n4932 vss.n579 585
R2182 vss.n5450 vss.n582 585
R2183 vss.n4935 vss.n565 585
R2184 vss.n5454 vss.n568 585
R2185 vss.n4938 vss.n551 585
R2186 vss.n5458 vss.n554 585
R2187 vss.n4941 vss.n537 585
R2188 vss.n5462 vss.n540 585
R2189 vss.n4944 vss.n523 585
R2190 vss.n5466 vss.n526 585
R2191 vss.n4947 vss.n509 585
R2192 vss.n5470 vss.n512 585
R2193 vss.n4950 vss.n495 585
R2194 vss.n5474 vss.n498 585
R2195 vss.n4953 vss.n481 585
R2196 vss.n5478 vss.n484 585
R2197 vss.n4956 vss.n467 585
R2198 vss.n5482 vss.n470 585
R2199 vss.n4959 vss.n453 585
R2200 vss.n5486 vss.n456 585
R2201 vss.n4962 vss.n439 585
R2202 vss.n5490 vss.n442 585
R2203 vss.n4965 vss.n425 585
R2204 vss.n5494 vss.n428 585
R2205 vss.n4968 vss.n411 585
R2206 vss.n5498 vss.n414 585
R2207 vss.n4971 vss.n397 585
R2208 vss.n5502 vss.n400 585
R2209 vss.n4974 vss.n383 585
R2210 vss.n5506 vss.n386 585
R2211 vss.n4977 vss.n369 585
R2212 vss.n5510 vss.n372 585
R2213 vss.n4980 vss.n355 585
R2214 vss.n5514 vss.n358 585
R2215 vss.n4983 vss.n341 585
R2216 vss.n5518 vss.n344 585
R2217 vss.n4986 vss.n327 585
R2218 vss.n5522 vss.n330 585
R2219 vss.n4989 vss.n313 585
R2220 vss.n5526 vss.n315 585
R2221 vss.n4992 vss.n308 585
R2222 vss.n5208 vss.n1015 585
R2223 vss.n4995 vss.n1009 585
R2224 vss.n5201 vss.n1028 585
R2225 vss.n4998 vss.n1021 585
R2226 vss.n5188 vss.n1040 585
R2227 vss.n5364 vss.n850 585
R2228 vss.n4876 vss.n834 585
R2229 vss.n5370 vss.n838 585
R2230 vss.n4879 vss.n815 585
R2231 vss.n5374 vss.n818 585
R2232 vss.n4882 vss.n799 585
R2233 vss.n5380 vss.n803 585
R2234 vss.n4885 vss.n782 585
R2235 vss.n5384 vss.n785 585
R2236 vss.n4888 vss.n766 585
R2237 vss.n5390 vss.n769 585
R2238 vss.n4891 vss.n754 585
R2239 vss.n5394 vss.n749 585
R2240 vss.n4896 vss.n4895 585
R2241 vss.n5406 vss.n731 585
R2242 vss.n4861 vss.n719 585
R2243 vss.n5410 vss.n717 585
R2244 vss.n4858 vss.n705 585
R2245 vss.n5414 vss.n703 585
R2246 vss.n4855 vss.n691 585
R2247 vss.n5418 vss.n689 585
R2248 vss.n4852 vss.n677 585
R2249 vss.n5422 vss.n675 585
R2250 vss.n4849 vss.n663 585
R2251 vss.n5426 vss.n661 585
R2252 vss.n4846 vss.n649 585
R2253 vss.n5430 vss.n647 585
R2254 vss.n4843 vss.n635 585
R2255 vss.n5434 vss.n633 585
R2256 vss.n4840 vss.n621 585
R2257 vss.n5438 vss.n619 585
R2258 vss.n4837 vss.n607 585
R2259 vss.n5442 vss.n605 585
R2260 vss.n4834 vss.n593 585
R2261 vss.n5446 vss.n591 585
R2262 vss.n4831 vss.n579 585
R2263 vss.n5450 vss.n577 585
R2264 vss.n4828 vss.n565 585
R2265 vss.n5454 vss.n563 585
R2266 vss.n4825 vss.n551 585
R2267 vss.n5458 vss.n549 585
R2268 vss.n4822 vss.n537 585
R2269 vss.n5462 vss.n535 585
R2270 vss.n4819 vss.n523 585
R2271 vss.n5466 vss.n521 585
R2272 vss.n4816 vss.n509 585
R2273 vss.n5470 vss.n507 585
R2274 vss.n4813 vss.n495 585
R2275 vss.n5474 vss.n493 585
R2276 vss.n4810 vss.n481 585
R2277 vss.n5478 vss.n479 585
R2278 vss.n4807 vss.n467 585
R2279 vss.n5482 vss.n465 585
R2280 vss.n4804 vss.n453 585
R2281 vss.n5486 vss.n451 585
R2282 vss.n4801 vss.n439 585
R2283 vss.n5490 vss.n437 585
R2284 vss.n4798 vss.n425 585
R2285 vss.n5494 vss.n423 585
R2286 vss.n4795 vss.n411 585
R2287 vss.n5498 vss.n409 585
R2288 vss.n4792 vss.n397 585
R2289 vss.n5502 vss.n395 585
R2290 vss.n4789 vss.n383 585
R2291 vss.n5506 vss.n381 585
R2292 vss.n4786 vss.n369 585
R2293 vss.n5510 vss.n367 585
R2294 vss.n4783 vss.n355 585
R2295 vss.n5514 vss.n353 585
R2296 vss.n4780 vss.n341 585
R2297 vss.n5518 vss.n339 585
R2298 vss.n4777 vss.n327 585
R2299 vss.n5522 vss.n325 585
R2300 vss.n4774 vss.n313 585
R2301 vss.n5526 vss.n311 585
R2302 vss.n4771 vss.n308 585
R2303 vss.n5208 vss.n1011 585
R2304 vss.n4768 vss.n1009 585
R2305 vss.n5201 vss.n1024 585
R2306 vss.n4765 vss.n1021 585
R2307 vss.n5188 vss.n1036 585
R2308 vss.n5364 vss.n844 585
R2309 vss.n985 vss.n834 585
R2310 vss.n5370 vss.n830 585
R2311 vss.n982 vss.n815 585
R2312 vss.n5374 vss.n811 585
R2313 vss.n979 vss.n799 585
R2314 vss.n5380 vss.n795 585
R2315 vss.n976 vss.n782 585
R2316 vss.n5384 vss.n779 585
R2317 vss.n973 vss.n766 585
R2318 vss.n5390 vss.n763 585
R2319 vss.n754 vss.n745 585
R2320 vss.n5395 vss.n5394 585
R2321 vss.n5397 vss.n5396 585
R2322 vss.n5406 vss.n736 585
R2323 vss.n5024 vss.n719 585
R2324 vss.n5410 vss.n723 585
R2325 vss.n5027 vss.n705 585
R2326 vss.n5414 vss.n709 585
R2327 vss.n5030 vss.n691 585
R2328 vss.n5418 vss.n695 585
R2329 vss.n5033 vss.n677 585
R2330 vss.n5422 vss.n681 585
R2331 vss.n5036 vss.n663 585
R2332 vss.n5426 vss.n667 585
R2333 vss.n5039 vss.n649 585
R2334 vss.n5430 vss.n653 585
R2335 vss.n5042 vss.n635 585
R2336 vss.n5434 vss.n639 585
R2337 vss.n5045 vss.n621 585
R2338 vss.n5438 vss.n625 585
R2339 vss.n5048 vss.n607 585
R2340 vss.n5442 vss.n611 585
R2341 vss.n5051 vss.n593 585
R2342 vss.n5446 vss.n597 585
R2343 vss.n5054 vss.n579 585
R2344 vss.n5450 vss.n583 585
R2345 vss.n5057 vss.n565 585
R2346 vss.n5454 vss.n569 585
R2347 vss.n5060 vss.n551 585
R2348 vss.n5458 vss.n555 585
R2349 vss.n5063 vss.n537 585
R2350 vss.n5462 vss.n541 585
R2351 vss.n5066 vss.n523 585
R2352 vss.n5466 vss.n527 585
R2353 vss.n5069 vss.n509 585
R2354 vss.n5470 vss.n513 585
R2355 vss.n5072 vss.n495 585
R2356 vss.n5474 vss.n499 585
R2357 vss.n5075 vss.n481 585
R2358 vss.n5478 vss.n485 585
R2359 vss.n5078 vss.n467 585
R2360 vss.n5482 vss.n471 585
R2361 vss.n5081 vss.n453 585
R2362 vss.n5486 vss.n457 585
R2363 vss.n5084 vss.n439 585
R2364 vss.n5490 vss.n443 585
R2365 vss.n5087 vss.n425 585
R2366 vss.n5494 vss.n429 585
R2367 vss.n5090 vss.n411 585
R2368 vss.n5498 vss.n415 585
R2369 vss.n5093 vss.n397 585
R2370 vss.n5502 vss.n401 585
R2371 vss.n5096 vss.n383 585
R2372 vss.n5506 vss.n387 585
R2373 vss.n5099 vss.n369 585
R2374 vss.n5510 vss.n373 585
R2375 vss.n5102 vss.n355 585
R2376 vss.n5514 vss.n359 585
R2377 vss.n5105 vss.n341 585
R2378 vss.n5518 vss.n345 585
R2379 vss.n5108 vss.n327 585
R2380 vss.n5522 vss.n331 585
R2381 vss.n5111 vss.n313 585
R2382 vss.n5526 vss.n316 585
R2383 vss.n5114 vss.n308 585
R2384 vss.n5208 vss.n1016 585
R2385 vss.n5117 vss.n1009 585
R2386 vss.n5201 vss.n1029 585
R2387 vss.n5120 vss.n1021 585
R2388 vss.n5188 vss.n1041 585
R2389 vss.n5364 vss.n851 585
R2390 vss.n5320 vss.n834 585
R2391 vss.n5370 vss.n839 585
R2392 vss.n5317 vss.n815 585
R2393 vss.n5374 vss.n819 585
R2394 vss.n5314 vss.n799 585
R2395 vss.n5380 vss.n804 585
R2396 vss.n5311 vss.n782 585
R2397 vss.n5384 vss.n786 585
R2398 vss.n5308 vss.n766 585
R2399 vss.n5390 vss.n770 585
R2400 vss.n5305 vss.n754 585
R2401 vss.n5394 vss.n748 585
R2402 vss.n5399 vss.n742 585
R2403 vss.n5406 vss.n730 585
R2404 vss.n5300 vss.n719 585
R2405 vss.n5410 vss.n716 585
R2406 vss.n5297 vss.n705 585
R2407 vss.n5414 vss.n702 585
R2408 vss.n5294 vss.n691 585
R2409 vss.n5418 vss.n688 585
R2410 vss.n5291 vss.n677 585
R2411 vss.n5422 vss.n674 585
R2412 vss.n5288 vss.n663 585
R2413 vss.n5426 vss.n660 585
R2414 vss.n5285 vss.n649 585
R2415 vss.n5430 vss.n646 585
R2416 vss.n5282 vss.n635 585
R2417 vss.n5434 vss.n632 585
R2418 vss.n5279 vss.n621 585
R2419 vss.n5438 vss.n618 585
R2420 vss.n5276 vss.n607 585
R2421 vss.n5442 vss.n604 585
R2422 vss.n5273 vss.n593 585
R2423 vss.n5446 vss.n590 585
R2424 vss.n5270 vss.n579 585
R2425 vss.n5450 vss.n576 585
R2426 vss.n5267 vss.n565 585
R2427 vss.n5454 vss.n562 585
R2428 vss.n5264 vss.n551 585
R2429 vss.n5458 vss.n548 585
R2430 vss.n5261 vss.n537 585
R2431 vss.n5462 vss.n534 585
R2432 vss.n5258 vss.n523 585
R2433 vss.n5466 vss.n520 585
R2434 vss.n5255 vss.n509 585
R2435 vss.n5470 vss.n506 585
R2436 vss.n5252 vss.n495 585
R2437 vss.n5474 vss.n492 585
R2438 vss.n5249 vss.n481 585
R2439 vss.n5478 vss.n478 585
R2440 vss.n5246 vss.n467 585
R2441 vss.n5482 vss.n464 585
R2442 vss.n5243 vss.n453 585
R2443 vss.n5486 vss.n450 585
R2444 vss.n5240 vss.n439 585
R2445 vss.n5490 vss.n436 585
R2446 vss.n5237 vss.n425 585
R2447 vss.n5494 vss.n422 585
R2448 vss.n5234 vss.n411 585
R2449 vss.n5498 vss.n408 585
R2450 vss.n5231 vss.n397 585
R2451 vss.n5502 vss.n394 585
R2452 vss.n5228 vss.n383 585
R2453 vss.n5506 vss.n380 585
R2454 vss.n5225 vss.n369 585
R2455 vss.n5510 vss.n366 585
R2456 vss.n5222 vss.n355 585
R2457 vss.n5514 vss.n352 585
R2458 vss.n5219 vss.n341 585
R2459 vss.n5518 vss.n338 585
R2460 vss.n5216 vss.n327 585
R2461 vss.n5522 vss.n324 585
R2462 vss.n5213 vss.n313 585
R2463 vss.n5526 vss.n310 585
R2464 vss.n5210 vss.n308 585
R2465 vss.n5209 vss.n5208 585
R2466 vss.n1009 vss.n1008 585
R2467 vss.n5201 vss.n1023 585
R2468 vss.n1264 vss.n1021 585
R2469 vss.n5188 vss.n1035 585
R2470 vss.n5364 vss.n843 585
R2471 vss.n955 vss.n834 585
R2472 vss.n5370 vss.n829 585
R2473 vss.n952 vss.n815 585
R2474 vss.n5374 vss.n810 585
R2475 vss.n949 vss.n799 585
R2476 vss.n5380 vss.n794 585
R2477 vss.n946 vss.n782 585
R2478 vss.n5384 vss.n778 585
R2479 vss.n766 vss.n761 585
R2480 vss.n5391 vss.n5390 585
R2481 vss.n5392 vss.n754 585
R2482 vss.n5394 vss.n5393 585
R2483 vss.n5400 vss.n728 585
R2484 vss.n5407 vss.n5406 585
R2485 vss.n5408 vss.n719 585
R2486 vss.n5410 vss.n5409 585
R2487 vss.n705 vss.n700 585
R2488 vss.n5415 vss.n5414 585
R2489 vss.n5416 vss.n691 585
R2490 vss.n5418 vss.n5417 585
R2491 vss.n677 vss.n672 585
R2492 vss.n5423 vss.n5422 585
R2493 vss.n5424 vss.n663 585
R2494 vss.n5426 vss.n5425 585
R2495 vss.n649 vss.n644 585
R2496 vss.n5431 vss.n5430 585
R2497 vss.n5432 vss.n635 585
R2498 vss.n5434 vss.n5433 585
R2499 vss.n621 vss.n616 585
R2500 vss.n5439 vss.n5438 585
R2501 vss.n5440 vss.n607 585
R2502 vss.n5442 vss.n5441 585
R2503 vss.n593 vss.n588 585
R2504 vss.n5447 vss.n5446 585
R2505 vss.n5448 vss.n579 585
R2506 vss.n5450 vss.n5449 585
R2507 vss.n565 vss.n560 585
R2508 vss.n5455 vss.n5454 585
R2509 vss.n5456 vss.n551 585
R2510 vss.n5458 vss.n5457 585
R2511 vss.n537 vss.n532 585
R2512 vss.n5463 vss.n5462 585
R2513 vss.n5464 vss.n523 585
R2514 vss.n5466 vss.n5465 585
R2515 vss.n509 vss.n504 585
R2516 vss.n5471 vss.n5470 585
R2517 vss.n5472 vss.n495 585
R2518 vss.n5474 vss.n5473 585
R2519 vss.n481 vss.n476 585
R2520 vss.n5479 vss.n5478 585
R2521 vss.n5480 vss.n467 585
R2522 vss.n5482 vss.n5481 585
R2523 vss.n453 vss.n448 585
R2524 vss.n5487 vss.n5486 585
R2525 vss.n5488 vss.n439 585
R2526 vss.n5490 vss.n5489 585
R2527 vss.n425 vss.n420 585
R2528 vss.n5495 vss.n5494 585
R2529 vss.n5496 vss.n411 585
R2530 vss.n5498 vss.n5497 585
R2531 vss.n397 vss.n392 585
R2532 vss.n5503 vss.n5502 585
R2533 vss.n5504 vss.n383 585
R2534 vss.n5506 vss.n5505 585
R2535 vss.n369 vss.n364 585
R2536 vss.n5511 vss.n5510 585
R2537 vss.n5512 vss.n355 585
R2538 vss.n5514 vss.n5513 585
R2539 vss.n341 vss.n336 585
R2540 vss.n5519 vss.n5518 585
R2541 vss.n5520 vss.n327 585
R2542 vss.n5522 vss.n5521 585
R2543 vss.n332 vss.n313 585
R2544 vss.n5526 vss.n317 585
R2545 vss.n5195 vss.n308 585
R2546 vss.n5208 vss.n1017 585
R2547 vss.n5199 vss.n1009 585
R2548 vss.n5201 vss.n5200 585
R2549 vss.n1030 vss.n1021 585
R2550 vss.n5189 vss.n5188 585
R2551 vss.n5364 vss.n852 585
R2552 vss.n1121 vss.n834 585
R2553 vss.n5370 vss.n840 585
R2554 vss.n1124 vss.n815 585
R2555 vss.n5374 vss.n820 585
R2556 vss.n1127 vss.n799 585
R2557 vss.n5380 vss.n805 585
R2558 vss.n1130 vss.n782 585
R2559 vss.n5384 vss.n787 585
R2560 vss.n1133 vss.n766 585
R2561 vss.n5390 vss.n771 585
R2562 vss.n1136 vss.n754 585
R2563 vss.n5394 vss.n747 585
R2564 vss.n5402 vss.n741 585
R2565 vss.n5406 vss.n729 585
R2566 vss.n1141 vss.n719 585
R2567 vss.n5410 vss.n715 585
R2568 vss.n1144 vss.n705 585
R2569 vss.n5414 vss.n701 585
R2570 vss.n1147 vss.n691 585
R2571 vss.n5418 vss.n687 585
R2572 vss.n1150 vss.n677 585
R2573 vss.n5422 vss.n673 585
R2574 vss.n1153 vss.n663 585
R2575 vss.n5426 vss.n659 585
R2576 vss.n1156 vss.n649 585
R2577 vss.n5430 vss.n645 585
R2578 vss.n1159 vss.n635 585
R2579 vss.n5434 vss.n631 585
R2580 vss.n1162 vss.n621 585
R2581 vss.n5438 vss.n617 585
R2582 vss.n1165 vss.n607 585
R2583 vss.n5442 vss.n603 585
R2584 vss.n1168 vss.n593 585
R2585 vss.n5446 vss.n589 585
R2586 vss.n1171 vss.n579 585
R2587 vss.n5450 vss.n575 585
R2588 vss.n1174 vss.n565 585
R2589 vss.n5454 vss.n561 585
R2590 vss.n1177 vss.n551 585
R2591 vss.n5458 vss.n547 585
R2592 vss.n1180 vss.n537 585
R2593 vss.n5462 vss.n533 585
R2594 vss.n1183 vss.n523 585
R2595 vss.n5466 vss.n519 585
R2596 vss.n1186 vss.n509 585
R2597 vss.n5470 vss.n505 585
R2598 vss.n1189 vss.n495 585
R2599 vss.n5474 vss.n491 585
R2600 vss.n1192 vss.n481 585
R2601 vss.n5478 vss.n477 585
R2602 vss.n1195 vss.n467 585
R2603 vss.n5482 vss.n463 585
R2604 vss.n1198 vss.n453 585
R2605 vss.n5486 vss.n449 585
R2606 vss.n1201 vss.n439 585
R2607 vss.n5490 vss.n435 585
R2608 vss.n1204 vss.n425 585
R2609 vss.n5494 vss.n421 585
R2610 vss.n1207 vss.n411 585
R2611 vss.n5498 vss.n407 585
R2612 vss.n1210 vss.n397 585
R2613 vss.n5502 vss.n393 585
R2614 vss.n1213 vss.n383 585
R2615 vss.n5506 vss.n379 585
R2616 vss.n1216 vss.n369 585
R2617 vss.n5510 vss.n365 585
R2618 vss.n1219 vss.n355 585
R2619 vss.n5514 vss.n351 585
R2620 vss.n1222 vss.n341 585
R2621 vss.n5518 vss.n337 585
R2622 vss.n1225 vss.n327 585
R2623 vss.n5522 vss.n323 585
R2624 vss.n1228 vss.n313 585
R2625 vss.n5526 vss.n309 585
R2626 vss.n1231 vss.n308 585
R2627 vss.n5208 vss.n1010 585
R2628 vss.n1234 vss.n1009 585
R2629 vss.n5201 vss.n1022 585
R2630 vss.n1237 vss.n1021 585
R2631 vss.n5188 vss.n1034 585
R2632 vss.n5364 vss.n842 585
R2633 vss.n929 vss.n834 585
R2634 vss.n5370 vss.n828 585
R2635 vss.n926 vss.n815 585
R2636 vss.n5374 vss.n809 585
R2637 vss.n923 vss.n799 585
R2638 vss.n5380 vss.n793 585
R2639 vss.n920 vss.n782 585
R2640 vss.n5384 vss.n777 585
R2641 vss.n917 vss.n766 585
R2642 vss.n5390 vss.n762 585
R2643 vss.n914 vss.n754 585
R2644 vss.n5394 vss.n740 585
R2645 vss.n5404 vss.n5403 585
R2646 vss.n5403 vss.n215 585
R2647 vss.n5406 vss.n5405 585
R2648 vss.n719 vss.n714 585
R2649 vss.n5411 vss.n5410 585
R2650 vss.n5412 vss.n705 585
R2651 vss.n5414 vss.n5413 585
R2652 vss.n691 vss.n686 585
R2653 vss.n5419 vss.n5418 585
R2654 vss.n5420 vss.n677 585
R2655 vss.n5422 vss.n5421 585
R2656 vss.n663 vss.n658 585
R2657 vss.n5427 vss.n5426 585
R2658 vss.n5428 vss.n649 585
R2659 vss.n5430 vss.n5429 585
R2660 vss.n635 vss.n630 585
R2661 vss.n5435 vss.n5434 585
R2662 vss.n5436 vss.n621 585
R2663 vss.n5438 vss.n5437 585
R2664 vss.n607 vss.n602 585
R2665 vss.n5443 vss.n5442 585
R2666 vss.n5444 vss.n593 585
R2667 vss.n5446 vss.n5445 585
R2668 vss.n579 vss.n574 585
R2669 vss.n5451 vss.n5450 585
R2670 vss.n5452 vss.n565 585
R2671 vss.n5454 vss.n5453 585
R2672 vss.n551 vss.n546 585
R2673 vss.n5459 vss.n5458 585
R2674 vss.n5460 vss.n537 585
R2675 vss.n5462 vss.n5461 585
R2676 vss.n523 vss.n518 585
R2677 vss.n5467 vss.n5466 585
R2678 vss.n5468 vss.n509 585
R2679 vss.n5470 vss.n5469 585
R2680 vss.n495 vss.n490 585
R2681 vss.n5475 vss.n5474 585
R2682 vss.n5476 vss.n481 585
R2683 vss.n5478 vss.n5477 585
R2684 vss.n467 vss.n462 585
R2685 vss.n5483 vss.n5482 585
R2686 vss.n5484 vss.n453 585
R2687 vss.n5486 vss.n5485 585
R2688 vss.n439 vss.n434 585
R2689 vss.n5491 vss.n5490 585
R2690 vss.n5492 vss.n425 585
R2691 vss.n5494 vss.n5493 585
R2692 vss.n411 vss.n406 585
R2693 vss.n5499 vss.n5498 585
R2694 vss.n5500 vss.n397 585
R2695 vss.n5502 vss.n5501 585
R2696 vss.n383 vss.n378 585
R2697 vss.n5507 vss.n5506 585
R2698 vss.n5508 vss.n369 585
R2699 vss.n5510 vss.n5509 585
R2700 vss.n355 vss.n350 585
R2701 vss.n5515 vss.n5514 585
R2702 vss.n5516 vss.n341 585
R2703 vss.n5518 vss.n5517 585
R2704 vss.n327 vss.n322 585
R2705 vss.n5523 vss.n5522 585
R2706 vss.n5524 vss.n313 585
R2707 vss.n5526 vss.n5525 585
R2708 vss.n318 vss.n308 585
R2709 vss.n5208 vss.n5207 585
R2710 vss.n1018 vss.n1009 585
R2711 vss.n5202 vss.n5201 585
R2712 vss.n1021 vss.n1020 585
R2713 vss.n5188 vss.n5187 585
R2714 vss.n4576 vss.n754 585
R2715 vss.n5390 vss.n772 585
R2716 vss.n788 vss.n766 585
R2717 vss.n5384 vss.n5383 585
R2718 vss.n5382 vss.n782 585
R2719 vss.n5381 vss.n5380 585
R2720 vss.n799 vss.n792 585
R2721 vss.n5374 vss.n5373 585
R2722 vss.n5372 vss.n815 585
R2723 vss.n5371 vss.n5370 585
R2724 vss.n834 vss.n827 585
R2725 vss.n5364 vss.n5363 585
R2726 vss.n2431 vss.n2387 585
R2727 vss.n2431 vss.n2430 585
R2728 vss.n2432 vss.n2381 585
R2729 vss.n2433 vss.n2432 585
R2730 vss.n2376 vss.n2372 585
R2731 vss.n2453 vss.n2372 585
R2732 vss.n2429 vss.n2428 585
R2733 vss.n2430 vss.n2429 585
R2734 vss.n2374 vss.n2373 585
R2735 vss.n2433 vss.n2373 585
R2736 vss.n2452 vss.n2451 585
R2737 vss.n2453 vss.n2452 585
R2738 vss.n5343 vss.n880 585
R2739 vss.n896 vss.n880 585
R2740 vss.n5342 vss.n881 585
R2741 vss.n5341 vss.n879 585
R2742 vss.n5340 vss.n882 585
R2743 vss.n896 vss.n882 585
R2744 vss.n5354 vss.n1004 585
R2745 vss.n5357 vss.n894 585
R2746 vss.n5357 vss.n896 585
R2747 vss.n5360 vss.n868 585
R2748 vss.n867 vss.n847 585
R2749 vss.n896 vss.n847 585
R2750 vss.n5347 vss.n880 585
R2751 vss.n5346 vss.n881 585
R2752 vss.n5345 vss.n879 585
R2753 vss.n5344 vss.n882 585
R2754 vss.n5354 vss.n1003 585
R2755 vss.n5357 vss.n892 585
R2756 vss.n5357 vss.n891 585
R2757 vss.n5360 vss.n865 585
R2758 vss.n864 vss.n847 585
R2759 vss.n891 vss.n847 585
R2760 vss.n898 vss.n880 585
R2761 vss.n4712 vss.n881 585
R2762 vss.n898 vss.n881 585
R2763 vss.n4713 vss.n879 585
R2764 vss.n898 vss.n879 585
R2765 vss.n4714 vss.n882 585
R2766 vss.n898 vss.n882 585
R2767 vss.n5354 vss.n1005 585
R2768 vss.n5357 vss.n897 585
R2769 vss.n5357 vss.n898 585
R2770 vss.n5360 vss.n870 585
R2771 vss.n4719 vss.n847 585
R2772 vss.n898 vss.n847 585
R2773 vss.n887 vss.n880 585
R2774 vss.n4238 vss.n881 585
R2775 vss.n887 vss.n881 585
R2776 vss.n4239 vss.n879 585
R2777 vss.n887 vss.n879 585
R2778 vss.n4240 vss.n882 585
R2779 vss.n887 vss.n882 585
R2780 vss.n5354 vss.n1001 585
R2781 vss.n5357 vss.n888 585
R2782 vss.n5357 vss.n887 585
R2783 vss.n5360 vss.n863 585
R2784 vss.n4245 vss.n847 585
R2785 vss.n887 vss.n847 585
R2786 vss.n900 vss.n880 585
R2787 vss.n4866 vss.n881 585
R2788 vss.n900 vss.n881 585
R2789 vss.n4867 vss.n879 585
R2790 vss.n900 vss.n879 585
R2791 vss.n4868 vss.n882 585
R2792 vss.n900 vss.n882 585
R2793 vss.n5354 vss.n1006 585
R2794 vss.n5357 vss.n899 585
R2795 vss.n5357 vss.n900 585
R2796 vss.n5360 vss.n872 585
R2797 vss.n4873 vss.n847 585
R2798 vss.n900 vss.n847 585
R2799 vss.n885 vss.n880 585
R2800 vss.n996 vss.n881 585
R2801 vss.n885 vss.n881 585
R2802 vss.n997 vss.n879 585
R2803 vss.n885 vss.n879 585
R2804 vss.n998 vss.n882 585
R2805 vss.n885 vss.n882 585
R2806 vss.n5354 vss.n999 585
R2807 vss.n5357 vss.n886 585
R2808 vss.n5357 vss.n885 585
R2809 vss.n5360 vss.n862 585
R2810 vss.n988 vss.n847 585
R2811 vss.n885 vss.n847 585
R2812 vss.n902 vss.n880 585
R2813 vss.n5331 vss.n881 585
R2814 vss.n902 vss.n881 585
R2815 vss.n5332 vss.n879 585
R2816 vss.n902 vss.n879 585
R2817 vss.n5333 vss.n882 585
R2818 vss.n902 vss.n882 585
R2819 vss.n5354 vss.n5334 585
R2820 vss.n5357 vss.n901 585
R2821 vss.n5357 vss.n902 585
R2822 vss.n5360 vss.n874 585
R2823 vss.n5323 vss.n847 585
R2824 vss.n902 vss.n847 585
R2825 vss.n5358 vss.n880 585
R2826 vss.n966 vss.n881 585
R2827 vss.n5358 vss.n881 585
R2828 vss.n967 vss.n879 585
R2829 vss.n5358 vss.n879 585
R2830 vss.n968 vss.n882 585
R2831 vss.n5358 vss.n882 585
R2832 vss.n5354 vss.n969 585
R2833 vss.n5357 vss.n884 585
R2834 vss.n5358 vss.n5357 585
R2835 vss.n5360 vss.n861 585
R2836 vss.n958 vss.n847 585
R2837 vss.n5358 vss.n847 585
R2838 vss.n880 vss.n877 585
R2839 vss.n908 vss.n881 585
R2840 vss.n881 vss.n877 585
R2841 vss.n909 vss.n879 585
R2842 vss.n879 vss.n877 585
R2843 vss.n910 vss.n882 585
R2844 vss.n882 vss.n877 585
R2845 vss.n5355 vss.n5354 585
R2846 vss.n5357 vss.n5356 585
R2847 vss.n5357 vss.n877 585
R2848 vss.n5360 vss.n876 585
R2849 vss.n1118 vss.n847 585
R2850 vss.n877 vss.n847 585
R2851 vss.n911 vss.n880 585
R2852 vss.n940 vss.n881 585
R2853 vss.n911 vss.n881 585
R2854 vss.n941 vss.n879 585
R2855 vss.n911 vss.n879 585
R2856 vss.n942 vss.n882 585
R2857 vss.n911 vss.n882 585
R2858 vss.n5354 vss.n943 585
R2859 vss.n5357 vss.n883 585
R2860 vss.n5360 vss.n860 585
R2861 vss.n932 vss.n847 585
R2862 vss.n911 vss.n847 585
R2863 vss.n5362 vss.n847 585
R2864 vss.n3026 vss.n847 585
R2865 vss.n5361 vss.n5360 585
R2866 vss.n5357 vss.n859 585
R2867 vss.n5354 vss.n5353 585
R2868 vss.n5352 vss.n882 585
R2869 vss.n3026 vss.n882 585
R2870 vss.n5351 vss.n879 585
R2871 vss.n3026 vss.n879 585
R2872 vss.n5350 vss.n881 585
R2873 vss.n3026 vss.n881 585
R2874 vss.n5349 vss.n880 585
R2875 vss.n3026 vss.n880 585
R2876 vss.n6009 vss.n133 585
R2877 vss.n5985 vss.n135 585
R2878 vss.n5986 vss.n141 585
R2879 vss.n5975 vss.n142 585
R2880 vss.n5993 vss.n140 585
R2881 vss.n5994 vss.n143 585
R2882 vss.n5970 vss.n139 585
R2883 vss.n6002 vss.n146 585
R2884 vss.n156 vss.n144 585
R2885 vss.n5962 vss.n158 585
R2886 vss.n5961 vss.n163 585
R2887 vss.n5957 vss.n162 585
R2888 vss.n173 vss.n167 585
R2889 vss.n5950 vss.n175 585
R2890 vss.n5949 vss.n179 585
R2891 vss.n183 vss.n178 585
R2892 vss.n5941 vss.n187 585
R2893 vss.n5940 vss.n190 585
R2894 vss.n194 vss.n189 585
R2895 vss.n5932 vss.n197 585
R2896 vss.n5931 vss.n200 585
R2897 vss.n204 vss.n199 585
R2898 vss.n5923 vss.n207 585
R2899 vss.n5922 vss.n5921 585
R2900 vss.n211 vss.n210 585
R2901 vss.n2764 vss.n2758 585
R2902 vss.n2775 vss.n2757 585
R2903 vss.n2776 vss.n2751 585
R2904 vss.n2748 vss.n2743 585
R2905 vss.n2784 vss.n2742 585
R2906 vss.n2785 vss.n2738 585
R2907 vss.n2732 vss.n2729 585
R2908 vss.n2793 vss.n2728 585
R2909 vss.n2794 vss.n2724 585
R2910 vss.n2718 vss.n2712 585
R2911 vss.n2800 vss.n2711 585
R2912 vss.n2801 vss.n2708 585
R2913 vss.n2702 vss.n2700 585
R2914 vss.n2809 vss.n2699 585
R2915 vss.n2810 vss.n2692 585
R2916 vss.n2689 vss.n2683 585
R2917 vss.n2818 vss.n2682 585
R2918 vss.n2819 vss.n2681 585
R2919 vss.n2672 vss.n2667 585
R2920 vss.n2826 vss.n2666 585
R2921 vss.n2827 vss.n2661 585
R2922 vss.n2828 vss.n2657 585
R2923 vss.n2656 vss.n2648 585
R2924 vss.n2835 vss.n2647 585
R2925 vss.n2836 vss.n2644 585
R2926 vss.n2637 vss.n2635 585
R2927 vss.n2844 vss.n2634 585
R2928 vss.n2845 vss.n2627 585
R2929 vss.n2624 vss.n2619 585
R2930 vss.n2853 vss.n2618 585
R2931 vss.n2854 vss.n2611 585
R2932 vss.n2607 vss.n2604 585
R2933 vss.n2860 vss.n2603 585
R2934 vss.n2861 vss.n2597 585
R2935 vss.n2594 vss.n2589 585
R2936 vss.n2869 vss.n2588 585
R2937 vss.n2870 vss.n2584 585
R2938 vss.n2578 vss.n2575 585
R2939 vss.n2878 vss.n2574 585
R2940 vss.n2879 vss.n2573 585
R2941 vss.n2566 vss.n2560 585
R2942 vss.n2886 vss.n2559 585
R2943 vss.n2887 vss.n2558 585
R2944 vss.n2549 vss.n2547 585
R2945 vss.n2893 vss.n2546 585
R2946 vss.n2894 vss.n2538 585
R2947 vss.n2535 vss.n2532 585
R2948 vss.n2902 vss.n2531 585
R2949 vss.n2903 vss.n2528 585
R2950 vss.n2522 vss.n2517 585
R2951 vss.n2910 vss.n2516 585
R2952 vss.n2911 vss.n2513 585
R2953 vss.n2507 vss.n2501 585
R2954 vss.n2919 vss.n2500 585
R2955 vss.n2920 vss.n2496 585
R2956 vss.n2921 vss.n2493 585
R2957 vss.n2487 vss.n2485 585
R2958 vss.n2929 vss.n2484 585
R2959 vss.n2930 vss.n2477 585
R2960 vss.n2474 vss.n2470 585
R2961 vss.n2938 vss.n2469 585
R2962 vss.n2939 vss.n2466 585
R2963 vss.n2462 vss.n2458 585
R2964 vss.n2947 vss.n2457 585
R2965 vss.n2948 vss.n2365 585
R2966 vss.n2371 vss.n2364 585
R2967 vss.n2363 vss.n2357 585
R2968 vss.n2956 vss.n2356 585
R2969 vss.n2957 vss.n2353 585
R2970 vss.n2352 vss.n2347 585
R2971 vss.n3005 vss.n2346 585
R2972 vss.n2964 vss.n2344 585
R2973 vss.n2997 vss.n2991 585
R2974 vss.n2996 vss.n1329 585
R2975 vss.n4203 vss.n1328 585
R2976 vss.n1335 vss.n1326 585
R2977 vss.n4195 vss.n1337 585
R2978 vss.n4194 vss.n4193 585
R2979 vss.n1342 vss.n1341 585
R2980 vss.n4186 vss.n1350 585
R2981 vss.n4185 vss.n1354 585
R2982 vss.n1353 vss.n1294 585
R2983 vss.n4177 vss.n1361 585
R2984 vss.n4176 vss.n1365 585
R2985 vss.n1369 vss.n1364 585
R2986 vss.n4168 vss.n1373 585
R2987 vss.n4167 vss.n1377 585
R2988 vss.n1381 vss.n1376 585
R2989 vss.n4159 vss.n1385 585
R2990 vss.n4158 vss.n4157 585
R2991 vss.n1389 vss.n1388 585
R2992 vss.n4150 vss.n1397 585
R2993 vss.n4149 vss.n1401 585
R2994 vss.n1405 vss.n1400 585
R2995 vss.n4141 vss.n1409 585
R2996 vss.n4140 vss.n1413 585
R2997 vss.n1417 vss.n1412 585
R2998 vss.n4132 vss.n1421 585
R2999 vss.n4131 vss.n1425 585
R3000 vss.n1429 vss.n1424 585
R3001 vss.n4124 vss.n1445 585
R3002 vss.n4120 vss.n1433 585
R3003 vss.n4119 vss.n1451 585
R3004 vss.n1455 vss.n1450 585
R3005 vss.n4111 vss.n1459 585
R3006 vss.n4110 vss.n1463 585
R3007 vss.n1467 vss.n1462 585
R3008 vss.n4102 vss.n1471 585
R3009 vss.n4101 vss.n1475 585
R3010 vss.n1479 vss.n1474 585
R3011 vss.n4093 vss.n1483 585
R3012 vss.n4092 vss.n4091 585
R3013 vss.n1487 vss.n1486 585
R3014 vss.n4084 vss.n1505 585
R3015 vss.n4083 vss.n1509 585
R3016 vss.n1513 vss.n1508 585
R3017 vss.n4075 vss.n1517 585
R3018 vss.n4074 vss.n1521 585
R3019 vss.n1525 vss.n1520 585
R3020 vss.n4066 vss.n1529 585
R3021 vss.n4065 vss.n1533 585
R3022 vss.n1537 vss.n1532 585
R3023 vss.n4057 vss.n1541 585
R3024 vss.n4056 vss.n4055 585
R3025 vss.n1545 vss.n1544 585
R3026 vss.n4048 vss.n1564 585
R3027 vss.n4047 vss.n1568 585
R3028 vss.n1572 vss.n1567 585
R3029 vss.n4039 vss.n1576 585
R3030 vss.n4038 vss.n1580 585
R3031 vss.n1584 vss.n1579 585
R3032 vss.n4030 vss.n1588 585
R3033 vss.n4029 vss.n1592 585
R3034 vss.n1596 vss.n1591 585
R3035 vss.n4022 vss.n1612 585
R3036 vss.n4018 vss.n1600 585
R3037 vss.n4017 vss.n1618 585
R3038 vss.n1622 vss.n1617 585
R3039 vss.n4009 vss.n1626 585
R3040 vss.n4008 vss.n1630 585
R3041 vss.n1634 vss.n1629 585
R3042 vss.n4000 vss.n1638 585
R3043 vss.n3999 vss.n1642 585
R3044 vss.n1646 vss.n1641 585
R3045 vss.n3991 vss.n1650 585
R3046 vss.n3990 vss.n3989 585
R3047 vss.n1654 vss.n1653 585
R3048 vss.n3982 vss.n1672 585
R3049 vss.n3981 vss.n1676 585
R3050 vss.n1680 vss.n1675 585
R3051 vss.n3973 vss.n1684 585
R3052 vss.n3972 vss.n1688 585
R3053 vss.n1692 vss.n1687 585
R3054 vss.n3964 vss.n1696 585
R3055 vss.n3963 vss.n1700 585
R3056 vss.n1704 vss.n1699 585
R3057 vss.n3955 vss.n1708 585
R3058 vss.n3954 vss.n3953 585
R3059 vss.n1712 vss.n1711 585
R3060 vss.n3946 vss.n1731 585
R3061 vss.n3945 vss.n1735 585
R3062 vss.n1739 vss.n1734 585
R3063 vss.n3937 vss.n1743 585
R3064 vss.n3936 vss.n1747 585
R3065 vss.n1751 vss.n1746 585
R3066 vss.n3928 vss.n1755 585
R3067 vss.n3927 vss.n1759 585
R3068 vss.n1763 vss.n1758 585
R3069 vss.n3920 vss.n1769 585
R3070 vss.n3916 vss.n1767 585
R3071 vss.n3915 vss.n1775 585
R3072 vss.n1779 vss.n1774 585
R3073 vss.n3907 vss.n1783 585
R3074 vss.n3906 vss.n1787 585
R3075 vss.n1791 vss.n1786 585
R3076 vss.n3898 vss.n1795 585
R3077 vss.n3897 vss.n1799 585
R3078 vss.n1803 vss.n1798 585
R3079 vss.n3889 vss.n1807 585
R3080 vss.n3888 vss.n1811 585
R3081 vss.n3884 vss.n1810 585
R3082 vss.n3880 vss.n1815 585
R3083 vss.n3879 vss.n1834 585
R3084 vss.n1838 vss.n1833 585
R3085 vss.n3871 vss.n1842 585
R3086 vss.n3870 vss.n1846 585
R3087 vss.n1850 vss.n1845 585
R3088 vss.n3862 vss.n1854 585
R3089 vss.n3861 vss.n1858 585
R3090 vss.n1862 vss.n1857 585
R3091 vss.n3853 vss.n1866 585
R3092 vss.n3852 vss.n3851 585
R3093 vss.n1870 vss.n1869 585
R3094 vss.n3844 vss.n1888 585
R3095 vss.n3843 vss.n1892 585
R3096 vss.n1896 vss.n1891 585
R3097 vss.n3835 vss.n1900 585
R3098 vss.n3834 vss.n1904 585
R3099 vss.n1908 vss.n1903 585
R3100 vss.n3826 vss.n1912 585
R3101 vss.n3825 vss.n1916 585
R3102 vss.n1920 vss.n1915 585
R3103 vss.n3818 vss.n1936 585
R3104 vss.n3814 vss.n1924 585
R3105 vss.n3813 vss.n1942 585
R3106 vss.n1946 vss.n1941 585
R3107 vss.n3805 vss.n1950 585
R3108 vss.n3804 vss.n1954 585
R3109 vss.n1958 vss.n1953 585
R3110 vss.n3796 vss.n1962 585
R3111 vss.n3795 vss.n1966 585
R3112 vss.n1970 vss.n1965 585
R3113 vss.n3787 vss.n1974 585
R3114 vss.n3786 vss.n1978 585
R3115 vss.n3782 vss.n1977 585
R3116 vss.n3778 vss.n1982 585
R3117 vss.n3777 vss.n2001 585
R3118 vss.n2005 vss.n2000 585
R3119 vss.n3769 vss.n2009 585
R3120 vss.n3768 vss.n2013 585
R3121 vss.n2017 vss.n2012 585
R3122 vss.n3760 vss.n2021 585
R3123 vss.n3759 vss.n2025 585
R3124 vss.n2029 vss.n2024 585
R3125 vss.n3751 vss.n2033 585
R3126 vss.n3750 vss.n3749 585
R3127 vss.n2037 vss.n2036 585
R3128 vss.n3742 vss.n2055 585
R3129 vss.n3741 vss.n2059 585
R3130 vss.n2063 vss.n2058 585
R3131 vss.n3733 vss.n2067 585
R3132 vss.n3732 vss.n2071 585
R3133 vss.n2075 vss.n2070 585
R3134 vss.n3724 vss.n2079 585
R3135 vss.n3723 vss.n2083 585
R3136 vss.n2087 vss.n2082 585
R3137 vss.n3716 vss.n2103 585
R3138 vss.n3712 vss.n2091 585
R3139 vss.n3711 vss.n2109 585
R3140 vss.n2113 vss.n2108 585
R3141 vss.n3703 vss.n2117 585
R3142 vss.n3702 vss.n2121 585
R3143 vss.n2125 vss.n2120 585
R3144 vss.n3694 vss.n2129 585
R3145 vss.n3693 vss.n2133 585
R3146 vss.n2137 vss.n2132 585
R3147 vss.n3685 vss.n2141 585
R3148 vss.n3684 vss.n2145 585
R3149 vss.n3680 vss.n2144 585
R3150 vss.n3676 vss.n2149 585
R3151 vss.n3675 vss.n2157 585
R3152 vss.n2161 vss.n2156 585
R3153 vss.n3667 vss.n2165 585
R3154 vss.n3666 vss.n2169 585
R3155 vss.n2173 vss.n2168 585
R3156 vss.n3658 vss.n2177 585
R3157 vss.n3657 vss.n2181 585
R3158 vss.n2185 vss.n2180 585
R3159 vss.n3649 vss.n2189 585
R3160 vss.n3648 vss.n3647 585
R3161 vss.n2193 vss.n2192 585
R3162 vss.n6009 vss.n131 585
R3163 vss.n5981 vss.n135 585
R3164 vss.n150 vss.n135 585
R3165 vss.n5982 vss.n141 585
R3166 vss.n5978 vss.n142 585
R3167 vss.n5976 vss.n140 585
R3168 vss.n5972 vss.n143 585
R3169 vss.n5968 vss.n139 585
R3170 vss.n6002 vss.n147 585
R3171 vss.n155 vss.n144 585
R3172 vss.n160 vss.n158 585
R3173 vss.n165 vss.n163 585
R3174 vss.n5957 vss.n5956 585
R3175 vss.n5955 vss.n167 585
R3176 vss.n175 vss.n170 585
R3177 vss.n181 vss.n179 585
R3178 vss.n185 vss.n183 585
R3179 vss.n188 vss.n187 585
R3180 vss.n192 vss.n190 585
R3181 vss.n195 vss.n194 585
R3182 vss.n198 vss.n197 585
R3183 vss.n202 vss.n200 585
R3184 vss.n205 vss.n204 585
R3185 vss.n209 vss.n207 585
R3186 vss.n5921 vss.n212 585
R3187 vss.n2767 vss.n211 585
R3188 vss.n2766 vss.n2764 585
R3189 vss.n2759 vss.n2757 585
R3190 vss.n2753 vss.n2751 585
R3191 vss.n2750 vss.n2748 585
R3192 vss.n2744 vss.n2742 585
R3193 vss.n2740 vss.n2738 585
R3194 vss.n2734 vss.n2732 585
R3195 vss.n2730 vss.n2728 585
R3196 vss.n2724 vss.n2722 585
R3197 vss.n2720 vss.n2718 585
R3198 vss.n2713 vss.n2711 585
R3199 vss.n2710 vss.n2708 585
R3200 vss.n2704 vss.n2702 585
R3201 vss.n2701 vss.n2699 585
R3202 vss.n2694 vss.n2692 585
R3203 vss.n2691 vss.n2689 585
R3204 vss.n2684 vss.n2682 585
R3205 vss.n2681 vss.n2676 585
R3206 vss.n2674 vss.n2672 585
R3207 vss.n2669 vss.n2666 585
R3208 vss.n2668 vss.n2661 585
R3209 vss.n2659 vss.n2657 585
R3210 vss.n2656 vss.n2651 585
R3211 vss.n2649 vss.n2647 585
R3212 vss.n2646 vss.n2644 585
R3213 vss.n2639 vss.n2637 585
R3214 vss.n2636 vss.n2634 585
R3215 vss.n2629 vss.n2627 585
R3216 vss.n2626 vss.n2624 585
R3217 vss.n2620 vss.n2618 585
R3218 vss.n2615 vss.n2611 585
R3219 vss.n2614 vss.n2607 585
R3220 vss.n2605 vss.n2603 585
R3221 vss.n2599 vss.n2597 585
R3222 vss.n2596 vss.n2594 585
R3223 vss.n2590 vss.n2588 585
R3224 vss.n2586 vss.n2584 585
R3225 vss.n2580 vss.n2578 585
R3226 vss.n2576 vss.n2574 585
R3227 vss.n2573 vss.n2570 585
R3228 vss.n2568 vss.n2566 585
R3229 vss.n2561 vss.n2559 585
R3230 vss.n2558 vss.n2553 585
R3231 vss.n2551 vss.n2549 585
R3232 vss.n2548 vss.n2546 585
R3233 vss.n2540 vss.n2538 585
R3234 vss.n2537 vss.n2535 585
R3235 vss.n2533 vss.n2531 585
R3236 vss.n2528 vss.n2526 585
R3237 vss.n2524 vss.n2522 585
R3238 vss.n2518 vss.n2516 585
R3239 vss.n2515 vss.n2513 585
R3240 vss.n2509 vss.n2507 585
R3241 vss.n2503 vss.n2500 585
R3242 vss.n2502 vss.n2496 585
R3243 vss.n2495 vss.n2493 585
R3244 vss.n2489 vss.n2487 585
R3245 vss.n2486 vss.n2484 585
R3246 vss.n2479 vss.n2477 585
R3247 vss.n2476 vss.n2474 585
R3248 vss.n2471 vss.n2469 585
R3249 vss.n2468 vss.n2466 585
R3250 vss.n2464 vss.n2462 585
R3251 vss.n2459 vss.n2457 585
R3252 vss.n2368 vss.n2365 585
R3253 vss.n2367 vss.n2364 585
R3254 vss.n2363 vss.n2360 585
R3255 vss.n2358 vss.n2356 585
R3256 vss.n2355 vss.n2353 585
R3257 vss.n2351 vss.n2347 585
R3258 vss.n3005 vss.n2348 585
R3259 vss.n2963 vss.n2344 585
R3260 vss.n2992 vss.n2991 585
R3261 vss.n2994 vss.n1329 585
R3262 vss.n4203 vss.n1330 585
R3263 vss.n1334 vss.n1326 585
R3264 vss.n1339 vss.n1337 585
R3265 vss.n4193 vss.n1344 585
R3266 vss.n1347 vss.n1342 585
R3267 vss.n1352 vss.n1350 585
R3268 vss.n1356 vss.n1354 585
R3269 vss.n1359 vss.n1294 585
R3270 vss.n1363 vss.n1361 585
R3271 vss.n1367 vss.n1365 585
R3272 vss.n1371 vss.n1369 585
R3273 vss.n1375 vss.n1373 585
R3274 vss.n1379 vss.n1377 585
R3275 vss.n1383 vss.n1381 585
R3276 vss.n1387 vss.n1385 585
R3277 vss.n4157 vss.n1391 585
R3278 vss.n1394 vss.n1389 585
R3279 vss.n1399 vss.n1397 585
R3280 vss.n1403 vss.n1401 585
R3281 vss.n1407 vss.n1405 585
R3282 vss.n1411 vss.n1409 585
R3283 vss.n1415 vss.n1413 585
R3284 vss.n1419 vss.n1417 585
R3285 vss.n1423 vss.n1421 585
R3286 vss.n1427 vss.n1425 585
R3287 vss.n1431 vss.n1429 585
R3288 vss.n4124 vss.n4123 585
R3289 vss.n4122 vss.n1433 585
R3290 vss.n1451 vss.n1446 585
R3291 vss.n1457 vss.n1455 585
R3292 vss.n1461 vss.n1459 585
R3293 vss.n1465 vss.n1463 585
R3294 vss.n1469 vss.n1467 585
R3295 vss.n1473 vss.n1471 585
R3296 vss.n1477 vss.n1475 585
R3297 vss.n1481 vss.n1479 585
R3298 vss.n1485 vss.n1483 585
R3299 vss.n4091 vss.n4090 585
R3300 vss.n4089 vss.n1487 585
R3301 vss.n1505 vss.n1500 585
R3302 vss.n1511 vss.n1509 585
R3303 vss.n1515 vss.n1513 585
R3304 vss.n1519 vss.n1517 585
R3305 vss.n1523 vss.n1521 585
R3306 vss.n1527 vss.n1525 585
R3307 vss.n1531 vss.n1529 585
R3308 vss.n1535 vss.n1533 585
R3309 vss.n1539 vss.n1537 585
R3310 vss.n1543 vss.n1541 585
R3311 vss.n4055 vss.n1558 585
R3312 vss.n1561 vss.n1545 585
R3313 vss.n1566 vss.n1564 585
R3314 vss.n1570 vss.n1568 585
R3315 vss.n1574 vss.n1572 585
R3316 vss.n1578 vss.n1576 585
R3317 vss.n1582 vss.n1580 585
R3318 vss.n1586 vss.n1584 585
R3319 vss.n1590 vss.n1588 585
R3320 vss.n1594 vss.n1592 585
R3321 vss.n1598 vss.n1596 585
R3322 vss.n4022 vss.n4021 585
R3323 vss.n4020 vss.n1600 585
R3324 vss.n1618 vss.n1613 585
R3325 vss.n1624 vss.n1622 585
R3326 vss.n1628 vss.n1626 585
R3327 vss.n1632 vss.n1630 585
R3328 vss.n1636 vss.n1634 585
R3329 vss.n1640 vss.n1638 585
R3330 vss.n1644 vss.n1642 585
R3331 vss.n1648 vss.n1646 585
R3332 vss.n1652 vss.n1650 585
R3333 vss.n3989 vss.n3988 585
R3334 vss.n3987 vss.n1654 585
R3335 vss.n1672 vss.n1667 585
R3336 vss.n1678 vss.n1676 585
R3337 vss.n1682 vss.n1680 585
R3338 vss.n1686 vss.n1684 585
R3339 vss.n1690 vss.n1688 585
R3340 vss.n1694 vss.n1692 585
R3341 vss.n1698 vss.n1696 585
R3342 vss.n1702 vss.n1700 585
R3343 vss.n1706 vss.n1704 585
R3344 vss.n1710 vss.n1708 585
R3345 vss.n3953 vss.n1725 585
R3346 vss.n1728 vss.n1712 585
R3347 vss.n1733 vss.n1731 585
R3348 vss.n1737 vss.n1735 585
R3349 vss.n1741 vss.n1739 585
R3350 vss.n1745 vss.n1743 585
R3351 vss.n1749 vss.n1747 585
R3352 vss.n1753 vss.n1751 585
R3353 vss.n1757 vss.n1755 585
R3354 vss.n1761 vss.n1759 585
R3355 vss.n1765 vss.n1763 585
R3356 vss.n3920 vss.n3919 585
R3357 vss.n3918 vss.n1767 585
R3358 vss.n1775 vss.n1770 585
R3359 vss.n1781 vss.n1779 585
R3360 vss.n1785 vss.n1783 585
R3361 vss.n1789 vss.n1787 585
R3362 vss.n1793 vss.n1791 585
R3363 vss.n1797 vss.n1795 585
R3364 vss.n1801 vss.n1799 585
R3365 vss.n1805 vss.n1803 585
R3366 vss.n1809 vss.n1807 585
R3367 vss.n1813 vss.n1811 585
R3368 vss.n3884 vss.n1828 585
R3369 vss.n1831 vss.n1815 585
R3370 vss.n1836 vss.n1834 585
R3371 vss.n1840 vss.n1838 585
R3372 vss.n1844 vss.n1842 585
R3373 vss.n1848 vss.n1846 585
R3374 vss.n1852 vss.n1850 585
R3375 vss.n1856 vss.n1854 585
R3376 vss.n1860 vss.n1858 585
R3377 vss.n1864 vss.n1862 585
R3378 vss.n1868 vss.n1866 585
R3379 vss.n3851 vss.n3850 585
R3380 vss.n3849 vss.n1870 585
R3381 vss.n1888 vss.n1883 585
R3382 vss.n1894 vss.n1892 585
R3383 vss.n1898 vss.n1896 585
R3384 vss.n1902 vss.n1900 585
R3385 vss.n1906 vss.n1904 585
R3386 vss.n1910 vss.n1908 585
R3387 vss.n1914 vss.n1912 585
R3388 vss.n1918 vss.n1916 585
R3389 vss.n1922 vss.n1920 585
R3390 vss.n3818 vss.n3817 585
R3391 vss.n3816 vss.n1924 585
R3392 vss.n1942 vss.n1937 585
R3393 vss.n1948 vss.n1946 585
R3394 vss.n1952 vss.n1950 585
R3395 vss.n1956 vss.n1954 585
R3396 vss.n1960 vss.n1958 585
R3397 vss.n1964 vss.n1962 585
R3398 vss.n1968 vss.n1966 585
R3399 vss.n1972 vss.n1970 585
R3400 vss.n1976 vss.n1974 585
R3401 vss.n1980 vss.n1978 585
R3402 vss.n3782 vss.n1995 585
R3403 vss.n1998 vss.n1982 585
R3404 vss.n2003 vss.n2001 585
R3405 vss.n2007 vss.n2005 585
R3406 vss.n2011 vss.n2009 585
R3407 vss.n2015 vss.n2013 585
R3408 vss.n2019 vss.n2017 585
R3409 vss.n2023 vss.n2021 585
R3410 vss.n2027 vss.n2025 585
R3411 vss.n2031 vss.n2029 585
R3412 vss.n2035 vss.n2033 585
R3413 vss.n3749 vss.n3748 585
R3414 vss.n3747 vss.n2037 585
R3415 vss.n2055 vss.n2050 585
R3416 vss.n2061 vss.n2059 585
R3417 vss.n2065 vss.n2063 585
R3418 vss.n2069 vss.n2067 585
R3419 vss.n2073 vss.n2071 585
R3420 vss.n2077 vss.n2075 585
R3421 vss.n2081 vss.n2079 585
R3422 vss.n2085 vss.n2083 585
R3423 vss.n2089 vss.n2087 585
R3424 vss.n3716 vss.n3715 585
R3425 vss.n3714 vss.n2091 585
R3426 vss.n2109 vss.n2104 585
R3427 vss.n2115 vss.n2113 585
R3428 vss.n2119 vss.n2117 585
R3429 vss.n2123 vss.n2121 585
R3430 vss.n2127 vss.n2125 585
R3431 vss.n2131 vss.n2129 585
R3432 vss.n2135 vss.n2133 585
R3433 vss.n2139 vss.n2137 585
R3434 vss.n2143 vss.n2141 585
R3435 vss.n2147 vss.n2145 585
R3436 vss.n3680 vss.n2151 585
R3437 vss.n2154 vss.n2149 585
R3438 vss.n2159 vss.n2157 585
R3439 vss.n2163 vss.n2161 585
R3440 vss.n2167 vss.n2165 585
R3441 vss.n2171 vss.n2169 585
R3442 vss.n2175 vss.n2173 585
R3443 vss.n2179 vss.n2177 585
R3444 vss.n2183 vss.n2181 585
R3445 vss.n2187 vss.n2185 585
R3446 vss.n2191 vss.n2189 585
R3447 vss.n3647 vss.n3646 585
R3448 vss.n3645 vss.n2193 585
R3449 vss.n3643 vss.n2193 585
R3450 vss.n3647 vss.n3041 585
R3451 vss.n2189 vss.n2184 585
R3452 vss.n3654 vss.n2185 585
R3453 vss.n3655 vss.n2181 585
R3454 vss.n2177 vss.n2172 585
R3455 vss.n3663 vss.n2173 585
R3456 vss.n3664 vss.n2169 585
R3457 vss.n2165 vss.n2160 585
R3458 vss.n3672 vss.n2161 585
R3459 vss.n3673 vss.n2157 585
R3460 vss.n2149 vss.n2148 585
R3461 vss.n3681 vss.n3680 585
R3462 vss.n3682 vss.n2145 585
R3463 vss.n2141 vss.n2136 585
R3464 vss.n3690 vss.n2137 585
R3465 vss.n3691 vss.n2133 585
R3466 vss.n2129 vss.n2124 585
R3467 vss.n3699 vss.n2125 585
R3468 vss.n3700 vss.n2121 585
R3469 vss.n2117 vss.n2112 585
R3470 vss.n3708 vss.n2113 585
R3471 vss.n3709 vss.n2109 585
R3472 vss.n2091 vss.n2090 585
R3473 vss.n3717 vss.n3716 585
R3474 vss.n3718 vss.n2087 585
R3475 vss.n2083 vss.n2078 585
R3476 vss.n3726 vss.n2079 585
R3477 vss.n3727 vss.n2075 585
R3478 vss.n2071 vss.n2066 585
R3479 vss.n3735 vss.n2067 585
R3480 vss.n3736 vss.n2063 585
R3481 vss.n2059 vss.n2054 585
R3482 vss.n3744 vss.n2055 585
R3483 vss.n3745 vss.n2037 585
R3484 vss.n3749 vss.n2049 585
R3485 vss.n2033 vss.n2028 585
R3486 vss.n3756 vss.n2029 585
R3487 vss.n3757 vss.n2025 585
R3488 vss.n2021 vss.n2016 585
R3489 vss.n3765 vss.n2017 585
R3490 vss.n3766 vss.n2013 585
R3491 vss.n2009 vss.n2004 585
R3492 vss.n3774 vss.n2005 585
R3493 vss.n3775 vss.n2001 585
R3494 vss.n1982 vss.n1981 585
R3495 vss.n3783 vss.n3782 585
R3496 vss.n3784 vss.n1978 585
R3497 vss.n1974 vss.n1969 585
R3498 vss.n3792 vss.n1970 585
R3499 vss.n3793 vss.n1966 585
R3500 vss.n1962 vss.n1957 585
R3501 vss.n3801 vss.n1958 585
R3502 vss.n3802 vss.n1954 585
R3503 vss.n1950 vss.n1945 585
R3504 vss.n3810 vss.n1946 585
R3505 vss.n3811 vss.n1942 585
R3506 vss.n1924 vss.n1923 585
R3507 vss.n3819 vss.n3818 585
R3508 vss.n3820 vss.n1920 585
R3509 vss.n1916 vss.n1911 585
R3510 vss.n3828 vss.n1912 585
R3511 vss.n3829 vss.n1908 585
R3512 vss.n1904 vss.n1899 585
R3513 vss.n3837 vss.n1900 585
R3514 vss.n3838 vss.n1896 585
R3515 vss.n1892 vss.n1887 585
R3516 vss.n3846 vss.n1888 585
R3517 vss.n3847 vss.n1870 585
R3518 vss.n3851 vss.n1882 585
R3519 vss.n1866 vss.n1861 585
R3520 vss.n3858 vss.n1862 585
R3521 vss.n3859 vss.n1858 585
R3522 vss.n1854 vss.n1849 585
R3523 vss.n3867 vss.n1850 585
R3524 vss.n3868 vss.n1846 585
R3525 vss.n1842 vss.n1837 585
R3526 vss.n3876 vss.n1838 585
R3527 vss.n3877 vss.n1834 585
R3528 vss.n1815 vss.n1814 585
R3529 vss.n3885 vss.n3884 585
R3530 vss.n3886 vss.n1811 585
R3531 vss.n1807 vss.n1802 585
R3532 vss.n3894 vss.n1803 585
R3533 vss.n3895 vss.n1799 585
R3534 vss.n1795 vss.n1790 585
R3535 vss.n3903 vss.n1791 585
R3536 vss.n3904 vss.n1787 585
R3537 vss.n1783 vss.n1778 585
R3538 vss.n3912 vss.n1779 585
R3539 vss.n3913 vss.n1775 585
R3540 vss.n1767 vss.n1766 585
R3541 vss.n3921 vss.n3920 585
R3542 vss.n3922 vss.n1763 585
R3543 vss.n1759 vss.n1754 585
R3544 vss.n3930 vss.n1755 585
R3545 vss.n3931 vss.n1751 585
R3546 vss.n1747 vss.n1742 585
R3547 vss.n3939 vss.n1743 585
R3548 vss.n3940 vss.n1739 585
R3549 vss.n1735 vss.n1730 585
R3550 vss.n3948 vss.n1731 585
R3551 vss.n3949 vss.n1712 585
R3552 vss.n3953 vss.n1707 585
R3553 vss.n3957 vss.n1708 585
R3554 vss.n3958 vss.n1704 585
R3555 vss.n1700 vss.n1695 585
R3556 vss.n3966 vss.n1696 585
R3557 vss.n3967 vss.n1692 585
R3558 vss.n1688 vss.n1683 585
R3559 vss.n3975 vss.n1684 585
R3560 vss.n3976 vss.n1680 585
R3561 vss.n1676 vss.n1671 585
R3562 vss.n3984 vss.n1672 585
R3563 vss.n3985 vss.n1654 585
R3564 vss.n3989 vss.n1666 585
R3565 vss.n1650 vss.n1645 585
R3566 vss.n3996 vss.n1646 585
R3567 vss.n3997 vss.n1642 585
R3568 vss.n1638 vss.n1633 585
R3569 vss.n4005 vss.n1634 585
R3570 vss.n4006 vss.n1630 585
R3571 vss.n1626 vss.n1621 585
R3572 vss.n4014 vss.n1622 585
R3573 vss.n4015 vss.n1618 585
R3574 vss.n1600 vss.n1599 585
R3575 vss.n4023 vss.n4022 585
R3576 vss.n4024 vss.n1596 585
R3577 vss.n1592 vss.n1587 585
R3578 vss.n4032 vss.n1588 585
R3579 vss.n4033 vss.n1584 585
R3580 vss.n1580 vss.n1575 585
R3581 vss.n4041 vss.n1576 585
R3582 vss.n4042 vss.n1572 585
R3583 vss.n1568 vss.n1563 585
R3584 vss.n4050 vss.n1564 585
R3585 vss.n4051 vss.n1545 585
R3586 vss.n4055 vss.n1540 585
R3587 vss.n4059 vss.n1541 585
R3588 vss.n4060 vss.n1537 585
R3589 vss.n1533 vss.n1528 585
R3590 vss.n4068 vss.n1529 585
R3591 vss.n4069 vss.n1525 585
R3592 vss.n1521 vss.n1516 585
R3593 vss.n4077 vss.n1517 585
R3594 vss.n4078 vss.n1513 585
R3595 vss.n1509 vss.n1504 585
R3596 vss.n4086 vss.n1505 585
R3597 vss.n4087 vss.n1487 585
R3598 vss.n4091 vss.n1499 585
R3599 vss.n1483 vss.n1478 585
R3600 vss.n4098 vss.n1479 585
R3601 vss.n4099 vss.n1475 585
R3602 vss.n1471 vss.n1466 585
R3603 vss.n4107 vss.n1467 585
R3604 vss.n4108 vss.n1463 585
R3605 vss.n1459 vss.n1454 585
R3606 vss.n4116 vss.n1455 585
R3607 vss.n4117 vss.n1451 585
R3608 vss.n1433 vss.n1432 585
R3609 vss.n4125 vss.n4124 585
R3610 vss.n4126 vss.n1429 585
R3611 vss.n1425 vss.n1420 585
R3612 vss.n4134 vss.n1421 585
R3613 vss.n4135 vss.n1417 585
R3614 vss.n1413 vss.n1408 585
R3615 vss.n4143 vss.n1409 585
R3616 vss.n4144 vss.n1405 585
R3617 vss.n1401 vss.n1396 585
R3618 vss.n4152 vss.n1397 585
R3619 vss.n4153 vss.n1389 585
R3620 vss.n4157 vss.n1384 585
R3621 vss.n4161 vss.n1385 585
R3622 vss.n4162 vss.n1381 585
R3623 vss.n1377 vss.n1372 585
R3624 vss.n4170 vss.n1373 585
R3625 vss.n4171 vss.n1369 585
R3626 vss.n1365 vss.n1360 585
R3627 vss.n4179 vss.n1361 585
R3628 vss.n4180 vss.n1294 585
R3629 vss.n1354 vss.n1349 585
R3630 vss.n4188 vss.n1350 585
R3631 vss.n4189 vss.n1342 585
R3632 vss.n4193 vss.n1336 585
R3633 vss.n4197 vss.n1337 585
R3634 vss.n4198 vss.n1326 585
R3635 vss.n4203 vss.n1327 585
R3636 vss.n2965 vss.n1329 585
R3637 vss.n2999 vss.n2991 585
R3638 vss.n3000 vss.n2344 585
R3639 vss.n3005 vss.n2345 585
R3640 vss.n2960 vss.n2347 585
R3641 vss.n2959 vss.n2353 585
R3642 vss.n2356 vss.n2354 585
R3643 vss.n2952 vss.n2363 585
R3644 vss.n2951 vss.n2364 585
R3645 vss.n2950 vss.n2365 585
R3646 vss.n2457 vss.n2366 585
R3647 vss.n2942 vss.n2462 585
R3648 vss.n2941 vss.n2466 585
R3649 vss.n2469 vss.n2467 585
R3650 vss.n2933 vss.n2474 585
R3651 vss.n2932 vss.n2477 585
R3652 vss.n2484 vss.n2478 585
R3653 vss.n2924 vss.n2487 585
R3654 vss.n2923 vss.n2493 585
R3655 vss.n2496 vss.n2494 585
R3656 vss.n2917 vss.n2500 585
R3657 vss.n2916 vss.n2507 585
R3658 vss.n2513 vss.n2508 585
R3659 vss.n2908 vss.n2516 585
R3660 vss.n2907 vss.n2522 585
R3661 vss.n2528 vss.n2523 585
R3662 vss.n2900 vss.n2531 585
R3663 vss.n2899 vss.n2535 585
R3664 vss.n2538 vss.n2536 585
R3665 vss.n2891 vss.n2546 585
R3666 vss.n2890 vss.n2549 585
R3667 vss.n2558 vss.n2550 585
R3668 vss.n2884 vss.n2559 585
R3669 vss.n2883 vss.n2566 585
R3670 vss.n2573 vss.n2567 585
R3671 vss.n2876 vss.n2574 585
R3672 vss.n2875 vss.n2578 585
R3673 vss.n2584 vss.n2579 585
R3674 vss.n2867 vss.n2588 585
R3675 vss.n2866 vss.n2594 585
R3676 vss.n2597 vss.n2595 585
R3677 vss.n2858 vss.n2603 585
R3678 vss.n2857 vss.n2607 585
R3679 vss.n2856 vss.n2611 585
R3680 vss.n2618 vss.n2612 585
R3681 vss.n2848 vss.n2624 585
R3682 vss.n2847 vss.n2627 585
R3683 vss.n2634 vss.n2628 585
R3684 vss.n2839 vss.n2637 585
R3685 vss.n2838 vss.n2644 585
R3686 vss.n2647 vss.n2645 585
R3687 vss.n2831 vss.n2656 585
R3688 vss.n2830 vss.n2657 585
R3689 vss.n2661 vss.n2658 585
R3690 vss.n2824 vss.n2666 585
R3691 vss.n2823 vss.n2672 585
R3692 vss.n2681 vss.n2673 585
R3693 vss.n2816 vss.n2682 585
R3694 vss.n2815 vss.n2689 585
R3695 vss.n2692 vss.n2690 585
R3696 vss.n2807 vss.n2699 585
R3697 vss.n2806 vss.n2702 585
R3698 vss.n2708 vss.n2703 585
R3699 vss.n2798 vss.n2711 585
R3700 vss.n2797 vss.n2718 585
R3701 vss.n2724 vss.n2719 585
R3702 vss.n2791 vss.n2728 585
R3703 vss.n2790 vss.n2732 585
R3704 vss.n2738 vss.n2733 585
R3705 vss.n2782 vss.n2742 585
R3706 vss.n2781 vss.n2748 585
R3707 vss.n2751 vss.n2749 585
R3708 vss.n2773 vss.n2757 585
R3709 vss.n2772 vss.n2764 585
R3710 vss.n2765 vss.n211 585
R3711 vss.n5921 vss.n206 585
R3712 vss.n5925 vss.n207 585
R3713 vss.n5926 vss.n204 585
R3714 vss.n200 vss.n196 585
R3715 vss.n5934 vss.n197 585
R3716 vss.n5935 vss.n194 585
R3717 vss.n190 vss.n186 585
R3718 vss.n5943 vss.n187 585
R3719 vss.n5944 vss.n183 585
R3720 vss.n179 vss.n174 585
R3721 vss.n5952 vss.n175 585
R3722 vss.n5953 vss.n167 585
R3723 vss.n5957 vss.n169 585
R3724 vss.n163 vss.n157 585
R3725 vss.n5964 vss.n158 585
R3726 vss.n5965 vss.n144 585
R3727 vss.n6002 vss.n145 585
R3728 vss.n6002 vss.n136 585
R3729 vss.n5997 vss.n139 585
R3730 vss.n139 vss.n136 585
R3731 vss.n5996 vss.n143 585
R3732 vss.n143 vss.n136 585
R3733 vss.n5971 vss.n140 585
R3734 vss.n140 vss.n136 585
R3735 vss.n5989 vss.n142 585
R3736 vss.n142 vss.n136 585
R3737 vss.n5988 vss.n141 585
R3738 vss.n141 vss.n136 585
R3739 vss.n135 vss.n134 585
R3740 vss.n6010 vss.n6009 585
R3741 vss.n6009 vss.n136 585
R3742 vss.n6009 vss.n132 585
R3743 vss.n6009 vss.n6008 585
R3744 vss.n5983 vss.n135 585
R3745 vss.n5984 vss.n141 585
R3746 vss.n6008 vss.n141 585
R3747 vss.n5979 vss.n142 585
R3748 vss.n6008 vss.n142 585
R3749 vss.n5977 vss.n140 585
R3750 vss.n6008 vss.n140 585
R3751 vss.n5973 vss.n143 585
R3752 vss.n6008 vss.n143 585
R3753 vss.n153 vss.n139 585
R3754 vss.n6008 vss.n139 585
R3755 vss.n6002 vss.n6001 585
R3756 vss.n152 vss.n144 585
R3757 vss.n161 vss.n158 585
R3758 vss.n5959 vss.n163 585
R3759 vss.n5958 vss.n5957 585
R3760 vss.n167 vss.n166 585
R3761 vss.n177 vss.n175 585
R3762 vss.n5947 vss.n179 585
R3763 vss.n5946 vss.n183 585
R3764 vss.n187 vss.n182 585
R3765 vss.n5938 vss.n190 585
R3766 vss.n5937 vss.n194 585
R3767 vss.n197 vss.n193 585
R3768 vss.n5929 vss.n200 585
R3769 vss.n5928 vss.n204 585
R3770 vss.n207 vss.n203 585
R3771 vss.n5921 vss.n213 585
R3772 vss.n2769 vss.n211 585
R3773 vss.n2770 vss.n2764 585
R3774 vss.n2757 vss.n2752 585
R3775 vss.n2778 vss.n2751 585
R3776 vss.n2779 vss.n2748 585
R3777 vss.n2742 vss.n2739 585
R3778 vss.n2787 vss.n2738 585
R3779 vss.n2788 vss.n2732 585
R3780 vss.n2731 vss.n2728 585
R3781 vss.n2724 vss.n2723 585
R3782 vss.n2721 vss.n2718 585
R3783 vss.n2711 vss.n2709 585
R3784 vss.n2803 vss.n2708 585
R3785 vss.n2804 vss.n2702 585
R3786 vss.n2699 vss.n2693 585
R3787 vss.n2812 vss.n2692 585
R3788 vss.n2813 vss.n2689 585
R3789 vss.n2685 vss.n2682 585
R3790 vss.n2681 vss.n2677 585
R3791 vss.n2675 vss.n2672 585
R3792 vss.n2671 vss.n2666 585
R3793 vss.n2670 vss.n2661 585
R3794 vss.n2660 vss.n2657 585
R3795 vss.n2656 vss.n2652 585
R3796 vss.n2650 vss.n2647 585
R3797 vss.n2644 vss.n2638 585
R3798 vss.n2841 vss.n2637 585
R3799 vss.n2842 vss.n2634 585
R3800 vss.n2627 vss.n2625 585
R3801 vss.n2850 vss.n2624 585
R3802 vss.n2851 vss.n2618 585
R3803 vss.n2617 vss.n2611 585
R3804 vss.n2616 vss.n2607 585
R3805 vss.n2603 vss.n2598 585
R3806 vss.n2863 vss.n2597 585
R3807 vss.n2864 vss.n2594 585
R3808 vss.n2588 vss.n2585 585
R3809 vss.n2872 vss.n2584 585
R3810 vss.n2873 vss.n2578 585
R3811 vss.n2577 vss.n2574 585
R3812 vss.n2573 vss.n2571 585
R3813 vss.n2569 vss.n2566 585
R3814 vss.n2562 vss.n2559 585
R3815 vss.n2558 vss.n2554 585
R3816 vss.n2552 vss.n2549 585
R3817 vss.n2546 vss.n2539 585
R3818 vss.n2896 vss.n2538 585
R3819 vss.n2897 vss.n2535 585
R3820 vss.n2534 vss.n2531 585
R3821 vss.n2528 vss.n2527 585
R3822 vss.n2525 vss.n2522 585
R3823 vss.n2516 vss.n2514 585
R3824 vss.n2913 vss.n2513 585
R3825 vss.n2914 vss.n2507 585
R3826 vss.n2505 vss.n2500 585
R3827 vss.n2504 vss.n2496 585
R3828 vss.n2493 vss.n2488 585
R3829 vss.n2926 vss.n2487 585
R3830 vss.n2927 vss.n2484 585
R3831 vss.n2477 vss.n2475 585
R3832 vss.n2935 vss.n2474 585
R3833 vss.n2936 vss.n2469 585
R3834 vss.n2466 vss.n2463 585
R3835 vss.n2944 vss.n2462 585
R3836 vss.n2945 vss.n2457 585
R3837 vss.n2370 vss.n2365 585
R3838 vss.n2369 vss.n2364 585
R3839 vss.n2363 vss.n2361 585
R3840 vss.n2359 vss.n2356 585
R3841 vss.n2353 vss.n2350 585
R3842 vss.n2962 vss.n2347 585
R3843 vss.n3005 vss.n3004 585
R3844 vss.n2349 vss.n2344 585
R3845 vss.n2993 vss.n2991 585
R3846 vss.n1332 vss.n1329 585
R3847 vss.n4203 vss.n4202 585
R3848 vss.n1331 vss.n1326 585
R3849 vss.n1340 vss.n1337 585
R3850 vss.n4193 vss.n4192 585
R3851 vss.n4191 vss.n1342 585
R3852 vss.n1350 vss.n1345 585
R3853 vss.n4183 vss.n1354 585
R3854 vss.n4182 vss.n1294 585
R3855 vss.n1361 vss.n1357 585
R3856 vss.n4174 vss.n1365 585
R3857 vss.n4173 vss.n1369 585
R3858 vss.n1373 vss.n1368 585
R3859 vss.n4165 vss.n1377 585
R3860 vss.n4164 vss.n1381 585
R3861 vss.n1385 vss.n1380 585
R3862 vss.n4157 vss.n4156 585
R3863 vss.n4155 vss.n1389 585
R3864 vss.n1397 vss.n1392 585
R3865 vss.n4147 vss.n1401 585
R3866 vss.n4146 vss.n1405 585
R3867 vss.n1409 vss.n1404 585
R3868 vss.n4138 vss.n1413 585
R3869 vss.n4137 vss.n1417 585
R3870 vss.n1421 vss.n1416 585
R3871 vss.n4129 vss.n1425 585
R3872 vss.n4128 vss.n1429 585
R3873 vss.n4124 vss.n1428 585
R3874 vss.n1448 vss.n1433 585
R3875 vss.n1453 vss.n1451 585
R3876 vss.n4114 vss.n1455 585
R3877 vss.n4113 vss.n1459 585
R3878 vss.n1463 vss.n1458 585
R3879 vss.n4105 vss.n1467 585
R3880 vss.n4104 vss.n1471 585
R3881 vss.n1475 vss.n1470 585
R3882 vss.n4096 vss.n1479 585
R3883 vss.n4095 vss.n1483 585
R3884 vss.n4091 vss.n1482 585
R3885 vss.n1502 vss.n1487 585
R3886 vss.n1507 vss.n1505 585
R3887 vss.n4081 vss.n1509 585
R3888 vss.n4080 vss.n1513 585
R3889 vss.n1517 vss.n1512 585
R3890 vss.n4072 vss.n1521 585
R3891 vss.n4071 vss.n1525 585
R3892 vss.n1529 vss.n1524 585
R3893 vss.n4063 vss.n1533 585
R3894 vss.n4062 vss.n1537 585
R3895 vss.n1541 vss.n1536 585
R3896 vss.n4055 vss.n4054 585
R3897 vss.n4053 vss.n1545 585
R3898 vss.n1564 vss.n1559 585
R3899 vss.n4045 vss.n1568 585
R3900 vss.n4044 vss.n1572 585
R3901 vss.n1576 vss.n1571 585
R3902 vss.n4036 vss.n1580 585
R3903 vss.n4035 vss.n1584 585
R3904 vss.n1588 vss.n1583 585
R3905 vss.n4027 vss.n1592 585
R3906 vss.n4026 vss.n1596 585
R3907 vss.n4022 vss.n1595 585
R3908 vss.n1615 vss.n1600 585
R3909 vss.n1620 vss.n1618 585
R3910 vss.n4012 vss.n1622 585
R3911 vss.n4011 vss.n1626 585
R3912 vss.n1630 vss.n1625 585
R3913 vss.n4003 vss.n1634 585
R3914 vss.n4002 vss.n1638 585
R3915 vss.n1642 vss.n1637 585
R3916 vss.n3994 vss.n1646 585
R3917 vss.n3993 vss.n1650 585
R3918 vss.n3989 vss.n1649 585
R3919 vss.n1669 vss.n1654 585
R3920 vss.n1674 vss.n1672 585
R3921 vss.n3979 vss.n1676 585
R3922 vss.n3978 vss.n1680 585
R3923 vss.n1684 vss.n1679 585
R3924 vss.n3970 vss.n1688 585
R3925 vss.n3969 vss.n1692 585
R3926 vss.n1696 vss.n1691 585
R3927 vss.n3961 vss.n1700 585
R3928 vss.n3960 vss.n1704 585
R3929 vss.n1708 vss.n1703 585
R3930 vss.n3953 vss.n3952 585
R3931 vss.n3951 vss.n1712 585
R3932 vss.n1731 vss.n1726 585
R3933 vss.n3943 vss.n1735 585
R3934 vss.n3942 vss.n1739 585
R3935 vss.n1743 vss.n1738 585
R3936 vss.n3934 vss.n1747 585
R3937 vss.n3933 vss.n1751 585
R3938 vss.n1755 vss.n1750 585
R3939 vss.n3925 vss.n1759 585
R3940 vss.n3924 vss.n1763 585
R3941 vss.n3920 vss.n1762 585
R3942 vss.n1772 vss.n1767 585
R3943 vss.n1777 vss.n1775 585
R3944 vss.n3910 vss.n1779 585
R3945 vss.n3909 vss.n1783 585
R3946 vss.n1787 vss.n1782 585
R3947 vss.n3901 vss.n1791 585
R3948 vss.n3900 vss.n1795 585
R3949 vss.n1799 vss.n1794 585
R3950 vss.n3892 vss.n1803 585
R3951 vss.n3891 vss.n1807 585
R3952 vss.n1811 vss.n1806 585
R3953 vss.n3884 vss.n3883 585
R3954 vss.n3882 vss.n1815 585
R3955 vss.n1834 vss.n1829 585
R3956 vss.n3874 vss.n1838 585
R3957 vss.n3873 vss.n1842 585
R3958 vss.n1846 vss.n1841 585
R3959 vss.n3865 vss.n1850 585
R3960 vss.n3864 vss.n1854 585
R3961 vss.n1858 vss.n1853 585
R3962 vss.n3856 vss.n1862 585
R3963 vss.n3855 vss.n1866 585
R3964 vss.n3851 vss.n1865 585
R3965 vss.n1885 vss.n1870 585
R3966 vss.n1890 vss.n1888 585
R3967 vss.n3841 vss.n1892 585
R3968 vss.n3840 vss.n1896 585
R3969 vss.n1900 vss.n1895 585
R3970 vss.n3832 vss.n1904 585
R3971 vss.n3831 vss.n1908 585
R3972 vss.n1912 vss.n1907 585
R3973 vss.n3823 vss.n1916 585
R3974 vss.n3822 vss.n1920 585
R3975 vss.n3818 vss.n1919 585
R3976 vss.n1939 vss.n1924 585
R3977 vss.n1944 vss.n1942 585
R3978 vss.n3808 vss.n1946 585
R3979 vss.n3807 vss.n1950 585
R3980 vss.n1954 vss.n1949 585
R3981 vss.n3799 vss.n1958 585
R3982 vss.n3798 vss.n1962 585
R3983 vss.n1966 vss.n1961 585
R3984 vss.n3790 vss.n1970 585
R3985 vss.n3789 vss.n1974 585
R3986 vss.n1978 vss.n1973 585
R3987 vss.n3782 vss.n3781 585
R3988 vss.n3780 vss.n1982 585
R3989 vss.n2001 vss.n1996 585
R3990 vss.n3772 vss.n2005 585
R3991 vss.n3771 vss.n2009 585
R3992 vss.n2013 vss.n2008 585
R3993 vss.n3763 vss.n2017 585
R3994 vss.n3762 vss.n2021 585
R3995 vss.n2025 vss.n2020 585
R3996 vss.n3754 vss.n2029 585
R3997 vss.n3753 vss.n2033 585
R3998 vss.n3749 vss.n2032 585
R3999 vss.n2052 vss.n2037 585
R4000 vss.n2057 vss.n2055 585
R4001 vss.n3739 vss.n2059 585
R4002 vss.n3738 vss.n2063 585
R4003 vss.n2067 vss.n2062 585
R4004 vss.n3730 vss.n2071 585
R4005 vss.n3729 vss.n2075 585
R4006 vss.n2079 vss.n2074 585
R4007 vss.n3721 vss.n2083 585
R4008 vss.n3720 vss.n2087 585
R4009 vss.n3716 vss.n2086 585
R4010 vss.n2106 vss.n2091 585
R4011 vss.n2111 vss.n2109 585
R4012 vss.n3706 vss.n2113 585
R4013 vss.n3705 vss.n2117 585
R4014 vss.n2121 vss.n2116 585
R4015 vss.n3697 vss.n2125 585
R4016 vss.n3696 vss.n2129 585
R4017 vss.n2133 vss.n2128 585
R4018 vss.n3688 vss.n2137 585
R4019 vss.n3687 vss.n2141 585
R4020 vss.n2145 vss.n2140 585
R4021 vss.n3680 vss.n3679 585
R4022 vss.n3678 vss.n2149 585
R4023 vss.n2157 vss.n2152 585
R4024 vss.n3670 vss.n2161 585
R4025 vss.n3669 vss.n2165 585
R4026 vss.n2169 vss.n2164 585
R4027 vss.n3661 vss.n2173 585
R4028 vss.n3660 vss.n2177 585
R4029 vss.n2181 vss.n2176 585
R4030 vss.n3652 vss.n2185 585
R4031 vss.n3651 vss.n2189 585
R4032 vss.n3647 vss.n2188 585
R4033 vss.n3044 vss.n2193 585
R4034 vss.n2287 vss.n2228 475.118
R4035 vss.n2308 vss.n1295 475.118
R4036 vss.n4232 vss.n1296 475.118
R4037 vss.n4228 vss.n1302 475.118
R4038 vss.n3023 vss.n1321 475.118
R4039 vss.n4207 vss.n1322 475.118
R4040 vss.n2988 vss.n2340 475.118
R4041 vss.n3008 vss.n2341 475.118
R4042 vss.n2420 vss.n2389 475.118
R4043 vss.n2429 vss.n2373 475.118
R4044 vss.n2285 vss.n2215 475.118
R4045 vss.n2311 vss.n2310 475.118
R4046 vss.n2212 vss.n1292 475.118
R4047 vss.n2195 vss.n1304 475.118
R4048 vss.n2199 vss.n2196 475.118
R4049 vss.n2980 vss.n1324 475.118
R4050 vss.n2982 vss.n2967 475.118
R4051 vss.n2394 vss.n2342 475.118
R4052 vss.n2422 vss.n2386 475.118
R4053 vss.n2432 vss.n2431 475.118
R4054 vss.n2287 vss.n2246 417.176
R4055 vss.n2308 vss.n2228 417.176
R4056 vss.n4232 vss.n1295 417.176
R4057 vss.n4228 vss.n1296 417.176
R4058 vss.n3023 vss.n1302 417.176
R4059 vss.n4207 vss.n1321 417.176
R4060 vss.n2988 vss.n1322 417.176
R4061 vss.n3008 vss.n2340 417.176
R4062 vss.n2420 vss.n2341 417.176
R4063 vss.n2429 vss.n2389 417.176
R4064 vss.n2452 vss.n2373 417.176
R4065 vss.n2285 vss.n2284 417.176
R4066 vss.n2310 vss.n2215 417.176
R4067 vss.n2311 vss.n1292 417.176
R4068 vss.n2212 vss.n1304 417.176
R4069 vss.n2196 vss.n2195 417.176
R4070 vss.n2199 vss.n1324 417.176
R4071 vss.n2980 vss.n2967 417.176
R4072 vss.n2982 vss.n2342 417.176
R4073 vss.n2422 vss.n2394 417.176
R4074 vss.n2431 vss.n2386 417.176
R4075 vss.n2432 vss.n2372 417.176
R4076 vss.n5916 vss.n5915 376.094
R4077 vss.n5917 vss.n5916 376.094
R4078 vss.n5918 vss.n218 322.55
R4079 vss.n5665 vss.n219 319.625
R4080 vss.n5916 vss.n219 319.625
R4081 vss.n5579 vss.n220 319.625
R4082 vss.n2413 vss.n2412 292.5
R4083 vss.t42 vss.n2413 292.5
R4084 vss.n3014 vss.n3013 292.5
R4085 vss.t41 vss.n3014 292.5
R4086 vss.n2201 vss.n1314 292.5
R4087 vss.t283 vss.n2201 292.5
R4088 vss.n2322 vss.n2321 292.5
R4089 vss.t7 vss.n2322 292.5
R4090 vss.n2302 vss.n2301 292.5
R4091 vss.n2301 vss.t284 292.5
R4092 vss.n2300 vss.n2299 292.5
R4093 vss.t284 vss.n2300 292.5
R4094 vss.n2324 vss.n2323 292.5
R4095 vss.n2323 vss.t7 292.5
R4096 vss.n3019 vss.n3018 292.5
R4097 vss.t283 vss.n3019 292.5
R4098 vss.n3016 vss.n3015 292.5
R4099 vss.n3015 vss.t41 292.5
R4100 vss.n2416 vss.n2415 292.5
R4101 vss.t42 vss.n2416 292.5
R4102 vss.n2447 vss.n305 292.5
R4103 vss.t4 vss.n305 292.5
R4104 vss.n304 vss.n303 292.5
R4105 vss.t4 vss.n304 292.5
R4106 vss.n891 vss.n890 288.024
R4107 vss.n891 vss.n889 288.024
R4108 vss.n3026 vss.n893 288.024
R4109 vss.n896 vss.n895 287.413
R4110 vss.n911 vss.n866 287.413
R4111 vss.n6006 vss.n6005 278.925
R4112 vss.n6006 vss.n6004 278.925
R4113 vss.n6006 vss.n6003 278.925
R4114 vss.n150 vss.n149 278.925
R4115 vss.n150 vss.n148 278.925
R4116 vss.n151 vss.n150 278.925
R4117 vss.n4742 vss.n4588 275.058
R4118 vss.n4898 vss.n4742 275.058
R4119 vss.n5400 vss.n5399 275.058
R4120 vss.n5403 vss.n5402 275.058
R4121 vss.n5360 vss.n869 264.132
R4122 vss.n5354 vss.n1002 264.132
R4123 vss.n5360 vss.n871 264.132
R4124 vss.n5354 vss.n1000 264.132
R4125 vss.n5360 vss.n873 264.132
R4126 vss.n5354 vss.n970 264.132
R4127 vss.n5360 vss.n875 264.132
R4128 vss.n5354 vss.n878 264.132
R4129 vss.n5360 vss.n5359 264.132
R4130 vss.n5354 vss.n912 264.132
R4131 vss.n6009 vss.n137 264.132
R4132 vss.n6007 vss.n6002 264.132
R4133 vss.n138 vss.n135 264.132
R4134 vss.n911 vss.n136 239.445
R4135 vss.n4587 vss.n215 236.826
R4136 vss.n4897 vss.n215 236.826
R4137 vss.n5398 vss.n215 236.826
R4138 vss.n5401 vss.n215 236.826
R4139 vss.n3029 vss.n2193 146.25
R4140 vss.n3647 vss.n3040 146.25
R4141 vss.n3039 vss.n2189 146.25
R4142 vss.n3038 vss.n2185 146.25
R4143 vss.n3037 vss.n2181 146.25
R4144 vss.n3036 vss.n2177 146.25
R4145 vss.n3035 vss.n2173 146.25
R4146 vss.n3034 vss.n2169 146.25
R4147 vss.n3033 vss.n2165 146.25
R4148 vss.n3032 vss.n2161 146.25
R4149 vss.n3031 vss.n2157 146.25
R4150 vss.n3030 vss.n2149 146.25
R4151 vss.n3680 vss.n2150 146.25
R4152 vss.n2263 vss.n2145 146.25
R4153 vss.n2264 vss.n2141 146.25
R4154 vss.n2265 vss.n2137 146.25
R4155 vss.n2266 vss.n2133 146.25
R4156 vss.n2267 vss.n2129 146.25
R4157 vss.n2268 vss.n2125 146.25
R4158 vss.n2273 vss.n2121 146.25
R4159 vss.n2272 vss.n2117 146.25
R4160 vss.n2271 vss.n2113 146.25
R4161 vss.n2270 vss.n2109 146.25
R4162 vss.n2269 vss.n2091 146.25
R4163 vss.n3716 vss.n2102 146.25
R4164 vss.n2101 vss.n2087 146.25
R4165 vss.n2100 vss.n2083 146.25
R4166 vss.n2099 vss.n2079 146.25
R4167 vss.n2098 vss.n2075 146.25
R4168 vss.n2097 vss.n2071 146.25
R4169 vss.n2096 vss.n2067 146.25
R4170 vss.n2095 vss.n2063 146.25
R4171 vss.n2094 vss.n2059 146.25
R4172 vss.n2093 vss.n2055 146.25
R4173 vss.n2092 vss.n2037 146.25
R4174 vss.n3749 vss.n2048 146.25
R4175 vss.n2047 vss.n2033 146.25
R4176 vss.n2046 vss.n2029 146.25
R4177 vss.n2045 vss.n2025 146.25
R4178 vss.n2044 vss.n2021 146.25
R4179 vss.n2043 vss.n2017 146.25
R4180 vss.n2042 vss.n2013 146.25
R4181 vss.n2041 vss.n2009 146.25
R4182 vss.n2040 vss.n2005 146.25
R4183 vss.n2039 vss.n2001 146.25
R4184 vss.n2038 vss.n1982 146.25
R4185 vss.n3782 vss.n1994 146.25
R4186 vss.n1993 vss.n1978 146.25
R4187 vss.n1992 vss.n1974 146.25
R4188 vss.n1991 vss.n1970 146.25
R4189 vss.n1990 vss.n1966 146.25
R4190 vss.n1989 vss.n1962 146.25
R4191 vss.n1988 vss.n1958 146.25
R4192 vss.n1987 vss.n1954 146.25
R4193 vss.n1986 vss.n1950 146.25
R4194 vss.n1985 vss.n1946 146.25
R4195 vss.n1984 vss.n1942 146.25
R4196 vss.n1983 vss.n1924 146.25
R4197 vss.n3818 vss.n1935 146.25
R4198 vss.n1934 vss.n1920 146.25
R4199 vss.n1933 vss.n1916 146.25
R4200 vss.n1932 vss.n1912 146.25
R4201 vss.n1931 vss.n1908 146.25
R4202 vss.n1930 vss.n1904 146.25
R4203 vss.n1929 vss.n1900 146.25
R4204 vss.n1928 vss.n1896 146.25
R4205 vss.n1927 vss.n1892 146.25
R4206 vss.n1926 vss.n1888 146.25
R4207 vss.n1925 vss.n1870 146.25
R4208 vss.n3851 vss.n1881 146.25
R4209 vss.n1880 vss.n1866 146.25
R4210 vss.n1879 vss.n1862 146.25
R4211 vss.n1878 vss.n1858 146.25
R4212 vss.n1877 vss.n1854 146.25
R4213 vss.n1876 vss.n1850 146.25
R4214 vss.n1875 vss.n1846 146.25
R4215 vss.n1874 vss.n1842 146.25
R4216 vss.n1873 vss.n1838 146.25
R4217 vss.n1872 vss.n1834 146.25
R4218 vss.n1871 vss.n1815 146.25
R4219 vss.n3884 vss.n1827 146.25
R4220 vss.n1826 vss.n1811 146.25
R4221 vss.n1825 vss.n1807 146.25
R4222 vss.n1824 vss.n1803 146.25
R4223 vss.n1823 vss.n1799 146.25
R4224 vss.n1822 vss.n1795 146.25
R4225 vss.n1821 vss.n1791 146.25
R4226 vss.n1820 vss.n1787 146.25
R4227 vss.n1819 vss.n1783 146.25
R4228 vss.n1818 vss.n1779 146.25
R4229 vss.n1817 vss.n1775 146.25
R4230 vss.n1816 vss.n1767 146.25
R4231 vss.n3920 vss.n1768 146.25
R4232 vss.n2251 vss.n1763 146.25
R4233 vss.n2252 vss.n1759 146.25
R4234 vss.n2253 vss.n1755 146.25
R4235 vss.n2260 vss.n1751 146.25
R4236 vss.n2259 vss.n1747 146.25
R4237 vss.n2258 vss.n1743 146.25
R4238 vss.n2257 vss.n1739 146.25
R4239 vss.n2256 vss.n1735 146.25
R4240 vss.n2255 vss.n1731 146.25
R4241 vss.n2254 vss.n1712 146.25
R4242 vss.n3953 vss.n1724 146.25
R4243 vss.n1723 vss.n1708 146.25
R4244 vss.n1722 vss.n1704 146.25
R4245 vss.n1721 vss.n1700 146.25
R4246 vss.n1720 vss.n1696 146.25
R4247 vss.n1719 vss.n1692 146.25
R4248 vss.n1718 vss.n1688 146.25
R4249 vss.n1717 vss.n1684 146.25
R4250 vss.n1716 vss.n1680 146.25
R4251 vss.n1715 vss.n1676 146.25
R4252 vss.n1714 vss.n1672 146.25
R4253 vss.n1713 vss.n1654 146.25
R4254 vss.n3989 vss.n1665 146.25
R4255 vss.n1664 vss.n1650 146.25
R4256 vss.n1663 vss.n1646 146.25
R4257 vss.n1662 vss.n1642 146.25
R4258 vss.n1661 vss.n1638 146.25
R4259 vss.n1660 vss.n1634 146.25
R4260 vss.n1659 vss.n1630 146.25
R4261 vss.n1658 vss.n1626 146.25
R4262 vss.n1657 vss.n1622 146.25
R4263 vss.n1656 vss.n1618 146.25
R4264 vss.n1655 vss.n1600 146.25
R4265 vss.n4022 vss.n1611 146.25
R4266 vss.n1610 vss.n1596 146.25
R4267 vss.n1609 vss.n1592 146.25
R4268 vss.n1608 vss.n1588 146.25
R4269 vss.n1607 vss.n1584 146.25
R4270 vss.n1606 vss.n1580 146.25
R4271 vss.n1605 vss.n1576 146.25
R4272 vss.n1604 vss.n1572 146.25
R4273 vss.n1603 vss.n1568 146.25
R4274 vss.n1602 vss.n1564 146.25
R4275 vss.n1601 vss.n1545 146.25
R4276 vss.n4055 vss.n1557 146.25
R4277 vss.n1556 vss.n1541 146.25
R4278 vss.n1555 vss.n1537 146.25
R4279 vss.n1554 vss.n1533 146.25
R4280 vss.n1553 vss.n1529 146.25
R4281 vss.n1552 vss.n1525 146.25
R4282 vss.n1551 vss.n1521 146.25
R4283 vss.n1550 vss.n1517 146.25
R4284 vss.n1549 vss.n1513 146.25
R4285 vss.n1548 vss.n1509 146.25
R4286 vss.n1547 vss.n1505 146.25
R4287 vss.n1546 vss.n1487 146.25
R4288 vss.n4091 vss.n1498 146.25
R4289 vss.n1497 vss.n1483 146.25
R4290 vss.n1496 vss.n1479 146.25
R4291 vss.n1495 vss.n1475 146.25
R4292 vss.n1494 vss.n1471 146.25
R4293 vss.n1493 vss.n1467 146.25
R4294 vss.n1492 vss.n1463 146.25
R4295 vss.n1491 vss.n1459 146.25
R4296 vss.n1490 vss.n1455 146.25
R4297 vss.n1489 vss.n1451 146.25
R4298 vss.n1488 vss.n1433 146.25
R4299 vss.n4124 vss.n1444 146.25
R4300 vss.n1443 vss.n1429 146.25
R4301 vss.n1442 vss.n1425 146.25
R4302 vss.n1441 vss.n1421 146.25
R4303 vss.n1440 vss.n1417 146.25
R4304 vss.n1439 vss.n1413 146.25
R4305 vss.n1438 vss.n1409 146.25
R4306 vss.n1437 vss.n1405 146.25
R4307 vss.n1436 vss.n1401 146.25
R4308 vss.n1435 vss.n1397 146.25
R4309 vss.n1434 vss.n1389 146.25
R4310 vss.n4157 vss.n1390 146.25
R4311 vss.n2249 vss.n1385 146.25
R4312 vss.n2281 vss.n1381 146.25
R4313 vss.n2247 vss.n1377 146.25
R4314 vss.n2233 vss.n1373 146.25
R4315 vss.n2216 vss.n1369 146.25
R4316 vss.n2227 vss.n1365 146.25
R4317 vss.n2217 vss.n1361 146.25
R4318 vss.n4233 vss.n1294 146.25
R4319 vss.n2205 vss.n1354 146.25
R4320 vss.n1350 vss.n1303 146.25
R4321 vss.n1342 vss.n1305 146.25
R4322 vss.n4193 vss.n1343 146.25
R4323 vss.n3020 vss.n1337 146.25
R4324 vss.n1326 vss.n1323 146.25
R4325 vss.n4204 vss.n4203 146.25
R4326 vss.n2966 vss.n1329 146.25
R4327 vss.n2991 vss.n2990 146.25
R4328 vss.n3006 vss.n3005 146.25
R4329 vss.n2399 vss.n2347 146.25
R4330 vss.n2419 vss.n2353 146.25
R4331 vss.n2395 vss.n2356 146.25
R4332 vss.n2388 vss.n2363 146.25
R4333 vss.n2434 vss.n2364 146.25
R4334 vss.n2454 vss.n2365 146.25
R4335 vss.n2457 vss.n2456 146.25
R4336 vss.n2462 vss.n2461 146.25
R4337 vss.n2466 vss.n306 146.25
R4338 vss.n2469 vss.n307 146.25
R4339 vss.n2474 vss.n2473 146.25
R4340 vss.n2481 vss.n2477 146.25
R4341 vss.n2484 vss.n2483 146.25
R4342 vss.n2490 vss.n2487 146.25
R4343 vss.n2493 vss.n2492 146.25
R4344 vss.n2497 vss.n2496 146.25
R4345 vss.n2500 vss.n2499 146.25
R4346 vss.n2513 vss.n2512 146.25
R4347 vss.n2519 vss.n2516 146.25
R4348 vss.n2522 vss.n2521 146.25
R4349 vss.n2529 vss.n2528 146.25
R4350 vss.n2542 vss.n2535 146.25
R4351 vss.n2543 vss.n2538 146.25
R4352 vss.n2546 vss.n2545 146.25
R4353 vss.n2555 vss.n2549 146.25
R4354 vss.n2558 vss.n2557 146.25
R4355 vss.n2563 vss.n2559 146.25
R4356 vss.n2566 vss.n2565 146.25
R4357 vss.n2573 vss.n2572 146.25
R4358 vss.n2574 vss.n224 146.25
R4359 vss.n2581 vss.n2578 146.25
R4360 vss.n2584 vss.n2583 146.25
R4361 vss.n2591 vss.n2588 146.25
R4362 vss.n2594 vss.n2593 146.25
R4363 vss.n2600 vss.n2597 146.25
R4364 vss.n2603 vss.n2602 146.25
R4365 vss.n2608 vss.n2607 146.25
R4366 vss.n2611 vss.n2610 146.25
R4367 vss.n2621 vss.n2618 146.25
R4368 vss.n2624 vss.n2623 146.25
R4369 vss.n2631 vss.n2627 146.25
R4370 vss.n2634 vss.n2633 146.25
R4371 vss.n2644 vss.n2643 146.25
R4372 vss.n2653 vss.n2647 146.25
R4373 vss.n2656 vss.n2655 146.25
R4374 vss.n2662 vss.n2657 146.25
R4375 vss.n2663 vss.n2661 146.25
R4376 vss.n2666 vss.n2665 146.25
R4377 vss.n2678 vss.n2672 146.25
R4378 vss.n2681 vss.n2680 146.25
R4379 vss.n2686 vss.n2682 146.25
R4380 vss.n2689 vss.n2688 146.25
R4381 vss.n2696 vss.n2692 146.25
R4382 vss.n2699 vss.n2698 146.25
R4383 vss.n2705 vss.n2702 146.25
R4384 vss.n2708 vss.n2707 146.25
R4385 vss.n2715 vss.n2711 146.25
R4386 vss.n2718 vss.n2717 146.25
R4387 vss.n2725 vss.n2724 146.25
R4388 vss.n2728 vss.n2727 146.25
R4389 vss.n2735 vss.n2732 146.25
R4390 vss.n2738 vss.n2737 146.25
R4391 vss.n2745 vss.n2742 146.25
R4392 vss.n2748 vss.n2747 146.25
R4393 vss.n2754 vss.n2751 146.25
R4394 vss.n2757 vss.n2756 146.25
R4395 vss.n2764 vss.n2763 146.25
R4396 vss.n2761 vss.n211 146.25
R4397 vss.n751 vss.n207 146.25
R4398 vss.n773 vss.n204 146.25
R4399 vss.n774 vss.n200 146.25
R4400 vss.n5388 vss.n194 146.25
R4401 vss.n5386 vss.n190 146.25
R4402 vss.n776 vss.n187 146.25
R4403 vss.n807 vss.n183 146.25
R4404 vss.n5378 vss.n179 146.25
R4405 vss.n5376 vss.n175 146.25
R4406 vss.n808 vss.n167 146.25
R4407 vss.n5957 vss.n168 146.25
R4408 vss.n5368 vss.n163 146.25
R4409 vss.n5366 vss.n158 146.25
R4410 vss.n841 vss.n144 146.25
R4411 vss.n5389 vss.n197 146.25
R4412 vss.n5921 vss.n5920 146.25
R4413 vss.n2641 vss.n2637 146.25
R4414 vss.n2531 vss.n2530 146.25
R4415 vss.n2510 vss.n2507 146.25
R4416 vss.n2344 vss.n1063 146.25
R4417 vss.n4896 vss.n746 137.529
R4418 vss.n2224 vss.n2223 117.001
R4419 vss.n2225 vss.n2224 117.001
R4420 vss.n4224 vss.n4223 117.001
R4421 vss.n4225 vss.n4224 117.001
R4422 vss.n2971 vss.n2970 117.001
R4423 vss.n2970 vss.n1325 117.001
R4424 vss.n2403 vss.n2402 117.001
R4425 vss.n2402 vss.n2401 117.001
R4426 vss.n2236 vss.n2232 117.001
R4427 vss.n2282 vss.n2232 117.001
R4428 vss.n2437 vss.n2436 117.001
R4429 vss.n2436 vss.n2435 117.001
R4430 vss.n5530 vss.n5529 117.001
R4431 vss.n5529 vss.n5528 117.001
R4432 vss.n5397 vss.n733 115.227
R4433 vss.n4898 vss.n4897 111.352
R4434 vss.n5398 vss.n5397 111.352
R4435 vss.n5401 vss.n5400 111.352
R4436 vss.n4588 vss.n4587 111.352
R4437 vss.n4897 vss.n4896 111.352
R4438 vss.n5399 vss.n5398 111.352
R4439 vss.n5402 vss.n5401 111.352
R4440 vss.n2530 vss.n2529 100.588
R4441 vss.n2543 vss.n2542 100.588
R4442 vss.n2663 vss.n2662 100.588
R4443 vss.n774 vss.n773 100.588
R4444 vss.n5389 vss.n5388 100.588
R4445 vss.n2678 vss.n595 97.8689
R4446 vss.n5389 vss.n775 97.8689
R4447 vss.n5920 vss.n215 95.1503
R4448 vss.n2655 vss.t23 93.7911
R4449 vss.n752 vss.n751 92.4318
R4450 vss.n5385 vss.n776 92.4318
R4451 vss.n2521 vss.n399 89.7132
R4452 vss.n2642 vss.n2641 89.7132
R4453 vss.n5387 vss.n5386 89.7132
R4454 vss.n2545 vss.t287 88.3539
R4455 vss.n2643 vss.n567 86.9946
R4456 vss.n2680 vss.n2679 86.9946
R4457 vss.n2763 vss.n2762 86.9946
R4458 vss.n2511 vss.n2510 84.2761
R4459 vss.n2557 vss.n2556 84.2761
R4460 vss.n2761 vss.n214 84.2761
R4461 vss.n5379 vss.n5378 84.2761
R4462 vss.n2512 vss.n385 81.5575
R4463 vss.n2632 vss.n2631 81.5575
R4464 vss.n807 vss.n806 81.5575
R4465 vss.n2572 vss.n455 78.8389
R4466 vss.n2633 vss.n553 78.8389
R4467 vss.n2688 vss.n2687 78.8389
R4468 vss.n2498 vss.n2497 76.1204
R4469 vss.n5375 vss.n808 76.1204
R4470 vss.n2499 vss.n371 73.4018
R4471 vss.n2705 vss.n637 73.4018
R4472 vss.n5377 vss.n5376 73.4018
R4473 vss.n2755 vss.t273 72.0425
R4474 vss.n2581 vss.n469 70.6832
R4475 vss.n2563 vss.t271 69.3239
R4476 vss.n2696 vss.t14 69.3239
R4477 vss.n2461 vss.n1014 67.9647
R4478 vss.n2491 vss.n2490 67.9647
R4479 vss.n2747 vss.n707 67.9647
R4480 vss.n5369 vss.n5368 67.9647
R4481 vss.n5531 vss.n303 66.8263
R4482 vss.t278 vss.n427 66.6054
R4483 vss.t19 vss.n2564 66.6054
R4484 vss.n2622 vss.t275 66.6054
R4485 vss.n2623 vss.t31 66.6054
R4486 vss.n2756 vss.t39 66.6054
R4487 vss.n2299 vss.n2298 66.3945
R4488 vss.n2492 vss.n357 65.2461
R4489 vss.n2715 vss.n651 65.2461
R4490 vss.n814 vss.n168 65.2461
R4491 vss.n2418 vss.n1033 65.0005
R4492 vss.n5182 vss.n1051 65.0005
R4493 vss.n2343 vss.n1045 65.0005
R4494 vss.n5176 vss.n1063 65.0005
R4495 vss.n2329 vss.n1057 65.0005
R4496 vss.n5170 vss.n1075 65.0005
R4497 vss.n4205 vss.n1069 65.0005
R4498 vss.n5164 vss.n1087 65.0005
R4499 vss.n3021 vss.n1081 65.0005
R4500 vss.n5158 vss.n1099 65.0005
R4501 vss.n4226 vss.n1093 65.0005
R4502 vss.n5152 vss.n1111 65.0005
R4503 vss.n1293 vss.n1105 65.0005
R4504 vss.n5146 vss.n4234 65.0005
R4505 vss.n2226 vss.n1115 65.0005
R4506 vss.n5406 vss.n214 65.0005
R4507 vss.n2762 vss.n719 65.0005
R4508 vss.n5410 vss.n721 65.0005
R4509 vss.n2755 vss.n705 65.0005
R4510 vss.n5414 vss.n707 65.0005
R4511 vss.n2746 vss.n691 65.0005
R4512 vss.n5418 vss.n693 65.0005
R4513 vss.n2736 vss.n677 65.0005
R4514 vss.n5422 vss.n679 65.0005
R4515 vss.n2726 vss.n663 65.0005
R4516 vss.n5426 vss.n665 65.0005
R4517 vss.n2716 vss.n649 65.0005
R4518 vss.n5430 vss.n651 65.0005
R4519 vss.n2706 vss.n635 65.0005
R4520 vss.n5434 vss.n637 65.0005
R4521 vss.n2697 vss.n621 65.0005
R4522 vss.n5438 vss.n623 65.0005
R4523 vss.n2687 vss.n607 65.0005
R4524 vss.n5442 vss.n609 65.0005
R4525 vss.n2679 vss.n593 65.0005
R4526 vss.n5446 vss.n595 65.0005
R4527 vss.n2664 vss.n579 65.0005
R4528 vss.n5450 vss.n581 65.0005
R4529 vss.n2654 vss.n565 65.0005
R4530 vss.n5454 vss.n567 65.0005
R4531 vss.n2642 vss.n551 65.0005
R4532 vss.n5458 vss.n553 65.0005
R4533 vss.n2632 vss.n537 65.0005
R4534 vss.n5462 vss.n539 65.0005
R4535 vss.n2622 vss.n523 65.0005
R4536 vss.n5466 vss.n525 65.0005
R4537 vss.n2609 vss.n509 65.0005
R4538 vss.n5470 vss.n511 65.0005
R4539 vss.n2601 vss.n495 65.0005
R4540 vss.n5474 vss.n497 65.0005
R4541 vss.n2592 vss.n481 65.0005
R4542 vss.n5478 vss.n483 65.0005
R4543 vss.n2582 vss.n467 65.0005
R4544 vss.n5482 vss.n469 65.0005
R4545 vss.n453 vss.n223 65.0005
R4546 vss.n5486 vss.n455 65.0005
R4547 vss.n2564 vss.n439 65.0005
R4548 vss.n5490 vss.n441 65.0005
R4549 vss.n2556 vss.n425 65.0005
R4550 vss.n5494 vss.n427 65.0005
R4551 vss.n2544 vss.n411 65.0005
R4552 vss.n5498 vss.n413 65.0005
R4553 vss.n2530 vss.n397 65.0005
R4554 vss.n5502 vss.n399 65.0005
R4555 vss.n2520 vss.n383 65.0005
R4556 vss.n5506 vss.n385 65.0005
R4557 vss.n2511 vss.n369 65.0005
R4558 vss.n5510 vss.n371 65.0005
R4559 vss.n2498 vss.n355 65.0005
R4560 vss.n5514 vss.n357 65.0005
R4561 vss.n2491 vss.n341 65.0005
R4562 vss.n5518 vss.n343 65.0005
R4563 vss.n2482 vss.n327 65.0005
R4564 vss.n5522 vss.n329 65.0005
R4565 vss.n2472 vss.n313 65.0005
R4566 vss.n5527 vss.n5526 65.0005
R4567 vss.n2460 vss.n308 65.0005
R4568 vss.n5208 vss.n1014 65.0005
R4569 vss.n2455 vss.n1009 65.0005
R4570 vss.n5201 vss.n1027 65.0005
R4571 vss.n2385 vss.n1021 65.0005
R4572 vss.n5188 vss.n1039 65.0005
R4573 vss.n2654 vss.t8 63.8868
R4574 vss.n2610 vss.n525 62.5275
R4575 vss.n2736 vss.n2735 62.5275
R4576 vss.t307 vss.n609 61.1682
R4577 vss.t12 vss.n2697 61.1682
R4578 vss.n5527 vss.n307 59.809
R4579 vss.n2482 vss.n2481 59.809
R4580 vss.n2583 vss.n2582 59.809
R4581 vss.n2737 vss.n693 59.809
R4582 vss.n5365 vss.n841 59.809
R4583 vss.n2299 vss.n2203 59.4829
R4584 vss.n2324 vss.n2203 59.4829
R4585 vss.n2325 vss.n2324 59.4829
R4586 vss.n3018 vss.n2325 59.4829
R4587 vss.n3018 vss.n3017 59.4829
R4588 vss.n3017 vss.n3016 59.4829
R4589 vss.n3016 vss.n2327 59.4829
R4590 vss.n2415 vss.n2327 59.4829
R4591 vss.n2415 vss.n2414 59.4829
R4592 vss.n2414 vss.n303 59.4829
R4593 vss.n5394 vss.n752 58.5005
R4594 vss.n2520 vss.t21 58.4497
R4595 vss.n2460 vss.n306 57.0904
R4596 vss.n2483 vss.n343 57.0904
R4597 vss.n2601 vss.n2600 57.0904
R4598 vss.n5367 vss.n5366 57.0904
R4599 vss.n3647 vss.n2193 56.9458
R4600 vss.n3647 vss.n2189 56.9458
R4601 vss.n2189 vss.n2185 56.9458
R4602 vss.n2185 vss.n2181 56.9458
R4603 vss.n2181 vss.n2177 56.9458
R4604 vss.n2177 vss.n2173 56.9458
R4605 vss.n2173 vss.n2169 56.9458
R4606 vss.n2169 vss.n2165 56.9458
R4607 vss.n2165 vss.n2161 56.9458
R4608 vss.n2161 vss.n2157 56.9458
R4609 vss.n2157 vss.n2149 56.9458
R4610 vss.n3680 vss.n2149 56.9458
R4611 vss.n3680 vss.n2145 56.9458
R4612 vss.n2145 vss.n2141 56.9458
R4613 vss.n2141 vss.n2137 56.9458
R4614 vss.n2137 vss.n2133 56.9458
R4615 vss.n2133 vss.n2129 56.9458
R4616 vss.n2129 vss.n2125 56.9458
R4617 vss.n2125 vss.n2121 56.9458
R4618 vss.n2121 vss.n2117 56.9458
R4619 vss.n2117 vss.n2113 56.9458
R4620 vss.n2113 vss.n2109 56.9458
R4621 vss.n2109 vss.n2091 56.9458
R4622 vss.n3716 vss.n2091 56.9458
R4623 vss.n3716 vss.n2087 56.9458
R4624 vss.n2087 vss.n2083 56.9458
R4625 vss.n2083 vss.n2079 56.9458
R4626 vss.n2079 vss.n2075 56.9458
R4627 vss.n2075 vss.n2071 56.9458
R4628 vss.n2071 vss.n2067 56.9458
R4629 vss.n2067 vss.n2063 56.9458
R4630 vss.n2063 vss.n2059 56.9458
R4631 vss.n2059 vss.n2055 56.9458
R4632 vss.n2055 vss.n2037 56.9458
R4633 vss.n3749 vss.n2037 56.9458
R4634 vss.n3749 vss.n2033 56.9458
R4635 vss.n2033 vss.n2029 56.9458
R4636 vss.n2029 vss.n2025 56.9458
R4637 vss.n2025 vss.n2021 56.9458
R4638 vss.n2021 vss.n2017 56.9458
R4639 vss.n2017 vss.n2013 56.9458
R4640 vss.n2013 vss.n2009 56.9458
R4641 vss.n2009 vss.n2005 56.9458
R4642 vss.n2005 vss.n2001 56.9458
R4643 vss.n2001 vss.n1982 56.9458
R4644 vss.n3782 vss.n1982 56.9458
R4645 vss.n3782 vss.n1978 56.9458
R4646 vss.n1978 vss.n1974 56.9458
R4647 vss.n1974 vss.n1970 56.9458
R4648 vss.n1970 vss.n1966 56.9458
R4649 vss.n1966 vss.n1962 56.9458
R4650 vss.n1962 vss.n1958 56.9458
R4651 vss.n1958 vss.n1954 56.9458
R4652 vss.n1954 vss.n1950 56.9458
R4653 vss.n1950 vss.n1946 56.9458
R4654 vss.n1946 vss.n1942 56.9458
R4655 vss.n1942 vss.n1924 56.9458
R4656 vss.n3818 vss.n1924 56.9458
R4657 vss.n3818 vss.n1920 56.9458
R4658 vss.n1920 vss.n1916 56.9458
R4659 vss.n1916 vss.n1912 56.9458
R4660 vss.n1912 vss.n1908 56.9458
R4661 vss.n1908 vss.n1904 56.9458
R4662 vss.n1904 vss.n1900 56.9458
R4663 vss.n1900 vss.n1896 56.9458
R4664 vss.n1896 vss.n1892 56.9458
R4665 vss.n1892 vss.n1888 56.9458
R4666 vss.n1888 vss.n1870 56.9458
R4667 vss.n3851 vss.n1870 56.9458
R4668 vss.n3851 vss.n1866 56.9458
R4669 vss.n1866 vss.n1862 56.9458
R4670 vss.n1862 vss.n1858 56.9458
R4671 vss.n1858 vss.n1854 56.9458
R4672 vss.n1854 vss.n1850 56.9458
R4673 vss.n1850 vss.n1846 56.9458
R4674 vss.n1846 vss.n1842 56.9458
R4675 vss.n1842 vss.n1838 56.9458
R4676 vss.n1838 vss.n1834 56.9458
R4677 vss.n1834 vss.n1815 56.9458
R4678 vss.n3884 vss.n1815 56.9458
R4679 vss.n3884 vss.n1811 56.9458
R4680 vss.n1811 vss.n1807 56.9458
R4681 vss.n1807 vss.n1803 56.9458
R4682 vss.n1803 vss.n1799 56.9458
R4683 vss.n1799 vss.n1795 56.9458
R4684 vss.n1795 vss.n1791 56.9458
R4685 vss.n1791 vss.n1787 56.9458
R4686 vss.n1787 vss.n1783 56.9458
R4687 vss.n1783 vss.n1779 56.9458
R4688 vss.n1779 vss.n1775 56.9458
R4689 vss.n1775 vss.n1767 56.9458
R4690 vss.n3920 vss.n1767 56.9458
R4691 vss.n3920 vss.n1763 56.9458
R4692 vss.n1763 vss.n1759 56.9458
R4693 vss.n1759 vss.n1755 56.9458
R4694 vss.n1755 vss.n1751 56.9458
R4695 vss.n1751 vss.n1747 56.9458
R4696 vss.n1747 vss.n1743 56.9458
R4697 vss.n1743 vss.n1739 56.9458
R4698 vss.n1739 vss.n1735 56.9458
R4699 vss.n1735 vss.n1731 56.9458
R4700 vss.n1731 vss.n1712 56.9458
R4701 vss.n3953 vss.n1712 56.9458
R4702 vss.n3953 vss.n1708 56.9458
R4703 vss.n1708 vss.n1704 56.9458
R4704 vss.n1704 vss.n1700 56.9458
R4705 vss.n1700 vss.n1696 56.9458
R4706 vss.n1696 vss.n1692 56.9458
R4707 vss.n1692 vss.n1688 56.9458
R4708 vss.n1688 vss.n1684 56.9458
R4709 vss.n1684 vss.n1680 56.9458
R4710 vss.n1680 vss.n1676 56.9458
R4711 vss.n1676 vss.n1672 56.9458
R4712 vss.n1672 vss.n1654 56.9458
R4713 vss.n3989 vss.n1654 56.9458
R4714 vss.n3989 vss.n1650 56.9458
R4715 vss.n1650 vss.n1646 56.9458
R4716 vss.n1646 vss.n1642 56.9458
R4717 vss.n1642 vss.n1638 56.9458
R4718 vss.n1638 vss.n1634 56.9458
R4719 vss.n1634 vss.n1630 56.9458
R4720 vss.n1630 vss.n1626 56.9458
R4721 vss.n1626 vss.n1622 56.9458
R4722 vss.n1622 vss.n1618 56.9458
R4723 vss.n1618 vss.n1600 56.9458
R4724 vss.n4022 vss.n1600 56.9458
R4725 vss.n4022 vss.n1596 56.9458
R4726 vss.n1596 vss.n1592 56.9458
R4727 vss.n1592 vss.n1588 56.9458
R4728 vss.n1588 vss.n1584 56.9458
R4729 vss.n1584 vss.n1580 56.9458
R4730 vss.n1580 vss.n1576 56.9458
R4731 vss.n1576 vss.n1572 56.9458
R4732 vss.n1572 vss.n1568 56.9458
R4733 vss.n1568 vss.n1564 56.9458
R4734 vss.n1564 vss.n1545 56.9458
R4735 vss.n4055 vss.n1545 56.9458
R4736 vss.n4055 vss.n1541 56.9458
R4737 vss.n1541 vss.n1537 56.9458
R4738 vss.n1537 vss.n1533 56.9458
R4739 vss.n1533 vss.n1529 56.9458
R4740 vss.n1529 vss.n1525 56.9458
R4741 vss.n1525 vss.n1521 56.9458
R4742 vss.n1521 vss.n1517 56.9458
R4743 vss.n1517 vss.n1513 56.9458
R4744 vss.n1513 vss.n1509 56.9458
R4745 vss.n1509 vss.n1505 56.9458
R4746 vss.n1505 vss.n1487 56.9458
R4747 vss.n4091 vss.n1487 56.9458
R4748 vss.n4091 vss.n1483 56.9458
R4749 vss.n1483 vss.n1479 56.9458
R4750 vss.n1479 vss.n1475 56.9458
R4751 vss.n1475 vss.n1471 56.9458
R4752 vss.n1471 vss.n1467 56.9458
R4753 vss.n1467 vss.n1463 56.9458
R4754 vss.n1463 vss.n1459 56.9458
R4755 vss.n1459 vss.n1455 56.9458
R4756 vss.n1455 vss.n1451 56.9458
R4757 vss.n1451 vss.n1433 56.9458
R4758 vss.n4124 vss.n1433 56.9458
R4759 vss.n4124 vss.n1429 56.9458
R4760 vss.n1429 vss.n1425 56.9458
R4761 vss.n1425 vss.n1421 56.9458
R4762 vss.n1421 vss.n1417 56.9458
R4763 vss.n1417 vss.n1413 56.9458
R4764 vss.n1413 vss.n1409 56.9458
R4765 vss.n1409 vss.n1405 56.9458
R4766 vss.n1405 vss.n1401 56.9458
R4767 vss.n1401 vss.n1397 56.9458
R4768 vss.n1397 vss.n1389 56.9458
R4769 vss.n4157 vss.n1389 56.9458
R4770 vss.n4157 vss.n1385 56.9458
R4771 vss.n1385 vss.n1381 56.9458
R4772 vss.n1381 vss.n1377 56.9458
R4773 vss.n1377 vss.n1373 56.9458
R4774 vss.n1373 vss.n1369 56.9458
R4775 vss.n1369 vss.n1365 56.9458
R4776 vss.n1365 vss.n1361 56.9458
R4777 vss.n1361 vss.n1294 56.9458
R4778 vss.n1354 vss.n1294 56.9458
R4779 vss.n1354 vss.n1350 56.9458
R4780 vss.n1350 vss.n1342 56.9458
R4781 vss.n4193 vss.n1342 56.9458
R4782 vss.n4193 vss.n1337 56.9458
R4783 vss.n1337 vss.n1326 56.9458
R4784 vss.n4203 vss.n1326 56.9458
R4785 vss.n4203 vss.n1329 56.9458
R4786 vss.n2991 vss.n1329 56.9458
R4787 vss.n2991 vss.n2344 56.9458
R4788 vss.n3005 vss.n2344 56.9458
R4789 vss.n3005 vss.n2347 56.9458
R4790 vss.n2353 vss.n2347 56.9458
R4791 vss.n2356 vss.n2353 56.9458
R4792 vss.n2363 vss.n2356 56.9458
R4793 vss.n2364 vss.n2363 56.9458
R4794 vss.n2365 vss.n2364 56.9458
R4795 vss.n2457 vss.n2365 56.9458
R4796 vss.n2462 vss.n2457 56.9458
R4797 vss.n2466 vss.n2462 56.9458
R4798 vss.n2469 vss.n2466 56.9458
R4799 vss.n2474 vss.n2469 56.9458
R4800 vss.n2477 vss.n2474 56.9458
R4801 vss.n2484 vss.n2477 56.9458
R4802 vss.n2487 vss.n2484 56.9458
R4803 vss.n2493 vss.n2487 56.9458
R4804 vss.n2496 vss.n2493 56.9458
R4805 vss.n2500 vss.n2496 56.9458
R4806 vss.n2507 vss.n2500 56.9458
R4807 vss.n2513 vss.n2507 56.9458
R4808 vss.n2516 vss.n2513 56.9458
R4809 vss.n2522 vss.n2516 56.9458
R4810 vss.n2528 vss.n2522 56.9458
R4811 vss.n2531 vss.n2528 56.9458
R4812 vss.n2535 vss.n2531 56.9458
R4813 vss.n2538 vss.n2535 56.9458
R4814 vss.n2546 vss.n2538 56.9458
R4815 vss.n2549 vss.n2546 56.9458
R4816 vss.n2558 vss.n2549 56.9458
R4817 vss.n2559 vss.n2558 56.9458
R4818 vss.n2566 vss.n2559 56.9458
R4819 vss.n2573 vss.n2566 56.9458
R4820 vss.n2574 vss.n2573 56.9458
R4821 vss.n2578 vss.n2574 56.9458
R4822 vss.n2584 vss.n2578 56.9458
R4823 vss.n2588 vss.n2584 56.9458
R4824 vss.n2594 vss.n2588 56.9458
R4825 vss.n2597 vss.n2594 56.9458
R4826 vss.n2603 vss.n2597 56.9458
R4827 vss.n2607 vss.n2603 56.9458
R4828 vss.n2611 vss.n2607 56.9458
R4829 vss.n2618 vss.n2611 56.9458
R4830 vss.n2624 vss.n2618 56.9458
R4831 vss.n2627 vss.n2624 56.9458
R4832 vss.n2634 vss.n2627 56.9458
R4833 vss.n2637 vss.n2634 56.9458
R4834 vss.n2644 vss.n2637 56.9458
R4835 vss.n2647 vss.n2644 56.9458
R4836 vss.n2656 vss.n2647 56.9458
R4837 vss.n2657 vss.n2656 56.9458
R4838 vss.n2661 vss.n2657 56.9458
R4839 vss.n2666 vss.n2661 56.9458
R4840 vss.n2672 vss.n2666 56.9458
R4841 vss.n2681 vss.n2672 56.9458
R4842 vss.n2682 vss.n2681 56.9458
R4843 vss.n2689 vss.n2682 56.9458
R4844 vss.n2692 vss.n2689 56.9458
R4845 vss.n2699 vss.n2692 56.9458
R4846 vss.n2702 vss.n2699 56.9458
R4847 vss.n2708 vss.n2702 56.9458
R4848 vss.n2711 vss.n2708 56.9458
R4849 vss.n2718 vss.n2711 56.9458
R4850 vss.n2724 vss.n2718 56.9458
R4851 vss.n2728 vss.n2724 56.9458
R4852 vss.n2732 vss.n2728 56.9458
R4853 vss.n2738 vss.n2732 56.9458
R4854 vss.n2742 vss.n2738 56.9458
R4855 vss.n2748 vss.n2742 56.9458
R4856 vss.n2751 vss.n2748 56.9458
R4857 vss.n2757 vss.n2751 56.9458
R4858 vss.n2764 vss.n2757 56.9458
R4859 vss.n2764 vss.n211 56.9458
R4860 vss.n5921 vss.n211 56.9458
R4861 vss.n5921 vss.n207 56.9458
R4862 vss.n207 vss.n204 56.9458
R4863 vss.n204 vss.n200 56.9458
R4864 vss.n200 vss.n197 56.9458
R4865 vss.n197 vss.n194 56.9458
R4866 vss.n194 vss.n190 56.9458
R4867 vss.n190 vss.n187 56.9458
R4868 vss.n187 vss.n183 56.9458
R4869 vss.n183 vss.n179 56.9458
R4870 vss.n179 vss.n175 56.9458
R4871 vss.n175 vss.n167 56.9458
R4872 vss.n5957 vss.n167 56.9458
R4873 vss.n5957 vss.n163 56.9458
R4874 vss.n163 vss.n158 56.9458
R4875 vss.n158 vss.n144 56.9458
R4876 vss.n6002 vss.n144 56.9458
R4877 vss.n6009 vss.n135 56.9458
R4878 vss.n896 vss.n869 56.7398
R4879 vss.n1002 vss.n891 56.7398
R4880 vss.n898 vss.n871 56.7398
R4881 vss.n1000 vss.n887 56.7398
R4882 vss.n900 vss.n873 56.7398
R4883 vss.n970 vss.n885 56.7398
R4884 vss.n902 vss.n875 56.7398
R4885 vss.n5358 vss.n878 56.7398
R4886 vss.n5359 vss.n877 56.7398
R4887 vss.n912 vss.n911 56.7398
R4888 vss.n6008 vss.n138 56.7398
R4889 vss.n6007 vss.n6006 56.7398
R4890 vss.n6006 vss.n137 56.7398
R4891 vss.n1002 vss.n896 56.7398
R4892 vss.n891 vss.n871 56.7398
R4893 vss.n1000 vss.n898 56.7398
R4894 vss.n887 vss.n873 56.7398
R4895 vss.n970 vss.n900 56.7398
R4896 vss.n885 vss.n875 56.7398
R4897 vss.n902 vss.n878 56.7398
R4898 vss.n5359 vss.n5358 56.7398
R4899 vss.n912 vss.n877 56.7398
R4900 vss.n3026 vss.n869 56.7398
R4901 vss.n150 vss.n137 56.7398
R4902 vss.n138 vss.n136 56.7398
R4903 vss.n6008 vss.n6007 56.7398
R4904 vss.t4 vss.n2455 55.7311
R4905 vss.n2600 vss.n497 54.3718
R4906 vss.n2602 vss.n511 54.3718
R4907 vss.n2717 vss.n2716 54.3718
R4908 vss.n2726 vss.n2725 54.3718
R4909 vss.n775 vss.n754 53.1823
R4910 vss.n5390 vss.n5389 53.1823
R4911 vss.n5387 vss.n766 53.1823
R4912 vss.n5385 vss.n5384 53.1823
R4913 vss.n806 vss.n782 53.1823
R4914 vss.n5380 vss.n5379 53.1823
R4915 vss.n5377 vss.n799 53.1823
R4916 vss.n5375 vss.n5374 53.1823
R4917 vss.n815 vss.n814 53.1823
R4918 vss.n5370 vss.n5369 53.1823
R4919 vss.n5367 vss.n834 53.1823
R4920 vss.n5365 vss.n5364 53.1823
R4921 vss.n2530 vss.t309 53.0125
R4922 vss.n2472 vss.n307 51.6533
R4923 vss.n2481 vss.n329 51.6533
R4924 vss.n2593 vss.n2592 51.6533
R4925 vss.t285 vss.n224 50.294
R4926 vss.n2707 vss.t10 50.294
R4927 vss.n2473 vss.n2472 48.9347
R4928 vss.n2473 vss.n329 48.9347
R4929 vss.n2592 vss.n2591 48.9347
R4930 vss.n2735 vss.n679 48.9347
R4931 vss.t27 vss.n2608 47.5754
R4932 vss.t299 vss.n2664 47.5754
R4933 vss.n2665 vss.t299 47.5754
R4934 vss.t296 vss.n2745 47.5754
R4935 vss.n2608 vss.n511 46.2161
R4936 vss.n2727 vss.n2726 46.2161
R4937 vss.t309 vss.n413 44.8568
R4938 vss.n2430 vss.n2388 43.4976
R4939 vss.n2461 vss.n2460 43.4976
R4940 vss.n2490 vss.n343 43.4976
R4941 vss.n2717 vss.n665 43.4976
R4942 vss.n5368 vss.n5367 43.4976
R4943 vss.n2430 vss.n1039 40.779
R4944 vss.n2433 vss.n2385 40.779
R4945 vss.n2453 vss.n1027 40.779
R4946 vss.n2483 vss.n2482 40.779
R4947 vss.n2745 vss.n693 40.779
R4948 vss.n5366 vss.n5365 40.779
R4949 vss.n2583 vss.n483 38.0604
R4950 vss.n2621 vss.n525 38.0604
R4951 vss.n2706 vss.n2705 38.0604
R4952 vss.n3605 vss.n3081 37.1593
R4953 vss.n3604 vss.n3081 37.1593
R4954 vss.n3081 vss.n3078 37.1593
R4955 vss.n3607 vss.n3081 37.1593
R4956 vss.n5528 vss.n5527 36.7011
R4957 vss.n2716 vss.t302 36.7011
R4958 vss.n299 vss.n296 36.4064
R4959 vss.n5574 vss.n276 36.4064
R4960 vss.n5806 vss.n5802 36.4064
R4961 vss.n5572 vss.n276 36.4064
R4962 vss.n276 vss.n272 36.4064
R4963 vss.n5539 vss.n299 36.4064
R4964 vss.n2454 vss.n2453 35.3419
R4965 vss.n2455 vss.n2454 35.3419
R4966 vss.n2497 vss.n357 35.3419
R4967 vss.n2610 vss.n2609 35.3419
R4968 vss.n2707 vss.n651 35.3419
R4969 vss.n814 vss.n808 35.3419
R4970 vss.n4369 vss.n4368 34.5783
R4971 vss.n4384 vss.n4383 34.5514
R4972 vss.n4370 vss.n4369 34.5141
R4973 vss.n4373 vss.n4364 34.5141
R4974 vss.n4376 vss.n4362 34.5141
R4975 vss.n4380 vss.n4325 34.5141
R4976 vss.n5803 vss.n5755 34.5082
R4977 vss.n4383 vss.n4322 34.4441
R4978 vss.n4380 vss.n4379 34.4354
R4979 vss.n4376 vss.n4375 34.4354
R4980 vss.n4374 vss.n4373 34.4354
R4981 vss.n4370 vss.n4363 34.4354
R4982 vss.n4368 vss.n4367 34.4354
R4983 vss.n5544 vss.n5543 34.4354
R4984 vss.n5578 vss.n5577 34.4346
R4985 vss.n286 vss.n274 34.4346
R4986 vss.n5575 vss.n269 34.4346
R4987 vss.n5540 vss.n295 34.4324
R4988 vss.n5582 vss.n269 34.4287
R4989 vss.n286 vss.n267 34.4287
R4990 vss.n2298 vss.n2297 34.2957
R4991 vss.t21 vss.n2519 33.9826
R4992 vss.t8 vss.n2653 33.9826
R4993 vss.n2456 vss.n1014 32.6233
R4994 vss.n2492 vss.n2491 32.6233
R4995 vss.n2572 vss.n223 32.6233
R4996 vss.n2754 vss.n707 32.6233
R4997 vss.n5369 vss.n168 32.6233
R4998 vss.n4491 vss.t35 31.838
R4999 vss.n4268 vss.t40 31.838
R5000 vss.n5753 vss.t319 31.6481
R5001 vss.n5659 vss.t32 31.6481
R5002 vss.n2582 vss.t269 31.264
R5003 vss.t33 vss.n483 31.264
R5004 vss.n2591 vss.t33 31.264
R5005 vss.t29 vss.n2601 31.264
R5006 vss.n2725 vss.t17 31.264
R5007 vss.n5147 vss.n1114 30.8711
R5008 vss.n5151 vss.n1092 30.8711
R5009 vss.n5159 vss.n1090 30.8711
R5010 vss.n5163 vss.n1068 30.8711
R5011 vss.n5171 vss.n1066 30.8711
R5012 vss.n5175 vss.n1044 30.8711
R5013 vss.n5183 vss.n1042 30.8711
R5014 vss.n5187 vss.n1020 30.8711
R5015 vss.n5202 vss.n1018 30.8711
R5016 vss.n5207 vss.n318 30.8711
R5017 vss.n5525 vss.n5524 30.8711
R5018 vss.n5523 vss.n322 30.8711
R5019 vss.n5517 vss.n5516 30.8711
R5020 vss.n5515 vss.n350 30.8711
R5021 vss.n5509 vss.n5508 30.8711
R5022 vss.n5507 vss.n378 30.8711
R5023 vss.n5501 vss.n5500 30.8711
R5024 vss.n5499 vss.n406 30.8711
R5025 vss.n5493 vss.n5492 30.8711
R5026 vss.n5491 vss.n434 30.8711
R5027 vss.n5485 vss.n5484 30.8711
R5028 vss.n5483 vss.n462 30.8711
R5029 vss.n5477 vss.n5476 30.8711
R5030 vss.n5475 vss.n490 30.8711
R5031 vss.n5469 vss.n5468 30.8711
R5032 vss.n5467 vss.n518 30.8711
R5033 vss.n5461 vss.n5460 30.8711
R5034 vss.n5459 vss.n546 30.8711
R5035 vss.n5453 vss.n5452 30.8711
R5036 vss.n5451 vss.n574 30.8711
R5037 vss.n5445 vss.n5444 30.8711
R5038 vss.n5443 vss.n602 30.8711
R5039 vss.n5437 vss.n5436 30.8711
R5040 vss.n5435 vss.n630 30.8711
R5041 vss.n5429 vss.n5428 30.8711
R5042 vss.n5427 vss.n658 30.8711
R5043 vss.n5421 vss.n5420 30.8711
R5044 vss.n5419 vss.n686 30.8711
R5045 vss.n5413 vss.n5412 30.8711
R5046 vss.n5411 vss.n714 30.8711
R5047 vss.n5405 vss.n5404 30.8711
R5048 vss.n914 vss.n740 30.8711
R5049 vss.n917 vss.n762 30.8711
R5050 vss.n920 vss.n777 30.8711
R5051 vss.n923 vss.n793 30.8711
R5052 vss.n926 vss.n809 30.8711
R5053 vss.n929 vss.n828 30.8711
R5054 vss.n932 vss.n842 30.8711
R5055 vss.n883 vss.n860 30.8711
R5056 vss.n943 vss.n942 30.8711
R5057 vss.n941 vss.n940 30.8711
R5058 vss.n1260 vss.n1259 30.8711
R5059 vss.n1255 vss.n1106 30.8711
R5060 vss.n1252 vss.n1094 30.8711
R5061 vss.n1249 vss.n1082 30.8711
R5062 vss.n1246 vss.n1070 30.8711
R5063 vss.n1243 vss.n1058 30.8711
R5064 vss.n1240 vss.n1046 30.8711
R5065 vss.n1237 vss.n1034 30.8711
R5066 vss.n1234 vss.n1022 30.8711
R5067 vss.n1231 vss.n1010 30.8711
R5068 vss.n1228 vss.n309 30.8711
R5069 vss.n1225 vss.n323 30.8711
R5070 vss.n1222 vss.n337 30.8711
R5071 vss.n1219 vss.n351 30.8711
R5072 vss.n1216 vss.n365 30.8711
R5073 vss.n1213 vss.n379 30.8711
R5074 vss.n1210 vss.n393 30.8711
R5075 vss.n1207 vss.n407 30.8711
R5076 vss.n1204 vss.n421 30.8711
R5077 vss.n1201 vss.n435 30.8711
R5078 vss.n1198 vss.n449 30.8711
R5079 vss.n1195 vss.n463 30.8711
R5080 vss.n1192 vss.n477 30.8711
R5081 vss.n1189 vss.n491 30.8711
R5082 vss.n1186 vss.n505 30.8711
R5083 vss.n1183 vss.n519 30.8711
R5084 vss.n1180 vss.n533 30.8711
R5085 vss.n1177 vss.n547 30.8711
R5086 vss.n1174 vss.n561 30.8711
R5087 vss.n1171 vss.n575 30.8711
R5088 vss.n1168 vss.n589 30.8711
R5089 vss.n1165 vss.n603 30.8711
R5090 vss.n1162 vss.n617 30.8711
R5091 vss.n1159 vss.n631 30.8711
R5092 vss.n1156 vss.n645 30.8711
R5093 vss.n1153 vss.n659 30.8711
R5094 vss.n1150 vss.n673 30.8711
R5095 vss.n1147 vss.n687 30.8711
R5096 vss.n1144 vss.n701 30.8711
R5097 vss.n1141 vss.n715 30.8711
R5098 vss.n741 vss.n729 30.8711
R5099 vss.n1136 vss.n747 30.8711
R5100 vss.n1133 vss.n771 30.8711
R5101 vss.n1130 vss.n787 30.8711
R5102 vss.n1127 vss.n805 30.8711
R5103 vss.n1124 vss.n820 30.8711
R5104 vss.n1121 vss.n840 30.8711
R5105 vss.n1118 vss.n852 30.8711
R5106 vss.n5356 vss.n876 30.8711
R5107 vss.n5355 vss.n910 30.8711
R5108 vss.n909 vss.n908 30.8711
R5109 vss.n5145 vss.n1104 30.8711
R5110 vss.n5153 vss.n1102 30.8711
R5111 vss.n5157 vss.n1080 30.8711
R5112 vss.n5165 vss.n1078 30.8711
R5113 vss.n5169 vss.n1056 30.8711
R5114 vss.n5177 vss.n1054 30.8711
R5115 vss.n5181 vss.n1032 30.8711
R5116 vss.n5189 vss.n1030 30.8711
R5117 vss.n5200 vss.n5199 30.8711
R5118 vss.n5195 vss.n1017 30.8711
R5119 vss.n332 vss.n317 30.8711
R5120 vss.n5521 vss.n5520 30.8711
R5121 vss.n5519 vss.n336 30.8711
R5122 vss.n5513 vss.n5512 30.8711
R5123 vss.n5511 vss.n364 30.8711
R5124 vss.n5505 vss.n5504 30.8711
R5125 vss.n5503 vss.n392 30.8711
R5126 vss.n5497 vss.n5496 30.8711
R5127 vss.n5495 vss.n420 30.8711
R5128 vss.n5489 vss.n5488 30.8711
R5129 vss.n5487 vss.n448 30.8711
R5130 vss.n5481 vss.n5480 30.8711
R5131 vss.n5479 vss.n476 30.8711
R5132 vss.n5473 vss.n5472 30.8711
R5133 vss.n5471 vss.n504 30.8711
R5134 vss.n5465 vss.n5464 30.8711
R5135 vss.n5463 vss.n532 30.8711
R5136 vss.n5457 vss.n5456 30.8711
R5137 vss.n5455 vss.n560 30.8711
R5138 vss.n5449 vss.n5448 30.8711
R5139 vss.n5447 vss.n588 30.8711
R5140 vss.n5441 vss.n5440 30.8711
R5141 vss.n5439 vss.n616 30.8711
R5142 vss.n5433 vss.n5432 30.8711
R5143 vss.n5431 vss.n644 30.8711
R5144 vss.n5425 vss.n5424 30.8711
R5145 vss.n5423 vss.n672 30.8711
R5146 vss.n5417 vss.n5416 30.8711
R5147 vss.n5415 vss.n700 30.8711
R5148 vss.n5409 vss.n5408 30.8711
R5149 vss.n5407 vss.n728 30.8711
R5150 vss.n5393 vss.n5392 30.8711
R5151 vss.n5391 vss.n761 30.8711
R5152 vss.n946 vss.n778 30.8711
R5153 vss.n949 vss.n794 30.8711
R5154 vss.n952 vss.n810 30.8711
R5155 vss.n955 vss.n829 30.8711
R5156 vss.n958 vss.n843 30.8711
R5157 vss.n884 vss.n861 30.8711
R5158 vss.n969 vss.n968 30.8711
R5159 vss.n967 vss.n966 30.8711
R5160 vss.n1287 vss.n1286 30.8711
R5161 vss.n1282 vss.n1107 30.8711
R5162 vss.n1279 vss.n1095 30.8711
R5163 vss.n1276 vss.n1083 30.8711
R5164 vss.n1273 vss.n1071 30.8711
R5165 vss.n1270 vss.n1059 30.8711
R5166 vss.n1267 vss.n1047 30.8711
R5167 vss.n1264 vss.n1035 30.8711
R5168 vss.n1023 vss.n1008 30.8711
R5169 vss.n5210 vss.n5209 30.8711
R5170 vss.n5213 vss.n310 30.8711
R5171 vss.n5216 vss.n324 30.8711
R5172 vss.n5219 vss.n338 30.8711
R5173 vss.n5222 vss.n352 30.8711
R5174 vss.n5225 vss.n366 30.8711
R5175 vss.n5228 vss.n380 30.8711
R5176 vss.n5231 vss.n394 30.8711
R5177 vss.n5234 vss.n408 30.8711
R5178 vss.n5237 vss.n422 30.8711
R5179 vss.n5240 vss.n436 30.8711
R5180 vss.n5243 vss.n450 30.8711
R5181 vss.n5246 vss.n464 30.8711
R5182 vss.n5249 vss.n478 30.8711
R5183 vss.n5252 vss.n492 30.8711
R5184 vss.n5255 vss.n506 30.8711
R5185 vss.n5258 vss.n520 30.8711
R5186 vss.n5261 vss.n534 30.8711
R5187 vss.n5264 vss.n548 30.8711
R5188 vss.n5267 vss.n562 30.8711
R5189 vss.n5270 vss.n576 30.8711
R5190 vss.n5273 vss.n590 30.8711
R5191 vss.n5276 vss.n604 30.8711
R5192 vss.n5279 vss.n618 30.8711
R5193 vss.n5282 vss.n632 30.8711
R5194 vss.n5285 vss.n646 30.8711
R5195 vss.n5288 vss.n660 30.8711
R5196 vss.n5291 vss.n674 30.8711
R5197 vss.n5294 vss.n688 30.8711
R5198 vss.n5297 vss.n702 30.8711
R5199 vss.n5300 vss.n716 30.8711
R5200 vss.n742 vss.n730 30.8711
R5201 vss.n5305 vss.n748 30.8711
R5202 vss.n5308 vss.n770 30.8711
R5203 vss.n5311 vss.n786 30.8711
R5204 vss.n5314 vss.n804 30.8711
R5205 vss.n5317 vss.n819 30.8711
R5206 vss.n5320 vss.n839 30.8711
R5207 vss.n5323 vss.n851 30.8711
R5208 vss.n901 vss.n874 30.8711
R5209 vss.n5334 vss.n5333 30.8711
R5210 vss.n5332 vss.n5331 30.8711
R5211 vss.n5143 vss.n5142 30.8711
R5212 vss.n5138 vss.n1113 30.8711
R5213 vss.n5135 vss.n1101 30.8711
R5214 vss.n5132 vss.n1089 30.8711
R5215 vss.n5129 vss.n1077 30.8711
R5216 vss.n5126 vss.n1065 30.8711
R5217 vss.n5123 vss.n1053 30.8711
R5218 vss.n5120 vss.n1041 30.8711
R5219 vss.n5117 vss.n1029 30.8711
R5220 vss.n5114 vss.n1016 30.8711
R5221 vss.n5111 vss.n316 30.8711
R5222 vss.n5108 vss.n331 30.8711
R5223 vss.n5105 vss.n345 30.8711
R5224 vss.n5102 vss.n359 30.8711
R5225 vss.n5099 vss.n373 30.8711
R5226 vss.n5096 vss.n387 30.8711
R5227 vss.n5093 vss.n401 30.8711
R5228 vss.n5090 vss.n415 30.8711
R5229 vss.n5087 vss.n429 30.8711
R5230 vss.n5084 vss.n443 30.8711
R5231 vss.n5081 vss.n457 30.8711
R5232 vss.n5078 vss.n471 30.8711
R5233 vss.n5075 vss.n485 30.8711
R5234 vss.n5072 vss.n499 30.8711
R5235 vss.n5069 vss.n513 30.8711
R5236 vss.n5066 vss.n527 30.8711
R5237 vss.n5063 vss.n541 30.8711
R5238 vss.n5060 vss.n555 30.8711
R5239 vss.n5057 vss.n569 30.8711
R5240 vss.n5054 vss.n583 30.8711
R5241 vss.n5051 vss.n597 30.8711
R5242 vss.n5048 vss.n611 30.8711
R5243 vss.n5045 vss.n625 30.8711
R5244 vss.n5042 vss.n639 30.8711
R5245 vss.n5039 vss.n653 30.8711
R5246 vss.n5036 vss.n667 30.8711
R5247 vss.n5033 vss.n681 30.8711
R5248 vss.n5030 vss.n695 30.8711
R5249 vss.n5027 vss.n709 30.8711
R5250 vss.n5024 vss.n723 30.8711
R5251 vss.n5396 vss.n736 30.8711
R5252 vss.n5395 vss.n745 30.8711
R5253 vss.n973 vss.n763 30.8711
R5254 vss.n976 vss.n779 30.8711
R5255 vss.n979 vss.n795 30.8711
R5256 vss.n982 vss.n811 30.8711
R5257 vss.n985 vss.n830 30.8711
R5258 vss.n988 vss.n844 30.8711
R5259 vss.n886 vss.n862 30.8711
R5260 vss.n999 vss.n998 30.8711
R5261 vss.n997 vss.n996 30.8711
R5262 vss.n4744 vss.n1288 30.8711
R5263 vss.n4747 vss.n1108 30.8711
R5264 vss.n4750 vss.n1096 30.8711
R5265 vss.n4753 vss.n1084 30.8711
R5266 vss.n4756 vss.n1072 30.8711
R5267 vss.n4759 vss.n1060 30.8711
R5268 vss.n4762 vss.n1048 30.8711
R5269 vss.n4765 vss.n1036 30.8711
R5270 vss.n4768 vss.n1024 30.8711
R5271 vss.n4771 vss.n1011 30.8711
R5272 vss.n4774 vss.n311 30.8711
R5273 vss.n4777 vss.n325 30.8711
R5274 vss.n4780 vss.n339 30.8711
R5275 vss.n4783 vss.n353 30.8711
R5276 vss.n4786 vss.n367 30.8711
R5277 vss.n4789 vss.n381 30.8711
R5278 vss.n4792 vss.n395 30.8711
R5279 vss.n4795 vss.n409 30.8711
R5280 vss.n4798 vss.n423 30.8711
R5281 vss.n4801 vss.n437 30.8711
R5282 vss.n4804 vss.n451 30.8711
R5283 vss.n4807 vss.n465 30.8711
R5284 vss.n4810 vss.n479 30.8711
R5285 vss.n4813 vss.n493 30.8711
R5286 vss.n4816 vss.n507 30.8711
R5287 vss.n4819 vss.n521 30.8711
R5288 vss.n4822 vss.n535 30.8711
R5289 vss.n4825 vss.n549 30.8711
R5290 vss.n4828 vss.n563 30.8711
R5291 vss.n4831 vss.n577 30.8711
R5292 vss.n4834 vss.n591 30.8711
R5293 vss.n4837 vss.n605 30.8711
R5294 vss.n4840 vss.n619 30.8711
R5295 vss.n4843 vss.n633 30.8711
R5296 vss.n4846 vss.n647 30.8711
R5297 vss.n4849 vss.n661 30.8711
R5298 vss.n4852 vss.n675 30.8711
R5299 vss.n4855 vss.n689 30.8711
R5300 vss.n4858 vss.n703 30.8711
R5301 vss.n4861 vss.n717 30.8711
R5302 vss.n4895 vss.n731 30.8711
R5303 vss.n4891 vss.n749 30.8711
R5304 vss.n4888 vss.n769 30.8711
R5305 vss.n4885 vss.n785 30.8711
R5306 vss.n4882 vss.n803 30.8711
R5307 vss.n4879 vss.n818 30.8711
R5308 vss.n4876 vss.n838 30.8711
R5309 vss.n4873 vss.n850 30.8711
R5310 vss.n899 vss.n872 30.8711
R5311 vss.n4868 vss.n1006 30.8711
R5312 vss.n4867 vss.n4866 30.8711
R5313 vss.n5021 vss.n5020 30.8711
R5314 vss.n5016 vss.n1112 30.8711
R5315 vss.n5013 vss.n1100 30.8711
R5316 vss.n5010 vss.n1088 30.8711
R5317 vss.n5007 vss.n1076 30.8711
R5318 vss.n5004 vss.n1064 30.8711
R5319 vss.n5001 vss.n1052 30.8711
R5320 vss.n4998 vss.n1040 30.8711
R5321 vss.n4995 vss.n1028 30.8711
R5322 vss.n4992 vss.n1015 30.8711
R5323 vss.n4989 vss.n315 30.8711
R5324 vss.n4986 vss.n330 30.8711
R5325 vss.n4983 vss.n344 30.8711
R5326 vss.n4980 vss.n358 30.8711
R5327 vss.n4977 vss.n372 30.8711
R5328 vss.n4974 vss.n386 30.8711
R5329 vss.n4971 vss.n400 30.8711
R5330 vss.n4968 vss.n414 30.8711
R5331 vss.n4965 vss.n428 30.8711
R5332 vss.n4962 vss.n442 30.8711
R5333 vss.n4959 vss.n456 30.8711
R5334 vss.n4956 vss.n470 30.8711
R5335 vss.n4953 vss.n484 30.8711
R5336 vss.n4950 vss.n498 30.8711
R5337 vss.n4947 vss.n512 30.8711
R5338 vss.n4944 vss.n526 30.8711
R5339 vss.n4941 vss.n540 30.8711
R5340 vss.n4938 vss.n554 30.8711
R5341 vss.n4935 vss.n568 30.8711
R5342 vss.n4932 vss.n582 30.8711
R5343 vss.n4929 vss.n596 30.8711
R5344 vss.n4926 vss.n610 30.8711
R5345 vss.n4923 vss.n624 30.8711
R5346 vss.n4920 vss.n638 30.8711
R5347 vss.n4917 vss.n652 30.8711
R5348 vss.n4914 vss.n666 30.8711
R5349 vss.n4911 vss.n680 30.8711
R5350 vss.n4908 vss.n694 30.8711
R5351 vss.n4905 vss.n708 30.8711
R5352 vss.n4902 vss.n722 30.8711
R5353 vss.n4899 vss.n735 30.8711
R5354 vss.n4263 vss.n756 30.8711
R5355 vss.n4260 vss.n764 30.8711
R5356 vss.n4257 vss.n780 30.8711
R5357 vss.n4254 vss.n796 30.8711
R5358 vss.n4251 vss.n812 30.8711
R5359 vss.n4248 vss.n831 30.8711
R5360 vss.n4245 vss.n845 30.8711
R5361 vss.n888 vss.n863 30.8711
R5362 vss.n4240 vss.n1001 30.8711
R5363 vss.n4239 vss.n4238 30.8711
R5364 vss.n4590 vss.n1289 30.8711
R5365 vss.n4593 vss.n1109 30.8711
R5366 vss.n4596 vss.n1097 30.8711
R5367 vss.n4599 vss.n1085 30.8711
R5368 vss.n4602 vss.n1073 30.8711
R5369 vss.n4605 vss.n1061 30.8711
R5370 vss.n4608 vss.n1049 30.8711
R5371 vss.n4611 vss.n1037 30.8711
R5372 vss.n4614 vss.n1025 30.8711
R5373 vss.n4617 vss.n1012 30.8711
R5374 vss.n4620 vss.n312 30.8711
R5375 vss.n4623 vss.n326 30.8711
R5376 vss.n4626 vss.n340 30.8711
R5377 vss.n4629 vss.n354 30.8711
R5378 vss.n4632 vss.n368 30.8711
R5379 vss.n4635 vss.n382 30.8711
R5380 vss.n4638 vss.n396 30.8711
R5381 vss.n4641 vss.n410 30.8711
R5382 vss.n4644 vss.n424 30.8711
R5383 vss.n4647 vss.n438 30.8711
R5384 vss.n4650 vss.n452 30.8711
R5385 vss.n4653 vss.n466 30.8711
R5386 vss.n4656 vss.n480 30.8711
R5387 vss.n4659 vss.n494 30.8711
R5388 vss.n4662 vss.n508 30.8711
R5389 vss.n4665 vss.n522 30.8711
R5390 vss.n4668 vss.n536 30.8711
R5391 vss.n4671 vss.n550 30.8711
R5392 vss.n4674 vss.n564 30.8711
R5393 vss.n4677 vss.n578 30.8711
R5394 vss.n4680 vss.n592 30.8711
R5395 vss.n4683 vss.n606 30.8711
R5396 vss.n4686 vss.n620 30.8711
R5397 vss.n4689 vss.n634 30.8711
R5398 vss.n4692 vss.n648 30.8711
R5399 vss.n4695 vss.n662 30.8711
R5400 vss.n4698 vss.n676 30.8711
R5401 vss.n4701 vss.n690 30.8711
R5402 vss.n4704 vss.n704 30.8711
R5403 vss.n4707 vss.n718 30.8711
R5404 vss.n4741 vss.n732 30.8711
R5405 vss.n4737 vss.n750 30.8711
R5406 vss.n4734 vss.n768 30.8711
R5407 vss.n4731 vss.n784 30.8711
R5408 vss.n4728 vss.n802 30.8711
R5409 vss.n4725 vss.n817 30.8711
R5410 vss.n4722 vss.n837 30.8711
R5411 vss.n4719 vss.n849 30.8711
R5412 vss.n897 vss.n870 30.8711
R5413 vss.n4714 vss.n1005 30.8711
R5414 vss.n4713 vss.n4712 30.8711
R5415 vss.n788 vss.n772 30.8711
R5416 vss.n5383 vss.n5382 30.8711
R5417 vss.n5381 vss.n792 30.8711
R5418 vss.n5373 vss.n5372 30.8711
R5419 vss.n5371 vss.n827 30.8711
R5420 vss.n5363 vss.n5362 30.8711
R5421 vss.n5361 vss.n859 30.8711
R5422 vss.n5353 vss.n5352 30.8711
R5423 vss.n5351 vss.n5350 30.8711
R5424 vss.n4581 vss.n753 30.8711
R5425 vss.n4577 vss.n767 30.8711
R5426 vss.n800 vss.n783 30.8711
R5427 vss.n821 vss.n801 30.8711
R5428 vss.n835 vss.n816 30.8711
R5429 vss.n853 vss.n836 30.8711
R5430 vss.n867 vss.n848 30.8711
R5431 vss.n894 vss.n868 30.8711
R5432 vss.n5340 vss.n1004 30.8711
R5433 vss.n5342 vss.n5341 30.8711
R5434 vss.n2293 vss.n2292 30.8711
R5435 vss.n2288 vss.n2229 30.8711
R5436 vss.n2307 vss.n1297 30.8711
R5437 vss.n4231 vss.n4230 30.8711
R5438 vss.n4229 vss.n1301 30.8711
R5439 vss.n3022 vss.n1319 30.8711
R5440 vss.n4208 vss.n1320 30.8711
R5441 vss.n2987 vss.n2338 30.8711
R5442 vss.n3009 vss.n2339 30.8711
R5443 vss.n2427 vss.n2390 30.8711
R5444 vss.n2428 vss.n2374 30.8711
R5445 vss.n2242 vss.n2241 30.8711
R5446 vss.n2312 vss.n2209 30.8711
R5447 vss.n2214 vss.n2213 30.8711
R5448 vss.n2210 vss.n1311 30.8711
R5449 vss.n2198 vss.n2197 30.8711
R5450 vss.n2981 vss.n1317 30.8711
R5451 vss.n2984 vss.n2983 30.8711
R5452 vss.n2392 vss.n2336 30.8711
R5453 vss.n2424 vss.n2423 30.8711
R5454 vss.n2387 vss.n2381 30.8711
R5455 vss.n2219 vss.n2207 30.8711
R5456 vss.n1313 vss.n1309 30.8711
R5457 vss.n2975 vss.n2974 30.8711
R5458 vss.n2405 vss.n2396 30.8711
R5459 vss.n2445 vss.n2378 30.8711
R5460 vss.n5535 vss.n5534 30.8711
R5461 vss.n4330 vss.n1290 30.8711
R5462 vss.n4333 vss.n1110 30.8711
R5463 vss.n4336 vss.n1098 30.8711
R5464 vss.n4339 vss.n1086 30.8711
R5465 vss.n4342 vss.n1074 30.8711
R5466 vss.n4345 vss.n1062 30.8711
R5467 vss.n4348 vss.n1050 30.8711
R5468 vss.n4327 vss.n1038 30.8711
R5469 vss.n4356 vss.n1026 30.8711
R5470 vss.n4387 vss.n1013 30.8711
R5471 vss.n4319 vss.n314 30.8711
R5472 vss.n4316 vss.n328 30.8711
R5473 vss.n4403 vss.n342 30.8711
R5474 vss.n4410 vss.n356 30.8711
R5475 vss.n4416 vss.n370 30.8711
R5476 vss.n4308 vss.n384 30.8711
R5477 vss.n4304 vss.n398 30.8711
R5478 vss.n4433 vss.n412 30.8711
R5479 vss.n4441 vss.n426 30.8711
R5480 vss.n4299 vss.n440 30.8711
R5481 vss.n4453 vss.n454 30.8711
R5482 vss.n4461 vss.n468 30.8711
R5483 vss.n4294 vss.n482 30.8711
R5484 vss.n4473 vss.n496 30.8711
R5485 vss.n4481 vss.n510 30.8711
R5486 vss.n4486 vss.n524 30.8711
R5487 vss.n4493 vss.n538 30.8711
R5488 vss.n4497 vss.n552 30.8711
R5489 vss.n4503 vss.n566 30.8711
R5490 vss.n4284 vss.n580 30.8711
R5491 vss.n4515 vss.n594 30.8711
R5492 vss.n4523 vss.n608 30.8711
R5493 vss.n4279 vss.n622 30.8711
R5494 vss.n4535 vss.n636 30.8711
R5495 vss.n4543 vss.n650 30.8711
R5496 vss.n4274 vss.n664 30.8711
R5497 vss.n4555 vss.n678 30.8711
R5498 vss.n4563 vss.n692 30.8711
R5499 vss.n4269 vss.n706 30.8711
R5500 vss.n4571 vss.n720 30.8711
R5501 vss.n4266 vss.n734 30.8711
R5502 vss.n4582 vss.n755 30.8711
R5503 vss.n4578 vss.n765 30.8711
R5504 vss.n797 vss.n781 30.8711
R5505 vss.n822 vss.n798 30.8711
R5506 vss.n832 vss.n813 30.8711
R5507 vss.n854 vss.n833 30.8711
R5508 vss.n864 vss.n846 30.8711
R5509 vss.n892 vss.n865 30.8711
R5510 vss.n5344 vss.n1003 30.8711
R5511 vss.n5346 vss.n5345 30.8711
R5512 vss.n469 vss.n224 29.9047
R5513 vss.n2631 vss.n539 29.9047
R5514 vss.n2697 vss.n2696 29.9047
R5515 vss.n2747 vss.n2746 29.9047
R5516 vss.n3040 vss.n3029 29.4426
R5517 vss.n3040 vss.n3039 29.4426
R5518 vss.n3039 vss.n3038 29.4426
R5519 vss.n3038 vss.n3037 29.4426
R5520 vss.n3037 vss.n3036 29.4426
R5521 vss.n3036 vss.n3035 29.4426
R5522 vss.n3035 vss.n3034 29.4426
R5523 vss.n3034 vss.n3033 29.4426
R5524 vss.n3033 vss.n3032 29.4426
R5525 vss.n3032 vss.n3031 29.4426
R5526 vss.n3031 vss.n3030 29.4426
R5527 vss.n3030 vss.n2150 29.4426
R5528 vss.n2263 vss.n2150 29.4426
R5529 vss.n2264 vss.n2263 29.4426
R5530 vss.n2265 vss.n2264 29.4426
R5531 vss.n2266 vss.n2265 29.4426
R5532 vss.n2267 vss.n2266 29.4426
R5533 vss.n2268 vss.n2267 29.4426
R5534 vss.n2273 vss.n2272 29.4426
R5535 vss.n2272 vss.n2271 29.4426
R5536 vss.n2270 vss.n2269 29.4426
R5537 vss.n2102 vss.n2101 29.4426
R5538 vss.n2100 vss.n2099 29.4426
R5539 vss.n2098 vss.n2097 29.4426
R5540 vss.n2096 vss.n2095 29.4426
R5541 vss.n2094 vss.n2093 29.4426
R5542 vss.n2092 vss.n2048 29.4426
R5543 vss.n2047 vss.n2046 29.4426
R5544 vss.n2045 vss.n2044 29.4426
R5545 vss.n2043 vss.n2042 29.4426
R5546 vss.n2041 vss.n2040 29.4426
R5547 vss.n2039 vss.n2038 29.4426
R5548 vss.n1994 vss.n1993 29.4426
R5549 vss.n1992 vss.n1991 29.4426
R5550 vss.n1990 vss.n1989 29.4426
R5551 vss.n1988 vss.n1987 29.4426
R5552 vss.n1986 vss.n1985 29.4426
R5553 vss.n1984 vss.n1983 29.4426
R5554 vss.n1935 vss.n1934 29.4426
R5555 vss.n1933 vss.n1932 29.4426
R5556 vss.n1931 vss.n1930 29.4426
R5557 vss.n1929 vss.n1928 29.4426
R5558 vss.n1927 vss.n1926 29.4426
R5559 vss.n1925 vss.n1881 29.4426
R5560 vss.n1880 vss.n1879 29.4426
R5561 vss.n1878 vss.n1877 29.4426
R5562 vss.n1876 vss.n1875 29.4426
R5563 vss.n1874 vss.n1873 29.4426
R5564 vss.n1872 vss.n1871 29.4426
R5565 vss.n1827 vss.n1826 29.4426
R5566 vss.n1825 vss.n1824 29.4426
R5567 vss.n1823 vss.n1822 29.4426
R5568 vss.n1821 vss.n1820 29.4426
R5569 vss.n1819 vss.n1818 29.4426
R5570 vss.n1817 vss.n1816 29.4426
R5571 vss.n2251 vss.n1768 29.4426
R5572 vss.n2253 vss.n2252 29.4426
R5573 vss.n2260 vss.n2259 29.4426
R5574 vss.n2258 vss.n2257 29.4426
R5575 vss.n2256 vss.n2255 29.4426
R5576 vss.n2254 vss.n1724 29.4426
R5577 vss.n1723 vss.n1722 29.4426
R5578 vss.n1721 vss.n1720 29.4426
R5579 vss.n1719 vss.n1718 29.4426
R5580 vss.n1717 vss.n1716 29.4426
R5581 vss.n1715 vss.n1714 29.4426
R5582 vss.n1713 vss.n1665 29.4426
R5583 vss.n1664 vss.n1663 29.4426
R5584 vss.n1662 vss.n1661 29.4426
R5585 vss.n1660 vss.n1659 29.4426
R5586 vss.n1658 vss.n1657 29.4426
R5587 vss.n1656 vss.n1655 29.4426
R5588 vss.n1611 vss.n1610 29.4426
R5589 vss.n1609 vss.n1608 29.4426
R5590 vss.n1607 vss.n1606 29.4426
R5591 vss.n1605 vss.n1604 29.4426
R5592 vss.n1603 vss.n1602 29.4426
R5593 vss.n1601 vss.n1557 29.4426
R5594 vss.n1556 vss.n1555 29.4426
R5595 vss.n1554 vss.n1553 29.4426
R5596 vss.n1552 vss.n1551 29.4426
R5597 vss.n1550 vss.n1549 29.4426
R5598 vss.n1548 vss.n1547 29.4426
R5599 vss.n1546 vss.n1498 29.4426
R5600 vss.n1497 vss.n1496 29.4426
R5601 vss.n1495 vss.n1494 29.4426
R5602 vss.n1493 vss.n1492 29.4426
R5603 vss.n1491 vss.n1490 29.4426
R5604 vss.n1489 vss.n1488 29.4426
R5605 vss.n1444 vss.n1443 29.4426
R5606 vss.n1442 vss.n1441 29.4426
R5607 vss.n1440 vss.n1439 29.4426
R5608 vss.n1438 vss.n1437 29.4426
R5609 vss.n1436 vss.n1435 29.4426
R5610 vss.n1434 vss.n1390 29.4426
R5611 vss.n2249 vss.n1390 29.4426
R5612 vss.n2281 vss.n2280 28.6469
R5613 vss.n2555 vss.t278 28.5454
R5614 vss.n2593 vss.t291 28.5454
R5615 vss.n2686 vss.t307 28.5454
R5616 vss.n2727 vss.t25 28.5454
R5617 vss.n3605 vss.n3073 27.8593
R5618 vss.n3614 vss.n3073 27.8593
R5619 vss.n3615 vss.n3614 27.8593
R5620 vss.n3616 vss.n3615 27.8593
R5621 vss.n3616 vss.n3064 27.8593
R5622 vss.n3624 vss.n3064 27.8593
R5623 vss.n3625 vss.n3624 27.8593
R5624 vss.n3625 vss.n3055 27.8593
R5625 vss.n3633 vss.n3055 27.8593
R5626 vss.n3634 vss.n3633 27.8593
R5627 vss.n3634 vss.n3046 27.8593
R5628 vss.n3642 vss.n3046 27.8593
R5629 vss.n3643 vss.n3642 27.8593
R5630 vss.n3643 vss.n3041 27.8593
R5631 vss.n3041 vss.n2184 27.8593
R5632 vss.n3654 vss.n2184 27.8593
R5633 vss.n3655 vss.n3654 27.8593
R5634 vss.n3655 vss.n2172 27.8593
R5635 vss.n3663 vss.n2172 27.8593
R5636 vss.n3664 vss.n3663 27.8593
R5637 vss.n3664 vss.n2160 27.8593
R5638 vss.n3672 vss.n2160 27.8593
R5639 vss.n3673 vss.n3672 27.8593
R5640 vss.n3673 vss.n2148 27.8593
R5641 vss.n3681 vss.n2148 27.8593
R5642 vss.n3682 vss.n3681 27.8593
R5643 vss.n3682 vss.n2136 27.8593
R5644 vss.n3690 vss.n2136 27.8593
R5645 vss.n3691 vss.n3690 27.8593
R5646 vss.n3691 vss.n2124 27.8593
R5647 vss.n3699 vss.n2124 27.8593
R5648 vss.n3700 vss.n3699 27.8593
R5649 vss.n3700 vss.n2112 27.8593
R5650 vss.n3708 vss.n2112 27.8593
R5651 vss.n3709 vss.n3708 27.8593
R5652 vss.n3709 vss.n2090 27.8593
R5653 vss.n3717 vss.n2090 27.8593
R5654 vss.n3718 vss.n3717 27.8593
R5655 vss.n3718 vss.n2078 27.8593
R5656 vss.n3726 vss.n2078 27.8593
R5657 vss.n3727 vss.n3726 27.8593
R5658 vss.n3727 vss.n2066 27.8593
R5659 vss.n3735 vss.n2066 27.8593
R5660 vss.n3736 vss.n3735 27.8593
R5661 vss.n3736 vss.n2054 27.8593
R5662 vss.n3744 vss.n2054 27.8593
R5663 vss.n3745 vss.n3744 27.8593
R5664 vss.n3745 vss.n2049 27.8593
R5665 vss.n2049 vss.n2028 27.8593
R5666 vss.n3756 vss.n2028 27.8593
R5667 vss.n3757 vss.n3756 27.8593
R5668 vss.n3757 vss.n2016 27.8593
R5669 vss.n3765 vss.n2016 27.8593
R5670 vss.n3766 vss.n3765 27.8593
R5671 vss.n3766 vss.n2004 27.8593
R5672 vss.n3774 vss.n2004 27.8593
R5673 vss.n3775 vss.n3774 27.8593
R5674 vss.n3775 vss.n1981 27.8593
R5675 vss.n3783 vss.n1981 27.8593
R5676 vss.n3784 vss.n3783 27.8593
R5677 vss.n3784 vss.n1969 27.8593
R5678 vss.n3792 vss.n1969 27.8593
R5679 vss.n3793 vss.n3792 27.8593
R5680 vss.n3793 vss.n1957 27.8593
R5681 vss.n3801 vss.n1957 27.8593
R5682 vss.n3802 vss.n3801 27.8593
R5683 vss.n3802 vss.n1945 27.8593
R5684 vss.n3810 vss.n1945 27.8593
R5685 vss.n3811 vss.n3810 27.8593
R5686 vss.n3811 vss.n1923 27.8593
R5687 vss.n3819 vss.n1923 27.8593
R5688 vss.n3820 vss.n3819 27.8593
R5689 vss.n3820 vss.n1911 27.8593
R5690 vss.n3828 vss.n1911 27.8593
R5691 vss.n3829 vss.n3828 27.8593
R5692 vss.n3829 vss.n1899 27.8593
R5693 vss.n3837 vss.n1899 27.8593
R5694 vss.n3838 vss.n3837 27.8593
R5695 vss.n3838 vss.n1887 27.8593
R5696 vss.n3846 vss.n1887 27.8593
R5697 vss.n3847 vss.n3846 27.8593
R5698 vss.n3847 vss.n1882 27.8593
R5699 vss.n1882 vss.n1861 27.8593
R5700 vss.n3858 vss.n1861 27.8593
R5701 vss.n3859 vss.n3858 27.8593
R5702 vss.n3859 vss.n1849 27.8593
R5703 vss.n3867 vss.n1849 27.8593
R5704 vss.n3868 vss.n3867 27.8593
R5705 vss.n3868 vss.n1837 27.8593
R5706 vss.n3876 vss.n1837 27.8593
R5707 vss.n3877 vss.n3876 27.8593
R5708 vss.n3877 vss.n1814 27.8593
R5709 vss.n3885 vss.n1814 27.8593
R5710 vss.n3886 vss.n3885 27.8593
R5711 vss.n3886 vss.n1802 27.8593
R5712 vss.n3894 vss.n1802 27.8593
R5713 vss.n3895 vss.n3894 27.8593
R5714 vss.n3895 vss.n1790 27.8593
R5715 vss.n3903 vss.n1790 27.8593
R5716 vss.n3904 vss.n3903 27.8593
R5717 vss.n3904 vss.n1778 27.8593
R5718 vss.n3912 vss.n1778 27.8593
R5719 vss.n3913 vss.n3912 27.8593
R5720 vss.n3913 vss.n1766 27.8593
R5721 vss.n3921 vss.n1766 27.8593
R5722 vss.n3922 vss.n3921 27.8593
R5723 vss.n3922 vss.n1754 27.8593
R5724 vss.n3930 vss.n1754 27.8593
R5725 vss.n3931 vss.n3930 27.8593
R5726 vss.n3931 vss.n1742 27.8593
R5727 vss.n3939 vss.n1742 27.8593
R5728 vss.n3940 vss.n3939 27.8593
R5729 vss.n3940 vss.n1730 27.8593
R5730 vss.n3948 vss.n1730 27.8593
R5731 vss.n3949 vss.n3948 27.8593
R5732 vss.n3949 vss.n1707 27.8593
R5733 vss.n3957 vss.n1707 27.8593
R5734 vss.n3958 vss.n3957 27.8593
R5735 vss.n3958 vss.n1695 27.8593
R5736 vss.n3966 vss.n1695 27.8593
R5737 vss.n3967 vss.n3966 27.8593
R5738 vss.n3967 vss.n1683 27.8593
R5739 vss.n3975 vss.n1683 27.8593
R5740 vss.n3976 vss.n3975 27.8593
R5741 vss.n3976 vss.n1671 27.8593
R5742 vss.n3984 vss.n1671 27.8593
R5743 vss.n3985 vss.n3984 27.8593
R5744 vss.n3985 vss.n1666 27.8593
R5745 vss.n1666 vss.n1645 27.8593
R5746 vss.n3996 vss.n1645 27.8593
R5747 vss.n3997 vss.n3996 27.8593
R5748 vss.n3997 vss.n1633 27.8593
R5749 vss.n4005 vss.n1633 27.8593
R5750 vss.n4006 vss.n4005 27.8593
R5751 vss.n4006 vss.n1621 27.8593
R5752 vss.n4014 vss.n1621 27.8593
R5753 vss.n4015 vss.n4014 27.8593
R5754 vss.n4015 vss.n1599 27.8593
R5755 vss.n4023 vss.n1599 27.8593
R5756 vss.n4024 vss.n4023 27.8593
R5757 vss.n4024 vss.n1587 27.8593
R5758 vss.n4032 vss.n1587 27.8593
R5759 vss.n4033 vss.n4032 27.8593
R5760 vss.n4033 vss.n1575 27.8593
R5761 vss.n4041 vss.n1575 27.8593
R5762 vss.n4042 vss.n4041 27.8593
R5763 vss.n4042 vss.n1563 27.8593
R5764 vss.n4050 vss.n1563 27.8593
R5765 vss.n4051 vss.n4050 27.8593
R5766 vss.n4051 vss.n1540 27.8593
R5767 vss.n4059 vss.n1540 27.8593
R5768 vss.n4060 vss.n4059 27.8593
R5769 vss.n4060 vss.n1528 27.8593
R5770 vss.n4068 vss.n1528 27.8593
R5771 vss.n4069 vss.n4068 27.8593
R5772 vss.n4069 vss.n1516 27.8593
R5773 vss.n4077 vss.n1516 27.8593
R5774 vss.n4078 vss.n4077 27.8593
R5775 vss.n4078 vss.n1504 27.8593
R5776 vss.n4086 vss.n1504 27.8593
R5777 vss.n4087 vss.n4086 27.8593
R5778 vss.n4087 vss.n1499 27.8593
R5779 vss.n1499 vss.n1478 27.8593
R5780 vss.n4098 vss.n1478 27.8593
R5781 vss.n4099 vss.n4098 27.8593
R5782 vss.n4099 vss.n1466 27.8593
R5783 vss.n4107 vss.n1466 27.8593
R5784 vss.n4108 vss.n4107 27.8593
R5785 vss.n4108 vss.n1454 27.8593
R5786 vss.n4116 vss.n1454 27.8593
R5787 vss.n4117 vss.n4116 27.8593
R5788 vss.n4117 vss.n1432 27.8593
R5789 vss.n4125 vss.n1432 27.8593
R5790 vss.n4126 vss.n4125 27.8593
R5791 vss.n4126 vss.n1420 27.8593
R5792 vss.n4134 vss.n1420 27.8593
R5793 vss.n4135 vss.n4134 27.8593
R5794 vss.n4135 vss.n1408 27.8593
R5795 vss.n4143 vss.n1408 27.8593
R5796 vss.n4144 vss.n4143 27.8593
R5797 vss.n4144 vss.n1396 27.8593
R5798 vss.n4152 vss.n1396 27.8593
R5799 vss.n4153 vss.n4152 27.8593
R5800 vss.n4153 vss.n1384 27.8593
R5801 vss.n4161 vss.n1384 27.8593
R5802 vss.n4162 vss.n4161 27.8593
R5803 vss.n4162 vss.n1372 27.8593
R5804 vss.n4170 vss.n1372 27.8593
R5805 vss.n4171 vss.n4170 27.8593
R5806 vss.n4171 vss.n1360 27.8593
R5807 vss.n4179 vss.n1360 27.8593
R5808 vss.n4180 vss.n4179 27.8593
R5809 vss.n4180 vss.n1349 27.8593
R5810 vss.n4188 vss.n1349 27.8593
R5811 vss.n4189 vss.n4188 27.8593
R5812 vss.n4189 vss.n1336 27.8593
R5813 vss.n4197 vss.n1336 27.8593
R5814 vss.n4198 vss.n4197 27.8593
R5815 vss.n4198 vss.n1327 27.8593
R5816 vss.n2965 vss.n1327 27.8593
R5817 vss.n2999 vss.n2965 27.8593
R5818 vss.n3000 vss.n2999 27.8593
R5819 vss.n3000 vss.n2345 27.8593
R5820 vss.n2960 vss.n2345 27.8593
R5821 vss.n2960 vss.n2959 27.8593
R5822 vss.n2959 vss.n2354 27.8593
R5823 vss.n2952 vss.n2354 27.8593
R5824 vss.n2952 vss.n2951 27.8593
R5825 vss.n2951 vss.n2950 27.8593
R5826 vss.n2950 vss.n2366 27.8593
R5827 vss.n2942 vss.n2366 27.8593
R5828 vss.n2942 vss.n2941 27.8593
R5829 vss.n2941 vss.n2467 27.8593
R5830 vss.n2933 vss.n2467 27.8593
R5831 vss.n2933 vss.n2932 27.8593
R5832 vss.n2932 vss.n2478 27.8593
R5833 vss.n2924 vss.n2478 27.8593
R5834 vss.n2924 vss.n2923 27.8593
R5835 vss.n2923 vss.n2494 27.8593
R5836 vss.n2917 vss.n2494 27.8593
R5837 vss.n2917 vss.n2916 27.8593
R5838 vss.n2916 vss.n2508 27.8593
R5839 vss.n2908 vss.n2508 27.8593
R5840 vss.n2908 vss.n2907 27.8593
R5841 vss.n2907 vss.n2523 27.8593
R5842 vss.n2900 vss.n2523 27.8593
R5843 vss.n2900 vss.n2899 27.8593
R5844 vss.n2899 vss.n2536 27.8593
R5845 vss.n2891 vss.n2536 27.8593
R5846 vss.n2891 vss.n2890 27.8593
R5847 vss.n2890 vss.n2550 27.8593
R5848 vss.n2884 vss.n2550 27.8593
R5849 vss.n2884 vss.n2883 27.8593
R5850 vss.n2883 vss.n2567 27.8593
R5851 vss.n2876 vss.n2567 27.8593
R5852 vss.n2876 vss.n2875 27.8593
R5853 vss.n2875 vss.n2579 27.8593
R5854 vss.n2867 vss.n2579 27.8593
R5855 vss.n2867 vss.n2866 27.8593
R5856 vss.n2866 vss.n2595 27.8593
R5857 vss.n2858 vss.n2595 27.8593
R5858 vss.n2858 vss.n2857 27.8593
R5859 vss.n2857 vss.n2856 27.8593
R5860 vss.n2856 vss.n2612 27.8593
R5861 vss.n2848 vss.n2612 27.8593
R5862 vss.n2848 vss.n2847 27.8593
R5863 vss.n2847 vss.n2628 27.8593
R5864 vss.n2839 vss.n2628 27.8593
R5865 vss.n2839 vss.n2838 27.8593
R5866 vss.n2838 vss.n2645 27.8593
R5867 vss.n2831 vss.n2645 27.8593
R5868 vss.n2831 vss.n2830 27.8593
R5869 vss.n2830 vss.n2658 27.8593
R5870 vss.n2824 vss.n2658 27.8593
R5871 vss.n2824 vss.n2823 27.8593
R5872 vss.n2823 vss.n2673 27.8593
R5873 vss.n2816 vss.n2673 27.8593
R5874 vss.n2816 vss.n2815 27.8593
R5875 vss.n2815 vss.n2690 27.8593
R5876 vss.n2807 vss.n2690 27.8593
R5877 vss.n2807 vss.n2806 27.8593
R5878 vss.n2806 vss.n2703 27.8593
R5879 vss.n2798 vss.n2703 27.8593
R5880 vss.n2798 vss.n2797 27.8593
R5881 vss.n2797 vss.n2719 27.8593
R5882 vss.n2791 vss.n2719 27.8593
R5883 vss.n2791 vss.n2790 27.8593
R5884 vss.n2790 vss.n2733 27.8593
R5885 vss.n2782 vss.n2733 27.8593
R5886 vss.n2782 vss.n2781 27.8593
R5887 vss.n2781 vss.n2749 27.8593
R5888 vss.n2773 vss.n2749 27.8593
R5889 vss.n2773 vss.n2772 27.8593
R5890 vss.n2772 vss.n2765 27.8593
R5891 vss.n2765 vss.n206 27.8593
R5892 vss.n5925 vss.n206 27.8593
R5893 vss.n5926 vss.n5925 27.8593
R5894 vss.n5926 vss.n196 27.8593
R5895 vss.n5934 vss.n196 27.8593
R5896 vss.n5935 vss.n5934 27.8593
R5897 vss.n5935 vss.n186 27.8593
R5898 vss.n5943 vss.n186 27.8593
R5899 vss.n5944 vss.n5943 27.8593
R5900 vss.n5944 vss.n174 27.8593
R5901 vss.n5952 vss.n174 27.8593
R5902 vss.n5953 vss.n5952 27.8593
R5903 vss.n5953 vss.n169 27.8593
R5904 vss.n169 vss.n157 27.8593
R5905 vss.n5964 vss.n157 27.8593
R5906 vss.n5965 vss.n5964 27.8593
R5907 vss.n5965 vss.n145 27.8593
R5908 vss.n5997 vss.n145 27.8593
R5909 vss.n5997 vss.n5996 27.8593
R5910 vss.n5996 vss.n5971 27.8593
R5911 vss.n5989 vss.n5971 27.8593
R5912 vss.n5989 vss.n5988 27.8593
R5913 vss.n5988 vss.n134 27.8593
R5914 vss.n6010 vss.n134 27.8593
R5915 vss.n3604 vss.n3080 27.8593
R5916 vss.n3080 vss.n3076 27.8593
R5917 vss.n3076 vss.n3075 27.8593
R5918 vss.n3075 vss.n3072 27.8593
R5919 vss.n3072 vss.n3069 27.8593
R5920 vss.n3069 vss.n3066 27.8593
R5921 vss.n3066 vss.n3063 27.8593
R5922 vss.n3063 vss.n3060 27.8593
R5923 vss.n3060 vss.n3057 27.8593
R5924 vss.n3057 vss.n3054 27.8593
R5925 vss.n3054 vss.n3051 27.8593
R5926 vss.n3051 vss.n3042 27.8593
R5927 vss.n3645 vss.n3042 27.8593
R5928 vss.n3646 vss.n3645 27.8593
R5929 vss.n3646 vss.n2191 27.8593
R5930 vss.n2191 vss.n2187 27.8593
R5931 vss.n2187 vss.n2183 27.8593
R5932 vss.n2183 vss.n2179 27.8593
R5933 vss.n2179 vss.n2175 27.8593
R5934 vss.n2175 vss.n2171 27.8593
R5935 vss.n2171 vss.n2167 27.8593
R5936 vss.n2167 vss.n2163 27.8593
R5937 vss.n2163 vss.n2159 27.8593
R5938 vss.n2159 vss.n2154 27.8593
R5939 vss.n2154 vss.n2151 27.8593
R5940 vss.n2151 vss.n2147 27.8593
R5941 vss.n2147 vss.n2143 27.8593
R5942 vss.n2143 vss.n2139 27.8593
R5943 vss.n2139 vss.n2135 27.8593
R5944 vss.n2135 vss.n2131 27.8593
R5945 vss.n2131 vss.n2127 27.8593
R5946 vss.n2127 vss.n2123 27.8593
R5947 vss.n2123 vss.n2119 27.8593
R5948 vss.n2119 vss.n2115 27.8593
R5949 vss.n2115 vss.n2104 27.8593
R5950 vss.n3714 vss.n2104 27.8593
R5951 vss.n3715 vss.n3714 27.8593
R5952 vss.n3715 vss.n2089 27.8593
R5953 vss.n2089 vss.n2085 27.8593
R5954 vss.n2085 vss.n2081 27.8593
R5955 vss.n2081 vss.n2077 27.8593
R5956 vss.n2077 vss.n2073 27.8593
R5957 vss.n2073 vss.n2069 27.8593
R5958 vss.n2069 vss.n2065 27.8593
R5959 vss.n2065 vss.n2061 27.8593
R5960 vss.n2061 vss.n2050 27.8593
R5961 vss.n3747 vss.n2050 27.8593
R5962 vss.n3748 vss.n3747 27.8593
R5963 vss.n3748 vss.n2035 27.8593
R5964 vss.n2035 vss.n2031 27.8593
R5965 vss.n2031 vss.n2027 27.8593
R5966 vss.n2027 vss.n2023 27.8593
R5967 vss.n2023 vss.n2019 27.8593
R5968 vss.n2019 vss.n2015 27.8593
R5969 vss.n2015 vss.n2011 27.8593
R5970 vss.n2011 vss.n2007 27.8593
R5971 vss.n2007 vss.n2003 27.8593
R5972 vss.n2003 vss.n1998 27.8593
R5973 vss.n1998 vss.n1995 27.8593
R5974 vss.n1995 vss.n1980 27.8593
R5975 vss.n1980 vss.n1976 27.8593
R5976 vss.n1976 vss.n1972 27.8593
R5977 vss.n1972 vss.n1968 27.8593
R5978 vss.n1968 vss.n1964 27.8593
R5979 vss.n1964 vss.n1960 27.8593
R5980 vss.n1960 vss.n1956 27.8593
R5981 vss.n1956 vss.n1952 27.8593
R5982 vss.n1952 vss.n1948 27.8593
R5983 vss.n1948 vss.n1937 27.8593
R5984 vss.n3816 vss.n1937 27.8593
R5985 vss.n3817 vss.n3816 27.8593
R5986 vss.n3817 vss.n1922 27.8593
R5987 vss.n1922 vss.n1918 27.8593
R5988 vss.n1918 vss.n1914 27.8593
R5989 vss.n1914 vss.n1910 27.8593
R5990 vss.n1910 vss.n1906 27.8593
R5991 vss.n1906 vss.n1902 27.8593
R5992 vss.n1902 vss.n1898 27.8593
R5993 vss.n1898 vss.n1894 27.8593
R5994 vss.n1894 vss.n1883 27.8593
R5995 vss.n3849 vss.n1883 27.8593
R5996 vss.n3850 vss.n3849 27.8593
R5997 vss.n3850 vss.n1868 27.8593
R5998 vss.n1868 vss.n1864 27.8593
R5999 vss.n1864 vss.n1860 27.8593
R6000 vss.n1860 vss.n1856 27.8593
R6001 vss.n1856 vss.n1852 27.8593
R6002 vss.n1852 vss.n1848 27.8593
R6003 vss.n1848 vss.n1844 27.8593
R6004 vss.n1844 vss.n1840 27.8593
R6005 vss.n1840 vss.n1836 27.8593
R6006 vss.n1836 vss.n1831 27.8593
R6007 vss.n1831 vss.n1828 27.8593
R6008 vss.n1828 vss.n1813 27.8593
R6009 vss.n1813 vss.n1809 27.8593
R6010 vss.n1809 vss.n1805 27.8593
R6011 vss.n1805 vss.n1801 27.8593
R6012 vss.n1801 vss.n1797 27.8593
R6013 vss.n1797 vss.n1793 27.8593
R6014 vss.n1793 vss.n1789 27.8593
R6015 vss.n1789 vss.n1785 27.8593
R6016 vss.n1785 vss.n1781 27.8593
R6017 vss.n1781 vss.n1770 27.8593
R6018 vss.n3918 vss.n1770 27.8593
R6019 vss.n3919 vss.n3918 27.8593
R6020 vss.n3919 vss.n1765 27.8593
R6021 vss.n1765 vss.n1761 27.8593
R6022 vss.n1761 vss.n1757 27.8593
R6023 vss.n1757 vss.n1753 27.8593
R6024 vss.n1753 vss.n1749 27.8593
R6025 vss.n1749 vss.n1745 27.8593
R6026 vss.n1745 vss.n1741 27.8593
R6027 vss.n1741 vss.n1737 27.8593
R6028 vss.n1737 vss.n1733 27.8593
R6029 vss.n1733 vss.n1728 27.8593
R6030 vss.n1728 vss.n1725 27.8593
R6031 vss.n1725 vss.n1710 27.8593
R6032 vss.n1710 vss.n1706 27.8593
R6033 vss.n1706 vss.n1702 27.8593
R6034 vss.n1702 vss.n1698 27.8593
R6035 vss.n1698 vss.n1694 27.8593
R6036 vss.n1694 vss.n1690 27.8593
R6037 vss.n1690 vss.n1686 27.8593
R6038 vss.n1686 vss.n1682 27.8593
R6039 vss.n1682 vss.n1678 27.8593
R6040 vss.n1678 vss.n1667 27.8593
R6041 vss.n3987 vss.n1667 27.8593
R6042 vss.n3988 vss.n3987 27.8593
R6043 vss.n3988 vss.n1652 27.8593
R6044 vss.n1652 vss.n1648 27.8593
R6045 vss.n1648 vss.n1644 27.8593
R6046 vss.n1644 vss.n1640 27.8593
R6047 vss.n1640 vss.n1636 27.8593
R6048 vss.n1636 vss.n1632 27.8593
R6049 vss.n1632 vss.n1628 27.8593
R6050 vss.n1628 vss.n1624 27.8593
R6051 vss.n1624 vss.n1613 27.8593
R6052 vss.n4020 vss.n1613 27.8593
R6053 vss.n4021 vss.n4020 27.8593
R6054 vss.n4021 vss.n1598 27.8593
R6055 vss.n1598 vss.n1594 27.8593
R6056 vss.n1594 vss.n1590 27.8593
R6057 vss.n1590 vss.n1586 27.8593
R6058 vss.n1586 vss.n1582 27.8593
R6059 vss.n1582 vss.n1578 27.8593
R6060 vss.n1578 vss.n1574 27.8593
R6061 vss.n1574 vss.n1570 27.8593
R6062 vss.n1570 vss.n1566 27.8593
R6063 vss.n1566 vss.n1561 27.8593
R6064 vss.n1561 vss.n1558 27.8593
R6065 vss.n1558 vss.n1543 27.8593
R6066 vss.n1543 vss.n1539 27.8593
R6067 vss.n1539 vss.n1535 27.8593
R6068 vss.n1535 vss.n1531 27.8593
R6069 vss.n1531 vss.n1527 27.8593
R6070 vss.n1527 vss.n1523 27.8593
R6071 vss.n1523 vss.n1519 27.8593
R6072 vss.n1519 vss.n1515 27.8593
R6073 vss.n1515 vss.n1511 27.8593
R6074 vss.n1511 vss.n1500 27.8593
R6075 vss.n4089 vss.n1500 27.8593
R6076 vss.n4090 vss.n4089 27.8593
R6077 vss.n4090 vss.n1485 27.8593
R6078 vss.n1485 vss.n1481 27.8593
R6079 vss.n1481 vss.n1477 27.8593
R6080 vss.n1477 vss.n1473 27.8593
R6081 vss.n1473 vss.n1469 27.8593
R6082 vss.n1469 vss.n1465 27.8593
R6083 vss.n1465 vss.n1461 27.8593
R6084 vss.n1461 vss.n1457 27.8593
R6085 vss.n1457 vss.n1446 27.8593
R6086 vss.n4122 vss.n1446 27.8593
R6087 vss.n4123 vss.n4122 27.8593
R6088 vss.n4123 vss.n1431 27.8593
R6089 vss.n1431 vss.n1427 27.8593
R6090 vss.n1427 vss.n1423 27.8593
R6091 vss.n1423 vss.n1419 27.8593
R6092 vss.n1419 vss.n1415 27.8593
R6093 vss.n1415 vss.n1411 27.8593
R6094 vss.n1411 vss.n1407 27.8593
R6095 vss.n1407 vss.n1403 27.8593
R6096 vss.n1403 vss.n1399 27.8593
R6097 vss.n1399 vss.n1394 27.8593
R6098 vss.n1394 vss.n1391 27.8593
R6099 vss.n1391 vss.n1387 27.8593
R6100 vss.n1387 vss.n1383 27.8593
R6101 vss.n1383 vss.n1379 27.8593
R6102 vss.n1379 vss.n1375 27.8593
R6103 vss.n1375 vss.n1371 27.8593
R6104 vss.n1371 vss.n1367 27.8593
R6105 vss.n1367 vss.n1363 27.8593
R6106 vss.n1363 vss.n1359 27.8593
R6107 vss.n1359 vss.n1356 27.8593
R6108 vss.n1356 vss.n1352 27.8593
R6109 vss.n1352 vss.n1347 27.8593
R6110 vss.n1347 vss.n1344 27.8593
R6111 vss.n1344 vss.n1339 27.8593
R6112 vss.n1339 vss.n1334 27.8593
R6113 vss.n1334 vss.n1330 27.8593
R6114 vss.n2994 vss.n1330 27.8593
R6115 vss.n2994 vss.n2992 27.8593
R6116 vss.n2992 vss.n2963 27.8593
R6117 vss.n2963 vss.n2348 27.8593
R6118 vss.n2351 vss.n2348 27.8593
R6119 vss.n2355 vss.n2351 27.8593
R6120 vss.n2358 vss.n2355 27.8593
R6121 vss.n2360 vss.n2358 27.8593
R6122 vss.n2367 vss.n2360 27.8593
R6123 vss.n2368 vss.n2367 27.8593
R6124 vss.n2459 vss.n2368 27.8593
R6125 vss.n2464 vss.n2459 27.8593
R6126 vss.n2468 vss.n2464 27.8593
R6127 vss.n2471 vss.n2468 27.8593
R6128 vss.n2476 vss.n2471 27.8593
R6129 vss.n2479 vss.n2476 27.8593
R6130 vss.n2486 vss.n2479 27.8593
R6131 vss.n2489 vss.n2486 27.8593
R6132 vss.n2495 vss.n2489 27.8593
R6133 vss.n2502 vss.n2495 27.8593
R6134 vss.n2503 vss.n2502 27.8593
R6135 vss.n2509 vss.n2503 27.8593
R6136 vss.n2515 vss.n2509 27.8593
R6137 vss.n2518 vss.n2515 27.8593
R6138 vss.n2524 vss.n2518 27.8593
R6139 vss.n2526 vss.n2524 27.8593
R6140 vss.n2533 vss.n2526 27.8593
R6141 vss.n2537 vss.n2533 27.8593
R6142 vss.n2540 vss.n2537 27.8593
R6143 vss.n2548 vss.n2540 27.8593
R6144 vss.n2551 vss.n2548 27.8593
R6145 vss.n2553 vss.n2551 27.8593
R6146 vss.n2561 vss.n2553 27.8593
R6147 vss.n2568 vss.n2561 27.8593
R6148 vss.n2570 vss.n2568 27.8593
R6149 vss.n2576 vss.n2570 27.8593
R6150 vss.n2580 vss.n2576 27.8593
R6151 vss.n2586 vss.n2580 27.8593
R6152 vss.n2590 vss.n2586 27.8593
R6153 vss.n2596 vss.n2590 27.8593
R6154 vss.n2599 vss.n2596 27.8593
R6155 vss.n2605 vss.n2599 27.8593
R6156 vss.n2614 vss.n2605 27.8593
R6157 vss.n2615 vss.n2614 27.8593
R6158 vss.n2620 vss.n2615 27.8593
R6159 vss.n2626 vss.n2620 27.8593
R6160 vss.n2629 vss.n2626 27.8593
R6161 vss.n2636 vss.n2629 27.8593
R6162 vss.n2639 vss.n2636 27.8593
R6163 vss.n2646 vss.n2639 27.8593
R6164 vss.n2649 vss.n2646 27.8593
R6165 vss.n2651 vss.n2649 27.8593
R6166 vss.n2659 vss.n2651 27.8593
R6167 vss.n2668 vss.n2659 27.8593
R6168 vss.n2669 vss.n2668 27.8593
R6169 vss.n2674 vss.n2669 27.8593
R6170 vss.n2676 vss.n2674 27.8593
R6171 vss.n2684 vss.n2676 27.8593
R6172 vss.n2691 vss.n2684 27.8593
R6173 vss.n2694 vss.n2691 27.8593
R6174 vss.n2701 vss.n2694 27.8593
R6175 vss.n2704 vss.n2701 27.8593
R6176 vss.n2710 vss.n2704 27.8593
R6177 vss.n2713 vss.n2710 27.8593
R6178 vss.n2720 vss.n2713 27.8593
R6179 vss.n2722 vss.n2720 27.8593
R6180 vss.n2730 vss.n2722 27.8593
R6181 vss.n2734 vss.n2730 27.8593
R6182 vss.n2740 vss.n2734 27.8593
R6183 vss.n2744 vss.n2740 27.8593
R6184 vss.n2750 vss.n2744 27.8593
R6185 vss.n2753 vss.n2750 27.8593
R6186 vss.n2759 vss.n2753 27.8593
R6187 vss.n2766 vss.n2759 27.8593
R6188 vss.n2767 vss.n2766 27.8593
R6189 vss.n2767 vss.n212 27.8593
R6190 vss.n212 vss.n209 27.8593
R6191 vss.n209 vss.n205 27.8593
R6192 vss.n205 vss.n202 27.8593
R6193 vss.n202 vss.n198 27.8593
R6194 vss.n198 vss.n195 27.8593
R6195 vss.n195 vss.n192 27.8593
R6196 vss.n192 vss.n188 27.8593
R6197 vss.n188 vss.n185 27.8593
R6198 vss.n185 vss.n181 27.8593
R6199 vss.n181 vss.n170 27.8593
R6200 vss.n5955 vss.n170 27.8593
R6201 vss.n5956 vss.n5955 27.8593
R6202 vss.n5956 vss.n165 27.8593
R6203 vss.n165 vss.n160 27.8593
R6204 vss.n160 vss.n155 27.8593
R6205 vss.n155 vss.n147 27.8593
R6206 vss.n5968 vss.n147 27.8593
R6207 vss.n5972 vss.n5968 27.8593
R6208 vss.n5976 vss.n5972 27.8593
R6209 vss.n5978 vss.n5976 27.8593
R6210 vss.n5982 vss.n5978 27.8593
R6211 vss.n5982 vss.n5981 27.8593
R6212 vss.n5981 vss.n131 27.8593
R6213 vss.n3610 vss.n3078 27.8593
R6214 vss.n3612 vss.n3610 27.8593
R6215 vss.n3612 vss.n3611 27.8593
R6216 vss.n3611 vss.n3067 27.8593
R6217 vss.n3621 vss.n3067 27.8593
R6218 vss.n3622 vss.n3621 27.8593
R6219 vss.n3622 vss.n3058 27.8593
R6220 vss.n3630 vss.n3058 27.8593
R6221 vss.n3631 vss.n3630 27.8593
R6222 vss.n3631 vss.n3049 27.8593
R6223 vss.n3639 vss.n3049 27.8593
R6224 vss.n3640 vss.n3639 27.8593
R6225 vss.n3640 vss.n2192 27.8593
R6226 vss.n3648 vss.n2192 27.8593
R6227 vss.n3649 vss.n3648 27.8593
R6228 vss.n3649 vss.n2180 27.8593
R6229 vss.n3657 vss.n2180 27.8593
R6230 vss.n3658 vss.n3657 27.8593
R6231 vss.n3658 vss.n2168 27.8593
R6232 vss.n3666 vss.n2168 27.8593
R6233 vss.n3667 vss.n3666 27.8593
R6234 vss.n3667 vss.n2156 27.8593
R6235 vss.n3675 vss.n2156 27.8593
R6236 vss.n3676 vss.n3675 27.8593
R6237 vss.n3676 vss.n2144 27.8593
R6238 vss.n3684 vss.n2144 27.8593
R6239 vss.n3685 vss.n3684 27.8593
R6240 vss.n3685 vss.n2132 27.8593
R6241 vss.n3693 vss.n2132 27.8593
R6242 vss.n3694 vss.n3693 27.8593
R6243 vss.n3694 vss.n2120 27.8593
R6244 vss.n3702 vss.n2120 27.8593
R6245 vss.n3703 vss.n3702 27.8593
R6246 vss.n3703 vss.n2108 27.8593
R6247 vss.n3711 vss.n2108 27.8593
R6248 vss.n3712 vss.n3711 27.8593
R6249 vss.n3712 vss.n2103 27.8593
R6250 vss.n2103 vss.n2082 27.8593
R6251 vss.n3723 vss.n2082 27.8593
R6252 vss.n3724 vss.n3723 27.8593
R6253 vss.n3724 vss.n2070 27.8593
R6254 vss.n3732 vss.n2070 27.8593
R6255 vss.n3733 vss.n3732 27.8593
R6256 vss.n3733 vss.n2058 27.8593
R6257 vss.n3741 vss.n2058 27.8593
R6258 vss.n3742 vss.n3741 27.8593
R6259 vss.n3742 vss.n2036 27.8593
R6260 vss.n3750 vss.n2036 27.8593
R6261 vss.n3751 vss.n3750 27.8593
R6262 vss.n3751 vss.n2024 27.8593
R6263 vss.n3759 vss.n2024 27.8593
R6264 vss.n3760 vss.n3759 27.8593
R6265 vss.n3760 vss.n2012 27.8593
R6266 vss.n3768 vss.n2012 27.8593
R6267 vss.n3769 vss.n3768 27.8593
R6268 vss.n3769 vss.n2000 27.8593
R6269 vss.n3777 vss.n2000 27.8593
R6270 vss.n3778 vss.n3777 27.8593
R6271 vss.n3778 vss.n1977 27.8593
R6272 vss.n3786 vss.n1977 27.8593
R6273 vss.n3787 vss.n3786 27.8593
R6274 vss.n3787 vss.n1965 27.8593
R6275 vss.n3795 vss.n1965 27.8593
R6276 vss.n3796 vss.n3795 27.8593
R6277 vss.n3796 vss.n1953 27.8593
R6278 vss.n3804 vss.n1953 27.8593
R6279 vss.n3805 vss.n3804 27.8593
R6280 vss.n3805 vss.n1941 27.8593
R6281 vss.n3813 vss.n1941 27.8593
R6282 vss.n3814 vss.n3813 27.8593
R6283 vss.n3814 vss.n1936 27.8593
R6284 vss.n1936 vss.n1915 27.8593
R6285 vss.n3825 vss.n1915 27.8593
R6286 vss.n3826 vss.n3825 27.8593
R6287 vss.n3826 vss.n1903 27.8593
R6288 vss.n3834 vss.n1903 27.8593
R6289 vss.n3835 vss.n3834 27.8593
R6290 vss.n3835 vss.n1891 27.8593
R6291 vss.n3843 vss.n1891 27.8593
R6292 vss.n3844 vss.n3843 27.8593
R6293 vss.n3844 vss.n1869 27.8593
R6294 vss.n3852 vss.n1869 27.8593
R6295 vss.n3853 vss.n3852 27.8593
R6296 vss.n3853 vss.n1857 27.8593
R6297 vss.n3861 vss.n1857 27.8593
R6298 vss.n3862 vss.n3861 27.8593
R6299 vss.n3862 vss.n1845 27.8593
R6300 vss.n3870 vss.n1845 27.8593
R6301 vss.n3871 vss.n3870 27.8593
R6302 vss.n3871 vss.n1833 27.8593
R6303 vss.n3879 vss.n1833 27.8593
R6304 vss.n3880 vss.n3879 27.8593
R6305 vss.n3880 vss.n1810 27.8593
R6306 vss.n3888 vss.n1810 27.8593
R6307 vss.n3889 vss.n3888 27.8593
R6308 vss.n3889 vss.n1798 27.8593
R6309 vss.n3897 vss.n1798 27.8593
R6310 vss.n3898 vss.n3897 27.8593
R6311 vss.n3898 vss.n1786 27.8593
R6312 vss.n3906 vss.n1786 27.8593
R6313 vss.n3907 vss.n3906 27.8593
R6314 vss.n3907 vss.n1774 27.8593
R6315 vss.n3915 vss.n1774 27.8593
R6316 vss.n3916 vss.n3915 27.8593
R6317 vss.n3916 vss.n1769 27.8593
R6318 vss.n1769 vss.n1758 27.8593
R6319 vss.n3927 vss.n1758 27.8593
R6320 vss.n3928 vss.n3927 27.8593
R6321 vss.n3928 vss.n1746 27.8593
R6322 vss.n3936 vss.n1746 27.8593
R6323 vss.n3937 vss.n3936 27.8593
R6324 vss.n3937 vss.n1734 27.8593
R6325 vss.n3945 vss.n1734 27.8593
R6326 vss.n3946 vss.n3945 27.8593
R6327 vss.n3946 vss.n1711 27.8593
R6328 vss.n3954 vss.n1711 27.8593
R6329 vss.n3955 vss.n3954 27.8593
R6330 vss.n3955 vss.n1699 27.8593
R6331 vss.n3963 vss.n1699 27.8593
R6332 vss.n3964 vss.n3963 27.8593
R6333 vss.n3964 vss.n1687 27.8593
R6334 vss.n3972 vss.n1687 27.8593
R6335 vss.n3973 vss.n3972 27.8593
R6336 vss.n3973 vss.n1675 27.8593
R6337 vss.n3981 vss.n1675 27.8593
R6338 vss.n3982 vss.n3981 27.8593
R6339 vss.n3982 vss.n1653 27.8593
R6340 vss.n3990 vss.n1653 27.8593
R6341 vss.n3991 vss.n3990 27.8593
R6342 vss.n3991 vss.n1641 27.8593
R6343 vss.n3999 vss.n1641 27.8593
R6344 vss.n4000 vss.n3999 27.8593
R6345 vss.n4000 vss.n1629 27.8593
R6346 vss.n4008 vss.n1629 27.8593
R6347 vss.n4009 vss.n4008 27.8593
R6348 vss.n4009 vss.n1617 27.8593
R6349 vss.n4017 vss.n1617 27.8593
R6350 vss.n4018 vss.n4017 27.8593
R6351 vss.n4018 vss.n1612 27.8593
R6352 vss.n1612 vss.n1591 27.8593
R6353 vss.n4029 vss.n1591 27.8593
R6354 vss.n4030 vss.n4029 27.8593
R6355 vss.n4030 vss.n1579 27.8593
R6356 vss.n4038 vss.n1579 27.8593
R6357 vss.n4039 vss.n4038 27.8593
R6358 vss.n4039 vss.n1567 27.8593
R6359 vss.n4047 vss.n1567 27.8593
R6360 vss.n4048 vss.n4047 27.8593
R6361 vss.n4048 vss.n1544 27.8593
R6362 vss.n4056 vss.n1544 27.8593
R6363 vss.n4057 vss.n4056 27.8593
R6364 vss.n4057 vss.n1532 27.8593
R6365 vss.n4065 vss.n1532 27.8593
R6366 vss.n4066 vss.n4065 27.8593
R6367 vss.n4066 vss.n1520 27.8593
R6368 vss.n4074 vss.n1520 27.8593
R6369 vss.n4075 vss.n4074 27.8593
R6370 vss.n4075 vss.n1508 27.8593
R6371 vss.n4083 vss.n1508 27.8593
R6372 vss.n4084 vss.n4083 27.8593
R6373 vss.n4084 vss.n1486 27.8593
R6374 vss.n4092 vss.n1486 27.8593
R6375 vss.n4093 vss.n4092 27.8593
R6376 vss.n4093 vss.n1474 27.8593
R6377 vss.n4101 vss.n1474 27.8593
R6378 vss.n4102 vss.n4101 27.8593
R6379 vss.n4102 vss.n1462 27.8593
R6380 vss.n4110 vss.n1462 27.8593
R6381 vss.n4111 vss.n4110 27.8593
R6382 vss.n4111 vss.n1450 27.8593
R6383 vss.n4119 vss.n1450 27.8593
R6384 vss.n4120 vss.n4119 27.8593
R6385 vss.n4120 vss.n1445 27.8593
R6386 vss.n1445 vss.n1424 27.8593
R6387 vss.n4131 vss.n1424 27.8593
R6388 vss.n4132 vss.n4131 27.8593
R6389 vss.n4132 vss.n1412 27.8593
R6390 vss.n4140 vss.n1412 27.8593
R6391 vss.n4141 vss.n4140 27.8593
R6392 vss.n4141 vss.n1400 27.8593
R6393 vss.n4149 vss.n1400 27.8593
R6394 vss.n4150 vss.n4149 27.8593
R6395 vss.n4150 vss.n1388 27.8593
R6396 vss.n4158 vss.n1388 27.8593
R6397 vss.n4159 vss.n4158 27.8593
R6398 vss.n4159 vss.n1376 27.8593
R6399 vss.n4167 vss.n1376 27.8593
R6400 vss.n4168 vss.n4167 27.8593
R6401 vss.n4168 vss.n1364 27.8593
R6402 vss.n4176 vss.n1364 27.8593
R6403 vss.n4177 vss.n4176 27.8593
R6404 vss.n4177 vss.n1353 27.8593
R6405 vss.n4185 vss.n1353 27.8593
R6406 vss.n4186 vss.n4185 27.8593
R6407 vss.n4186 vss.n1341 27.8593
R6408 vss.n4194 vss.n1341 27.8593
R6409 vss.n4195 vss.n4194 27.8593
R6410 vss.n4195 vss.n1335 27.8593
R6411 vss.n1335 vss.n1328 27.8593
R6412 vss.n2996 vss.n1328 27.8593
R6413 vss.n2997 vss.n2996 27.8593
R6414 vss.n2997 vss.n2964 27.8593
R6415 vss.n2964 vss.n2346 27.8593
R6416 vss.n2352 vss.n2346 27.8593
R6417 vss.n2957 vss.n2352 27.8593
R6418 vss.n2957 vss.n2956 27.8593
R6419 vss.n2956 vss.n2357 27.8593
R6420 vss.n2371 vss.n2357 27.8593
R6421 vss.n2948 vss.n2371 27.8593
R6422 vss.n2948 vss.n2947 27.8593
R6423 vss.n2947 vss.n2458 27.8593
R6424 vss.n2939 vss.n2458 27.8593
R6425 vss.n2939 vss.n2938 27.8593
R6426 vss.n2938 vss.n2470 27.8593
R6427 vss.n2930 vss.n2470 27.8593
R6428 vss.n2930 vss.n2929 27.8593
R6429 vss.n2929 vss.n2485 27.8593
R6430 vss.n2921 vss.n2485 27.8593
R6431 vss.n2921 vss.n2920 27.8593
R6432 vss.n2920 vss.n2919 27.8593
R6433 vss.n2919 vss.n2501 27.8593
R6434 vss.n2911 vss.n2501 27.8593
R6435 vss.n2911 vss.n2910 27.8593
R6436 vss.n2910 vss.n2517 27.8593
R6437 vss.n2903 vss.n2517 27.8593
R6438 vss.n2903 vss.n2902 27.8593
R6439 vss.n2902 vss.n2532 27.8593
R6440 vss.n2894 vss.n2532 27.8593
R6441 vss.n2894 vss.n2893 27.8593
R6442 vss.n2893 vss.n2547 27.8593
R6443 vss.n2887 vss.n2547 27.8593
R6444 vss.n2887 vss.n2886 27.8593
R6445 vss.n2886 vss.n2560 27.8593
R6446 vss.n2879 vss.n2560 27.8593
R6447 vss.n2879 vss.n2878 27.8593
R6448 vss.n2878 vss.n2575 27.8593
R6449 vss.n2870 vss.n2575 27.8593
R6450 vss.n2870 vss.n2869 27.8593
R6451 vss.n2869 vss.n2589 27.8593
R6452 vss.n2861 vss.n2589 27.8593
R6453 vss.n2861 vss.n2860 27.8593
R6454 vss.n2860 vss.n2604 27.8593
R6455 vss.n2854 vss.n2604 27.8593
R6456 vss.n2854 vss.n2853 27.8593
R6457 vss.n2853 vss.n2619 27.8593
R6458 vss.n2845 vss.n2619 27.8593
R6459 vss.n2845 vss.n2844 27.8593
R6460 vss.n2844 vss.n2635 27.8593
R6461 vss.n2836 vss.n2635 27.8593
R6462 vss.n2836 vss.n2835 27.8593
R6463 vss.n2835 vss.n2648 27.8593
R6464 vss.n2828 vss.n2648 27.8593
R6465 vss.n2828 vss.n2827 27.8593
R6466 vss.n2827 vss.n2826 27.8593
R6467 vss.n2826 vss.n2667 27.8593
R6468 vss.n2819 vss.n2667 27.8593
R6469 vss.n2819 vss.n2818 27.8593
R6470 vss.n2818 vss.n2683 27.8593
R6471 vss.n2810 vss.n2683 27.8593
R6472 vss.n2810 vss.n2809 27.8593
R6473 vss.n2809 vss.n2700 27.8593
R6474 vss.n2801 vss.n2700 27.8593
R6475 vss.n2801 vss.n2800 27.8593
R6476 vss.n2800 vss.n2712 27.8593
R6477 vss.n2794 vss.n2712 27.8593
R6478 vss.n2794 vss.n2793 27.8593
R6479 vss.n2793 vss.n2729 27.8593
R6480 vss.n2785 vss.n2729 27.8593
R6481 vss.n2785 vss.n2784 27.8593
R6482 vss.n2784 vss.n2743 27.8593
R6483 vss.n2776 vss.n2743 27.8593
R6484 vss.n2776 vss.n2775 27.8593
R6485 vss.n2775 vss.n2758 27.8593
R6486 vss.n2758 vss.n210 27.8593
R6487 vss.n5922 vss.n210 27.8593
R6488 vss.n5923 vss.n5922 27.8593
R6489 vss.n5923 vss.n199 27.8593
R6490 vss.n5931 vss.n199 27.8593
R6491 vss.n5932 vss.n5931 27.8593
R6492 vss.n5932 vss.n189 27.8593
R6493 vss.n5940 vss.n189 27.8593
R6494 vss.n5941 vss.n5940 27.8593
R6495 vss.n5941 vss.n178 27.8593
R6496 vss.n5949 vss.n178 27.8593
R6497 vss.n5950 vss.n5949 27.8593
R6498 vss.n5950 vss.n173 27.8593
R6499 vss.n173 vss.n162 27.8593
R6500 vss.n5961 vss.n162 27.8593
R6501 vss.n5962 vss.n5961 27.8593
R6502 vss.n5962 vss.n156 27.8593
R6503 vss.n156 vss.n146 27.8593
R6504 vss.n5970 vss.n146 27.8593
R6505 vss.n5994 vss.n5970 27.8593
R6506 vss.n5994 vss.n5993 27.8593
R6507 vss.n5993 vss.n5975 27.8593
R6508 vss.n5986 vss.n5975 27.8593
R6509 vss.n5986 vss.n5985 27.8593
R6510 vss.n5985 vss.n133 27.8593
R6511 vss.n3608 vss.n3607 27.8593
R6512 vss.n3608 vss.n3077 27.8593
R6513 vss.n3077 vss.n3070 27.8593
R6514 vss.n3618 vss.n3070 27.8593
R6515 vss.n3619 vss.n3618 27.8593
R6516 vss.n3619 vss.n3061 27.8593
R6517 vss.n3627 vss.n3061 27.8593
R6518 vss.n3628 vss.n3627 27.8593
R6519 vss.n3628 vss.n3052 27.8593
R6520 vss.n3636 vss.n3052 27.8593
R6521 vss.n3637 vss.n3636 27.8593
R6522 vss.n3637 vss.n3048 27.8593
R6523 vss.n3048 vss.n3044 27.8593
R6524 vss.n3044 vss.n2188 27.8593
R6525 vss.n3651 vss.n2188 27.8593
R6526 vss.n3652 vss.n3651 27.8593
R6527 vss.n3652 vss.n2176 27.8593
R6528 vss.n3660 vss.n2176 27.8593
R6529 vss.n3661 vss.n3660 27.8593
R6530 vss.n3661 vss.n2164 27.8593
R6531 vss.n3669 vss.n2164 27.8593
R6532 vss.n3670 vss.n3669 27.8593
R6533 vss.n3670 vss.n2152 27.8593
R6534 vss.n3678 vss.n2152 27.8593
R6535 vss.n3679 vss.n3678 27.8593
R6536 vss.n3679 vss.n2140 27.8593
R6537 vss.n3687 vss.n2140 27.8593
R6538 vss.n3688 vss.n3687 27.8593
R6539 vss.n3688 vss.n2128 27.8593
R6540 vss.n3696 vss.n2128 27.8593
R6541 vss.n3697 vss.n3696 27.8593
R6542 vss.n3697 vss.n2116 27.8593
R6543 vss.n3705 vss.n2116 27.8593
R6544 vss.n3706 vss.n3705 27.8593
R6545 vss.n3706 vss.n2111 27.8593
R6546 vss.n2111 vss.n2106 27.8593
R6547 vss.n2106 vss.n2086 27.8593
R6548 vss.n3720 vss.n2086 27.8593
R6549 vss.n3721 vss.n3720 27.8593
R6550 vss.n3721 vss.n2074 27.8593
R6551 vss.n3729 vss.n2074 27.8593
R6552 vss.n3730 vss.n3729 27.8593
R6553 vss.n3730 vss.n2062 27.8593
R6554 vss.n3738 vss.n2062 27.8593
R6555 vss.n3739 vss.n3738 27.8593
R6556 vss.n3739 vss.n2057 27.8593
R6557 vss.n2057 vss.n2052 27.8593
R6558 vss.n2052 vss.n2032 27.8593
R6559 vss.n3753 vss.n2032 27.8593
R6560 vss.n3754 vss.n3753 27.8593
R6561 vss.n3754 vss.n2020 27.8593
R6562 vss.n3762 vss.n2020 27.8593
R6563 vss.n3763 vss.n3762 27.8593
R6564 vss.n3763 vss.n2008 27.8593
R6565 vss.n3771 vss.n2008 27.8593
R6566 vss.n3772 vss.n3771 27.8593
R6567 vss.n3772 vss.n1996 27.8593
R6568 vss.n3780 vss.n1996 27.8593
R6569 vss.n3781 vss.n3780 27.8593
R6570 vss.n3781 vss.n1973 27.8593
R6571 vss.n3789 vss.n1973 27.8593
R6572 vss.n3790 vss.n3789 27.8593
R6573 vss.n3790 vss.n1961 27.8593
R6574 vss.n3798 vss.n1961 27.8593
R6575 vss.n3799 vss.n3798 27.8593
R6576 vss.n3799 vss.n1949 27.8593
R6577 vss.n3807 vss.n1949 27.8593
R6578 vss.n3808 vss.n3807 27.8593
R6579 vss.n3808 vss.n1944 27.8593
R6580 vss.n1944 vss.n1939 27.8593
R6581 vss.n1939 vss.n1919 27.8593
R6582 vss.n3822 vss.n1919 27.8593
R6583 vss.n3823 vss.n3822 27.8593
R6584 vss.n3823 vss.n1907 27.8593
R6585 vss.n3831 vss.n1907 27.8593
R6586 vss.n3832 vss.n3831 27.8593
R6587 vss.n3832 vss.n1895 27.8593
R6588 vss.n3840 vss.n1895 27.8593
R6589 vss.n3841 vss.n3840 27.8593
R6590 vss.n3841 vss.n1890 27.8593
R6591 vss.n1890 vss.n1885 27.8593
R6592 vss.n1885 vss.n1865 27.8593
R6593 vss.n3855 vss.n1865 27.8593
R6594 vss.n3856 vss.n3855 27.8593
R6595 vss.n3856 vss.n1853 27.8593
R6596 vss.n3864 vss.n1853 27.8593
R6597 vss.n3865 vss.n3864 27.8593
R6598 vss.n3865 vss.n1841 27.8593
R6599 vss.n3873 vss.n1841 27.8593
R6600 vss.n3874 vss.n3873 27.8593
R6601 vss.n3874 vss.n1829 27.8593
R6602 vss.n3882 vss.n1829 27.8593
R6603 vss.n3883 vss.n3882 27.8593
R6604 vss.n3883 vss.n1806 27.8593
R6605 vss.n3891 vss.n1806 27.8593
R6606 vss.n3892 vss.n3891 27.8593
R6607 vss.n3892 vss.n1794 27.8593
R6608 vss.n3900 vss.n1794 27.8593
R6609 vss.n3901 vss.n3900 27.8593
R6610 vss.n3901 vss.n1782 27.8593
R6611 vss.n3909 vss.n1782 27.8593
R6612 vss.n3910 vss.n3909 27.8593
R6613 vss.n3910 vss.n1777 27.8593
R6614 vss.n1777 vss.n1772 27.8593
R6615 vss.n1772 vss.n1762 27.8593
R6616 vss.n3924 vss.n1762 27.8593
R6617 vss.n3925 vss.n3924 27.8593
R6618 vss.n3925 vss.n1750 27.8593
R6619 vss.n3933 vss.n1750 27.8593
R6620 vss.n3934 vss.n3933 27.8593
R6621 vss.n3934 vss.n1738 27.8593
R6622 vss.n3942 vss.n1738 27.8593
R6623 vss.n3943 vss.n3942 27.8593
R6624 vss.n3943 vss.n1726 27.8593
R6625 vss.n3951 vss.n1726 27.8593
R6626 vss.n3952 vss.n3951 27.8593
R6627 vss.n3952 vss.n1703 27.8593
R6628 vss.n3960 vss.n1703 27.8593
R6629 vss.n3961 vss.n3960 27.8593
R6630 vss.n3961 vss.n1691 27.8593
R6631 vss.n3969 vss.n1691 27.8593
R6632 vss.n3970 vss.n3969 27.8593
R6633 vss.n3970 vss.n1679 27.8593
R6634 vss.n3978 vss.n1679 27.8593
R6635 vss.n3979 vss.n3978 27.8593
R6636 vss.n3979 vss.n1674 27.8593
R6637 vss.n1674 vss.n1669 27.8593
R6638 vss.n1669 vss.n1649 27.8593
R6639 vss.n3993 vss.n1649 27.8593
R6640 vss.n3994 vss.n3993 27.8593
R6641 vss.n3994 vss.n1637 27.8593
R6642 vss.n4002 vss.n1637 27.8593
R6643 vss.n4003 vss.n4002 27.8593
R6644 vss.n4003 vss.n1625 27.8593
R6645 vss.n4011 vss.n1625 27.8593
R6646 vss.n4012 vss.n4011 27.8593
R6647 vss.n4012 vss.n1620 27.8593
R6648 vss.n1620 vss.n1615 27.8593
R6649 vss.n1615 vss.n1595 27.8593
R6650 vss.n4026 vss.n1595 27.8593
R6651 vss.n4027 vss.n4026 27.8593
R6652 vss.n4027 vss.n1583 27.8593
R6653 vss.n4035 vss.n1583 27.8593
R6654 vss.n4036 vss.n4035 27.8593
R6655 vss.n4036 vss.n1571 27.8593
R6656 vss.n4044 vss.n1571 27.8593
R6657 vss.n4045 vss.n4044 27.8593
R6658 vss.n4045 vss.n1559 27.8593
R6659 vss.n4053 vss.n1559 27.8593
R6660 vss.n4054 vss.n4053 27.8593
R6661 vss.n4054 vss.n1536 27.8593
R6662 vss.n4062 vss.n1536 27.8593
R6663 vss.n4063 vss.n4062 27.8593
R6664 vss.n4063 vss.n1524 27.8593
R6665 vss.n4071 vss.n1524 27.8593
R6666 vss.n4072 vss.n4071 27.8593
R6667 vss.n4072 vss.n1512 27.8593
R6668 vss.n4080 vss.n1512 27.8593
R6669 vss.n4081 vss.n4080 27.8593
R6670 vss.n4081 vss.n1507 27.8593
R6671 vss.n1507 vss.n1502 27.8593
R6672 vss.n1502 vss.n1482 27.8593
R6673 vss.n4095 vss.n1482 27.8593
R6674 vss.n4096 vss.n4095 27.8593
R6675 vss.n4096 vss.n1470 27.8593
R6676 vss.n4104 vss.n1470 27.8593
R6677 vss.n4105 vss.n4104 27.8593
R6678 vss.n4105 vss.n1458 27.8593
R6679 vss.n4113 vss.n1458 27.8593
R6680 vss.n4114 vss.n4113 27.8593
R6681 vss.n4114 vss.n1453 27.8593
R6682 vss.n1453 vss.n1448 27.8593
R6683 vss.n1448 vss.n1428 27.8593
R6684 vss.n4128 vss.n1428 27.8593
R6685 vss.n4129 vss.n4128 27.8593
R6686 vss.n4129 vss.n1416 27.8593
R6687 vss.n4137 vss.n1416 27.8593
R6688 vss.n4138 vss.n4137 27.8593
R6689 vss.n4138 vss.n1404 27.8593
R6690 vss.n4146 vss.n1404 27.8593
R6691 vss.n4147 vss.n4146 27.8593
R6692 vss.n4147 vss.n1392 27.8593
R6693 vss.n4155 vss.n1392 27.8593
R6694 vss.n4156 vss.n4155 27.8593
R6695 vss.n4156 vss.n1380 27.8593
R6696 vss.n4164 vss.n1380 27.8593
R6697 vss.n4165 vss.n4164 27.8593
R6698 vss.n4165 vss.n1368 27.8593
R6699 vss.n4173 vss.n1368 27.8593
R6700 vss.n4174 vss.n4173 27.8593
R6701 vss.n4174 vss.n1357 27.8593
R6702 vss.n4182 vss.n1357 27.8593
R6703 vss.n4183 vss.n4182 27.8593
R6704 vss.n4183 vss.n1345 27.8593
R6705 vss.n4191 vss.n1345 27.8593
R6706 vss.n4192 vss.n4191 27.8593
R6707 vss.n4192 vss.n1340 27.8593
R6708 vss.n1340 vss.n1331 27.8593
R6709 vss.n4202 vss.n1331 27.8593
R6710 vss.n4202 vss.n1332 27.8593
R6711 vss.n2993 vss.n1332 27.8593
R6712 vss.n2993 vss.n2349 27.8593
R6713 vss.n3004 vss.n2349 27.8593
R6714 vss.n3004 vss.n2962 27.8593
R6715 vss.n2962 vss.n2350 27.8593
R6716 vss.n2359 vss.n2350 27.8593
R6717 vss.n2361 vss.n2359 27.8593
R6718 vss.n2369 vss.n2361 27.8593
R6719 vss.n2370 vss.n2369 27.8593
R6720 vss.n2945 vss.n2370 27.8593
R6721 vss.n2945 vss.n2944 27.8593
R6722 vss.n2944 vss.n2463 27.8593
R6723 vss.n2936 vss.n2463 27.8593
R6724 vss.n2936 vss.n2935 27.8593
R6725 vss.n2935 vss.n2475 27.8593
R6726 vss.n2927 vss.n2475 27.8593
R6727 vss.n2927 vss.n2926 27.8593
R6728 vss.n2926 vss.n2488 27.8593
R6729 vss.n2504 vss.n2488 27.8593
R6730 vss.n2505 vss.n2504 27.8593
R6731 vss.n2914 vss.n2505 27.8593
R6732 vss.n2914 vss.n2913 27.8593
R6733 vss.n2913 vss.n2514 27.8593
R6734 vss.n2525 vss.n2514 27.8593
R6735 vss.n2527 vss.n2525 27.8593
R6736 vss.n2534 vss.n2527 27.8593
R6737 vss.n2897 vss.n2534 27.8593
R6738 vss.n2897 vss.n2896 27.8593
R6739 vss.n2896 vss.n2539 27.8593
R6740 vss.n2552 vss.n2539 27.8593
R6741 vss.n2554 vss.n2552 27.8593
R6742 vss.n2562 vss.n2554 27.8593
R6743 vss.n2569 vss.n2562 27.8593
R6744 vss.n2571 vss.n2569 27.8593
R6745 vss.n2577 vss.n2571 27.8593
R6746 vss.n2873 vss.n2577 27.8593
R6747 vss.n2873 vss.n2872 27.8593
R6748 vss.n2872 vss.n2585 27.8593
R6749 vss.n2864 vss.n2585 27.8593
R6750 vss.n2864 vss.n2863 27.8593
R6751 vss.n2863 vss.n2598 27.8593
R6752 vss.n2616 vss.n2598 27.8593
R6753 vss.n2617 vss.n2616 27.8593
R6754 vss.n2851 vss.n2617 27.8593
R6755 vss.n2851 vss.n2850 27.8593
R6756 vss.n2850 vss.n2625 27.8593
R6757 vss.n2842 vss.n2625 27.8593
R6758 vss.n2842 vss.n2841 27.8593
R6759 vss.n2841 vss.n2638 27.8593
R6760 vss.n2650 vss.n2638 27.8593
R6761 vss.n2652 vss.n2650 27.8593
R6762 vss.n2660 vss.n2652 27.8593
R6763 vss.n2670 vss.n2660 27.8593
R6764 vss.n2671 vss.n2670 27.8593
R6765 vss.n2675 vss.n2671 27.8593
R6766 vss.n2677 vss.n2675 27.8593
R6767 vss.n2685 vss.n2677 27.8593
R6768 vss.n2813 vss.n2685 27.8593
R6769 vss.n2813 vss.n2812 27.8593
R6770 vss.n2812 vss.n2693 27.8593
R6771 vss.n2804 vss.n2693 27.8593
R6772 vss.n2804 vss.n2803 27.8593
R6773 vss.n2803 vss.n2709 27.8593
R6774 vss.n2721 vss.n2709 27.8593
R6775 vss.n2723 vss.n2721 27.8593
R6776 vss.n2731 vss.n2723 27.8593
R6777 vss.n2788 vss.n2731 27.8593
R6778 vss.n2788 vss.n2787 27.8593
R6779 vss.n2787 vss.n2739 27.8593
R6780 vss.n2779 vss.n2739 27.8593
R6781 vss.n2779 vss.n2778 27.8593
R6782 vss.n2778 vss.n2752 27.8593
R6783 vss.n2770 vss.n2752 27.8593
R6784 vss.n2770 vss.n2769 27.8593
R6785 vss.n2769 vss.n213 27.8593
R6786 vss.n213 vss.n203 27.8593
R6787 vss.n5928 vss.n203 27.8593
R6788 vss.n5929 vss.n5928 27.8593
R6789 vss.n5929 vss.n193 27.8593
R6790 vss.n5937 vss.n193 27.8593
R6791 vss.n5938 vss.n5937 27.8593
R6792 vss.n5938 vss.n182 27.8593
R6793 vss.n5946 vss.n182 27.8593
R6794 vss.n5947 vss.n5946 27.8593
R6795 vss.n5947 vss.n177 27.8593
R6796 vss.n177 vss.n166 27.8593
R6797 vss.n5958 vss.n166 27.8593
R6798 vss.n5959 vss.n5958 27.8593
R6799 vss.n5959 vss.n161 27.8593
R6800 vss.n161 vss.n152 27.8593
R6801 vss.n6001 vss.n152 27.8593
R6802 vss.n6001 vss.n153 27.8593
R6803 vss.n5973 vss.n153 27.8593
R6804 vss.n5977 vss.n5973 27.8593
R6805 vss.n5979 vss.n5977 27.8593
R6806 vss.n5984 vss.n5979 27.8593
R6807 vss.n5984 vss.n5983 27.8593
R6808 vss.n5983 vss.n132 27.8593
R6809 vss.n2274 vss.n2268 27.8511
R6810 vss.n2294 vss.n2293 27.4829
R6811 vss.n2222 vss.n2219 27.4829
R6812 vss.n4222 vss.n1309 27.4829
R6813 vss.n2975 vss.n2972 27.4829
R6814 vss.n2405 vss.n2404 27.4829
R6815 vss.n2438 vss.n2378 27.4829
R6816 vss.n2291 vss.n2231 27.4829
R6817 vss.n2304 vss.n2303 27.4829
R6818 vss.n2317 vss.n2315 27.4829
R6819 vss.n2320 vss.n2318 27.4829
R6820 vss.n4216 vss.n4215 27.4829
R6821 vss.n4212 vss.n4211 27.4829
R6822 vss.n4211 vss.n1316 27.4829
R6823 vss.n2973 vss.n2333 27.4829
R6824 vss.n3012 vss.n2334 27.4829
R6825 vss.n2411 vss.n2410 27.4829
R6826 vss.n2444 vss.n2379 27.4829
R6827 vss.n2448 vss.n2446 27.4829
R6828 vss.n5536 vss.n300 27.4829
R6829 vss.n5536 vss.n5535 27.4829
R6830 vss.n5534 vss.n302 27.4829
R6831 vss.n2388 vss.n2385 27.1862
R6832 vss.n2510 vss.n371 27.1862
R6833 vss.n2623 vss.n2622 27.1862
R6834 vss.n2698 vss.n637 27.1862
R6835 vss.n5378 vss.n5377 27.1862
R6836 vss.n151 vss.n139 27.1522
R6837 vss.n6003 vss.n139 27.1522
R6838 vss.n148 vss.n140 27.1522
R6839 vss.n6004 vss.n140 27.1522
R6840 vss.n149 vss.n141 27.1522
R6841 vss.n6005 vss.n141 27.1522
R6842 vss.n6005 vss.n135 27.1522
R6843 vss.n6004 vss.n142 27.1522
R6844 vss.n6003 vss.n143 27.1522
R6845 vss.n149 vss.n142 27.1522
R6846 vss.n148 vss.n143 27.1522
R6847 vss.n6002 vss.n151 27.1522
R6848 vss.n5151 vss.n1114 27.1064
R6849 vss.n5159 vss.n1092 27.1064
R6850 vss.n5163 vss.n1090 27.1064
R6851 vss.n5171 vss.n1068 27.1064
R6852 vss.n5175 vss.n1066 27.1064
R6853 vss.n5183 vss.n1044 27.1064
R6854 vss.n5187 vss.n1042 27.1064
R6855 vss.n5202 vss.n1020 27.1064
R6856 vss.n5207 vss.n1018 27.1064
R6857 vss.n5525 vss.n318 27.1064
R6858 vss.n5524 vss.n5523 27.1064
R6859 vss.n5517 vss.n322 27.1064
R6860 vss.n5516 vss.n5515 27.1064
R6861 vss.n5509 vss.n350 27.1064
R6862 vss.n5508 vss.n5507 27.1064
R6863 vss.n5501 vss.n378 27.1064
R6864 vss.n5500 vss.n5499 27.1064
R6865 vss.n5493 vss.n406 27.1064
R6866 vss.n5492 vss.n5491 27.1064
R6867 vss.n5485 vss.n434 27.1064
R6868 vss.n5484 vss.n5483 27.1064
R6869 vss.n5477 vss.n462 27.1064
R6870 vss.n5476 vss.n5475 27.1064
R6871 vss.n5469 vss.n490 27.1064
R6872 vss.n5468 vss.n5467 27.1064
R6873 vss.n5461 vss.n518 27.1064
R6874 vss.n5460 vss.n5459 27.1064
R6875 vss.n5453 vss.n546 27.1064
R6876 vss.n5452 vss.n5451 27.1064
R6877 vss.n5445 vss.n574 27.1064
R6878 vss.n5444 vss.n5443 27.1064
R6879 vss.n5437 vss.n602 27.1064
R6880 vss.n5436 vss.n5435 27.1064
R6881 vss.n5429 vss.n630 27.1064
R6882 vss.n5428 vss.n5427 27.1064
R6883 vss.n5421 vss.n658 27.1064
R6884 vss.n5420 vss.n5419 27.1064
R6885 vss.n5413 vss.n686 27.1064
R6886 vss.n5412 vss.n5411 27.1064
R6887 vss.n5405 vss.n714 27.1064
R6888 vss.n5404 vss.n740 27.1064
R6889 vss.n914 vss.n762 27.1064
R6890 vss.n917 vss.n777 27.1064
R6891 vss.n920 vss.n793 27.1064
R6892 vss.n923 vss.n809 27.1064
R6893 vss.n926 vss.n828 27.1064
R6894 vss.n929 vss.n842 27.1064
R6895 vss.n932 vss.n860 27.1064
R6896 vss.n943 vss.n883 27.1064
R6897 vss.n942 vss.n941 27.1064
R6898 vss.n1259 vss.n1106 27.1064
R6899 vss.n1255 vss.n1094 27.1064
R6900 vss.n1252 vss.n1082 27.1064
R6901 vss.n1249 vss.n1070 27.1064
R6902 vss.n1246 vss.n1058 27.1064
R6903 vss.n1243 vss.n1046 27.1064
R6904 vss.n1240 vss.n1034 27.1064
R6905 vss.n1237 vss.n1022 27.1064
R6906 vss.n1234 vss.n1010 27.1064
R6907 vss.n1231 vss.n309 27.1064
R6908 vss.n1228 vss.n323 27.1064
R6909 vss.n1225 vss.n337 27.1064
R6910 vss.n1222 vss.n351 27.1064
R6911 vss.n1219 vss.n365 27.1064
R6912 vss.n1216 vss.n379 27.1064
R6913 vss.n1213 vss.n393 27.1064
R6914 vss.n1210 vss.n407 27.1064
R6915 vss.n1207 vss.n421 27.1064
R6916 vss.n1204 vss.n435 27.1064
R6917 vss.n1201 vss.n449 27.1064
R6918 vss.n1198 vss.n463 27.1064
R6919 vss.n1195 vss.n477 27.1064
R6920 vss.n1192 vss.n491 27.1064
R6921 vss.n1189 vss.n505 27.1064
R6922 vss.n1186 vss.n519 27.1064
R6923 vss.n1183 vss.n533 27.1064
R6924 vss.n1180 vss.n547 27.1064
R6925 vss.n1177 vss.n561 27.1064
R6926 vss.n1174 vss.n575 27.1064
R6927 vss.n1171 vss.n589 27.1064
R6928 vss.n1168 vss.n603 27.1064
R6929 vss.n1165 vss.n617 27.1064
R6930 vss.n1162 vss.n631 27.1064
R6931 vss.n1159 vss.n645 27.1064
R6932 vss.n1156 vss.n659 27.1064
R6933 vss.n1153 vss.n673 27.1064
R6934 vss.n1150 vss.n687 27.1064
R6935 vss.n1147 vss.n701 27.1064
R6936 vss.n1144 vss.n715 27.1064
R6937 vss.n1141 vss.n729 27.1064
R6938 vss.n747 vss.n741 27.1064
R6939 vss.n1136 vss.n771 27.1064
R6940 vss.n1133 vss.n787 27.1064
R6941 vss.n1130 vss.n805 27.1064
R6942 vss.n1127 vss.n820 27.1064
R6943 vss.n1124 vss.n840 27.1064
R6944 vss.n1121 vss.n852 27.1064
R6945 vss.n1118 vss.n876 27.1064
R6946 vss.n5356 vss.n5355 27.1064
R6947 vss.n910 vss.n909 27.1064
R6948 vss.n5153 vss.n1104 27.1064
R6949 vss.n5157 vss.n1102 27.1064
R6950 vss.n5165 vss.n1080 27.1064
R6951 vss.n5169 vss.n1078 27.1064
R6952 vss.n5177 vss.n1056 27.1064
R6953 vss.n5181 vss.n1054 27.1064
R6954 vss.n5189 vss.n1032 27.1064
R6955 vss.n5200 vss.n1030 27.1064
R6956 vss.n5199 vss.n1017 27.1064
R6957 vss.n5195 vss.n317 27.1064
R6958 vss.n5521 vss.n332 27.1064
R6959 vss.n5520 vss.n5519 27.1064
R6960 vss.n5513 vss.n336 27.1064
R6961 vss.n5512 vss.n5511 27.1064
R6962 vss.n5505 vss.n364 27.1064
R6963 vss.n5504 vss.n5503 27.1064
R6964 vss.n5497 vss.n392 27.1064
R6965 vss.n5496 vss.n5495 27.1064
R6966 vss.n5489 vss.n420 27.1064
R6967 vss.n5488 vss.n5487 27.1064
R6968 vss.n5481 vss.n448 27.1064
R6969 vss.n5480 vss.n5479 27.1064
R6970 vss.n5473 vss.n476 27.1064
R6971 vss.n5472 vss.n5471 27.1064
R6972 vss.n5465 vss.n504 27.1064
R6973 vss.n5464 vss.n5463 27.1064
R6974 vss.n5457 vss.n532 27.1064
R6975 vss.n5456 vss.n5455 27.1064
R6976 vss.n5449 vss.n560 27.1064
R6977 vss.n5448 vss.n5447 27.1064
R6978 vss.n5441 vss.n588 27.1064
R6979 vss.n5440 vss.n5439 27.1064
R6980 vss.n5433 vss.n616 27.1064
R6981 vss.n5432 vss.n5431 27.1064
R6982 vss.n5425 vss.n644 27.1064
R6983 vss.n5424 vss.n5423 27.1064
R6984 vss.n5417 vss.n672 27.1064
R6985 vss.n5416 vss.n5415 27.1064
R6986 vss.n5409 vss.n700 27.1064
R6987 vss.n5408 vss.n5407 27.1064
R6988 vss.n5393 vss.n728 27.1064
R6989 vss.n5392 vss.n5391 27.1064
R6990 vss.n778 vss.n761 27.1064
R6991 vss.n946 vss.n794 27.1064
R6992 vss.n949 vss.n810 27.1064
R6993 vss.n952 vss.n829 27.1064
R6994 vss.n955 vss.n843 27.1064
R6995 vss.n958 vss.n861 27.1064
R6996 vss.n969 vss.n884 27.1064
R6997 vss.n968 vss.n967 27.1064
R6998 vss.n1286 vss.n1107 27.1064
R6999 vss.n1282 vss.n1095 27.1064
R7000 vss.n1279 vss.n1083 27.1064
R7001 vss.n1276 vss.n1071 27.1064
R7002 vss.n1273 vss.n1059 27.1064
R7003 vss.n1270 vss.n1047 27.1064
R7004 vss.n1267 vss.n1035 27.1064
R7005 vss.n1264 vss.n1023 27.1064
R7006 vss.n5209 vss.n1008 27.1064
R7007 vss.n5210 vss.n310 27.1064
R7008 vss.n5213 vss.n324 27.1064
R7009 vss.n5216 vss.n338 27.1064
R7010 vss.n5219 vss.n352 27.1064
R7011 vss.n5222 vss.n366 27.1064
R7012 vss.n5225 vss.n380 27.1064
R7013 vss.n5228 vss.n394 27.1064
R7014 vss.n5231 vss.n408 27.1064
R7015 vss.n5234 vss.n422 27.1064
R7016 vss.n5237 vss.n436 27.1064
R7017 vss.n5240 vss.n450 27.1064
R7018 vss.n5243 vss.n464 27.1064
R7019 vss.n5246 vss.n478 27.1064
R7020 vss.n5249 vss.n492 27.1064
R7021 vss.n5252 vss.n506 27.1064
R7022 vss.n5255 vss.n520 27.1064
R7023 vss.n5258 vss.n534 27.1064
R7024 vss.n5261 vss.n548 27.1064
R7025 vss.n5264 vss.n562 27.1064
R7026 vss.n5267 vss.n576 27.1064
R7027 vss.n5270 vss.n590 27.1064
R7028 vss.n5273 vss.n604 27.1064
R7029 vss.n5276 vss.n618 27.1064
R7030 vss.n5279 vss.n632 27.1064
R7031 vss.n5282 vss.n646 27.1064
R7032 vss.n5285 vss.n660 27.1064
R7033 vss.n5288 vss.n674 27.1064
R7034 vss.n5291 vss.n688 27.1064
R7035 vss.n5294 vss.n702 27.1064
R7036 vss.n5297 vss.n716 27.1064
R7037 vss.n5300 vss.n730 27.1064
R7038 vss.n748 vss.n742 27.1064
R7039 vss.n5305 vss.n770 27.1064
R7040 vss.n5308 vss.n786 27.1064
R7041 vss.n5311 vss.n804 27.1064
R7042 vss.n5314 vss.n819 27.1064
R7043 vss.n5317 vss.n839 27.1064
R7044 vss.n5320 vss.n851 27.1064
R7045 vss.n5323 vss.n874 27.1064
R7046 vss.n5334 vss.n901 27.1064
R7047 vss.n5333 vss.n5332 27.1064
R7048 vss.n5142 vss.n1113 27.1064
R7049 vss.n5138 vss.n1101 27.1064
R7050 vss.n5135 vss.n1089 27.1064
R7051 vss.n5132 vss.n1077 27.1064
R7052 vss.n5129 vss.n1065 27.1064
R7053 vss.n5126 vss.n1053 27.1064
R7054 vss.n5123 vss.n1041 27.1064
R7055 vss.n5120 vss.n1029 27.1064
R7056 vss.n5117 vss.n1016 27.1064
R7057 vss.n5114 vss.n316 27.1064
R7058 vss.n5111 vss.n331 27.1064
R7059 vss.n5108 vss.n345 27.1064
R7060 vss.n5105 vss.n359 27.1064
R7061 vss.n5102 vss.n373 27.1064
R7062 vss.n5099 vss.n387 27.1064
R7063 vss.n5096 vss.n401 27.1064
R7064 vss.n5093 vss.n415 27.1064
R7065 vss.n5090 vss.n429 27.1064
R7066 vss.n5087 vss.n443 27.1064
R7067 vss.n5084 vss.n457 27.1064
R7068 vss.n5081 vss.n471 27.1064
R7069 vss.n5078 vss.n485 27.1064
R7070 vss.n5075 vss.n499 27.1064
R7071 vss.n5072 vss.n513 27.1064
R7072 vss.n5069 vss.n527 27.1064
R7073 vss.n5066 vss.n541 27.1064
R7074 vss.n5063 vss.n555 27.1064
R7075 vss.n5060 vss.n569 27.1064
R7076 vss.n5057 vss.n583 27.1064
R7077 vss.n5054 vss.n597 27.1064
R7078 vss.n5051 vss.n611 27.1064
R7079 vss.n5048 vss.n625 27.1064
R7080 vss.n5045 vss.n639 27.1064
R7081 vss.n5042 vss.n653 27.1064
R7082 vss.n5039 vss.n667 27.1064
R7083 vss.n5036 vss.n681 27.1064
R7084 vss.n5033 vss.n695 27.1064
R7085 vss.n5030 vss.n709 27.1064
R7086 vss.n5027 vss.n723 27.1064
R7087 vss.n5024 vss.n736 27.1064
R7088 vss.n5396 vss.n5395 27.1064
R7089 vss.n763 vss.n745 27.1064
R7090 vss.n973 vss.n779 27.1064
R7091 vss.n976 vss.n795 27.1064
R7092 vss.n979 vss.n811 27.1064
R7093 vss.n982 vss.n830 27.1064
R7094 vss.n985 vss.n844 27.1064
R7095 vss.n988 vss.n862 27.1064
R7096 vss.n999 vss.n886 27.1064
R7097 vss.n998 vss.n997 27.1064
R7098 vss.n4744 vss.n1108 27.1064
R7099 vss.n4747 vss.n1096 27.1064
R7100 vss.n4750 vss.n1084 27.1064
R7101 vss.n4753 vss.n1072 27.1064
R7102 vss.n4756 vss.n1060 27.1064
R7103 vss.n4759 vss.n1048 27.1064
R7104 vss.n4762 vss.n1036 27.1064
R7105 vss.n4765 vss.n1024 27.1064
R7106 vss.n4768 vss.n1011 27.1064
R7107 vss.n4771 vss.n311 27.1064
R7108 vss.n4774 vss.n325 27.1064
R7109 vss.n4777 vss.n339 27.1064
R7110 vss.n4780 vss.n353 27.1064
R7111 vss.n4783 vss.n367 27.1064
R7112 vss.n4786 vss.n381 27.1064
R7113 vss.n4789 vss.n395 27.1064
R7114 vss.n4792 vss.n409 27.1064
R7115 vss.n4795 vss.n423 27.1064
R7116 vss.n4798 vss.n437 27.1064
R7117 vss.n4801 vss.n451 27.1064
R7118 vss.n4804 vss.n465 27.1064
R7119 vss.n4807 vss.n479 27.1064
R7120 vss.n4810 vss.n493 27.1064
R7121 vss.n4813 vss.n507 27.1064
R7122 vss.n4816 vss.n521 27.1064
R7123 vss.n4819 vss.n535 27.1064
R7124 vss.n4822 vss.n549 27.1064
R7125 vss.n4825 vss.n563 27.1064
R7126 vss.n4828 vss.n577 27.1064
R7127 vss.n4831 vss.n591 27.1064
R7128 vss.n4834 vss.n605 27.1064
R7129 vss.n4837 vss.n619 27.1064
R7130 vss.n4840 vss.n633 27.1064
R7131 vss.n4843 vss.n647 27.1064
R7132 vss.n4846 vss.n661 27.1064
R7133 vss.n4849 vss.n675 27.1064
R7134 vss.n4852 vss.n689 27.1064
R7135 vss.n4855 vss.n703 27.1064
R7136 vss.n4858 vss.n717 27.1064
R7137 vss.n4861 vss.n731 27.1064
R7138 vss.n4895 vss.n749 27.1064
R7139 vss.n4891 vss.n769 27.1064
R7140 vss.n4888 vss.n785 27.1064
R7141 vss.n4885 vss.n803 27.1064
R7142 vss.n4882 vss.n818 27.1064
R7143 vss.n4879 vss.n838 27.1064
R7144 vss.n4876 vss.n850 27.1064
R7145 vss.n4873 vss.n872 27.1064
R7146 vss.n1006 vss.n899 27.1064
R7147 vss.n4868 vss.n4867 27.1064
R7148 vss.n5020 vss.n1112 27.1064
R7149 vss.n5016 vss.n1100 27.1064
R7150 vss.n5013 vss.n1088 27.1064
R7151 vss.n5010 vss.n1076 27.1064
R7152 vss.n5007 vss.n1064 27.1064
R7153 vss.n5004 vss.n1052 27.1064
R7154 vss.n5001 vss.n1040 27.1064
R7155 vss.n4998 vss.n1028 27.1064
R7156 vss.n4995 vss.n1015 27.1064
R7157 vss.n4992 vss.n315 27.1064
R7158 vss.n4989 vss.n330 27.1064
R7159 vss.n4986 vss.n344 27.1064
R7160 vss.n4983 vss.n358 27.1064
R7161 vss.n4980 vss.n372 27.1064
R7162 vss.n4977 vss.n386 27.1064
R7163 vss.n4974 vss.n400 27.1064
R7164 vss.n4971 vss.n414 27.1064
R7165 vss.n4968 vss.n428 27.1064
R7166 vss.n4965 vss.n442 27.1064
R7167 vss.n4962 vss.n456 27.1064
R7168 vss.n4959 vss.n470 27.1064
R7169 vss.n4956 vss.n484 27.1064
R7170 vss.n4953 vss.n498 27.1064
R7171 vss.n4950 vss.n512 27.1064
R7172 vss.n4947 vss.n526 27.1064
R7173 vss.n4944 vss.n540 27.1064
R7174 vss.n4941 vss.n554 27.1064
R7175 vss.n4938 vss.n568 27.1064
R7176 vss.n4935 vss.n582 27.1064
R7177 vss.n4932 vss.n596 27.1064
R7178 vss.n4929 vss.n610 27.1064
R7179 vss.n4926 vss.n624 27.1064
R7180 vss.n4923 vss.n638 27.1064
R7181 vss.n4920 vss.n652 27.1064
R7182 vss.n4917 vss.n666 27.1064
R7183 vss.n4914 vss.n680 27.1064
R7184 vss.n4911 vss.n694 27.1064
R7185 vss.n4908 vss.n708 27.1064
R7186 vss.n4905 vss.n722 27.1064
R7187 vss.n4902 vss.n735 27.1064
R7188 vss.n4899 vss.n756 27.1064
R7189 vss.n4263 vss.n764 27.1064
R7190 vss.n4260 vss.n780 27.1064
R7191 vss.n4257 vss.n796 27.1064
R7192 vss.n4254 vss.n812 27.1064
R7193 vss.n4251 vss.n831 27.1064
R7194 vss.n4248 vss.n845 27.1064
R7195 vss.n4245 vss.n863 27.1064
R7196 vss.n1001 vss.n888 27.1064
R7197 vss.n4240 vss.n4239 27.1064
R7198 vss.n4590 vss.n1109 27.1064
R7199 vss.n4593 vss.n1097 27.1064
R7200 vss.n4596 vss.n1085 27.1064
R7201 vss.n4599 vss.n1073 27.1064
R7202 vss.n4602 vss.n1061 27.1064
R7203 vss.n4605 vss.n1049 27.1064
R7204 vss.n4608 vss.n1037 27.1064
R7205 vss.n4611 vss.n1025 27.1064
R7206 vss.n4614 vss.n1012 27.1064
R7207 vss.n4617 vss.n312 27.1064
R7208 vss.n4620 vss.n326 27.1064
R7209 vss.n4623 vss.n340 27.1064
R7210 vss.n4626 vss.n354 27.1064
R7211 vss.n4629 vss.n368 27.1064
R7212 vss.n4632 vss.n382 27.1064
R7213 vss.n4635 vss.n396 27.1064
R7214 vss.n4638 vss.n410 27.1064
R7215 vss.n4641 vss.n424 27.1064
R7216 vss.n4644 vss.n438 27.1064
R7217 vss.n4647 vss.n452 27.1064
R7218 vss.n4650 vss.n466 27.1064
R7219 vss.n4653 vss.n480 27.1064
R7220 vss.n4656 vss.n494 27.1064
R7221 vss.n4659 vss.n508 27.1064
R7222 vss.n4662 vss.n522 27.1064
R7223 vss.n4665 vss.n536 27.1064
R7224 vss.n4668 vss.n550 27.1064
R7225 vss.n4671 vss.n564 27.1064
R7226 vss.n4674 vss.n578 27.1064
R7227 vss.n4677 vss.n592 27.1064
R7228 vss.n4680 vss.n606 27.1064
R7229 vss.n4683 vss.n620 27.1064
R7230 vss.n4686 vss.n634 27.1064
R7231 vss.n4689 vss.n648 27.1064
R7232 vss.n4692 vss.n662 27.1064
R7233 vss.n4695 vss.n676 27.1064
R7234 vss.n4698 vss.n690 27.1064
R7235 vss.n4701 vss.n704 27.1064
R7236 vss.n4704 vss.n718 27.1064
R7237 vss.n4707 vss.n732 27.1064
R7238 vss.n4741 vss.n750 27.1064
R7239 vss.n4737 vss.n768 27.1064
R7240 vss.n4734 vss.n784 27.1064
R7241 vss.n4731 vss.n802 27.1064
R7242 vss.n4728 vss.n817 27.1064
R7243 vss.n4725 vss.n837 27.1064
R7244 vss.n4722 vss.n849 27.1064
R7245 vss.n4719 vss.n870 27.1064
R7246 vss.n1005 vss.n897 27.1064
R7247 vss.n4714 vss.n4713 27.1064
R7248 vss.n4576 vss.n772 27.1064
R7249 vss.n5383 vss.n788 27.1064
R7250 vss.n5382 vss.n5381 27.1064
R7251 vss.n5373 vss.n792 27.1064
R7252 vss.n5372 vss.n5371 27.1064
R7253 vss.n5363 vss.n827 27.1064
R7254 vss.n5362 vss.n5361 27.1064
R7255 vss.n5353 vss.n859 27.1064
R7256 vss.n5352 vss.n5351 27.1064
R7257 vss.n5350 vss.n5349 27.1064
R7258 vss.n4586 vss.n753 27.1064
R7259 vss.n4581 vss.n767 27.1064
R7260 vss.n4577 vss.n783 27.1064
R7261 vss.n801 vss.n800 27.1064
R7262 vss.n821 vss.n816 27.1064
R7263 vss.n836 vss.n835 27.1064
R7264 vss.n853 vss.n848 27.1064
R7265 vss.n868 vss.n867 27.1064
R7266 vss.n1004 vss.n894 27.1064
R7267 vss.n5341 vss.n5340 27.1064
R7268 vss.n5343 vss.n5342 27.1064
R7269 vss.n2288 vss.n2245 27.1064
R7270 vss.n2307 vss.n2229 27.1064
R7271 vss.n4231 vss.n1297 27.1064
R7272 vss.n4230 vss.n4229 27.1064
R7273 vss.n3022 vss.n1301 27.1064
R7274 vss.n4208 vss.n1319 27.1064
R7275 vss.n2987 vss.n1320 27.1064
R7276 vss.n3009 vss.n2338 27.1064
R7277 vss.n2390 vss.n2339 27.1064
R7278 vss.n2428 vss.n2427 27.1064
R7279 vss.n2451 vss.n2374 27.1064
R7280 vss.n2248 vss.n2241 27.1064
R7281 vss.n2242 vss.n2209 27.1064
R7282 vss.n2312 vss.n2214 27.1064
R7283 vss.n2213 vss.n2210 27.1064
R7284 vss.n2197 vss.n1311 27.1064
R7285 vss.n2198 vss.n1317 27.1064
R7286 vss.n2984 vss.n2981 27.1064
R7287 vss.n2983 vss.n2336 27.1064
R7288 vss.n2423 vss.n2392 27.1064
R7289 vss.n2424 vss.n2387 27.1064
R7290 vss.n2381 vss.n2376 27.1064
R7291 vss.n5543 vss.n296 27.1064
R7292 vss.n5575 vss.n5574 27.1064
R7293 vss.n5583 vss.n5582 27.1064
R7294 vss.n5583 vss.n261 27.1064
R7295 vss.n5592 vss.n261 27.1064
R7296 vss.n5593 vss.n5592 27.1064
R7297 vss.n5594 vss.n5593 27.1064
R7298 vss.n5594 vss.n255 27.1064
R7299 vss.n5602 vss.n255 27.1064
R7300 vss.n5603 vss.n5602 27.1064
R7301 vss.n5603 vss.n249 27.1064
R7302 vss.n5611 vss.n249 27.1064
R7303 vss.n5613 vss.n5611 27.1064
R7304 vss.n5613 vss.n5612 27.1064
R7305 vss.n5612 vss.n231 27.1064
R7306 vss.n5909 vss.n231 27.1064
R7307 vss.n5909 vss.n5908 27.1064
R7308 vss.n5908 vss.n5907 27.1064
R7309 vss.n5907 vss.n232 27.1064
R7310 vss.n5631 vss.n232 27.1064
R7311 vss.n5897 vss.n5631 27.1064
R7312 vss.n5897 vss.n5896 27.1064
R7313 vss.n5896 vss.n5632 27.1064
R7314 vss.n5646 vss.n5632 27.1064
R7315 vss.n5885 vss.n5646 27.1064
R7316 vss.n5885 vss.n5884 27.1064
R7317 vss.n5884 vss.n5647 27.1064
R7318 vss.n5878 vss.n5647 27.1064
R7319 vss.n5878 vss.n5877 27.1064
R7320 vss.n5877 vss.n5655 27.1064
R7321 vss.n5870 vss.n5655 27.1064
R7322 vss.n5870 vss.n5869 27.1064
R7323 vss.n5869 vss.n5668 27.1064
R7324 vss.n5682 vss.n5668 27.1064
R7325 vss.n5859 vss.n5682 27.1064
R7326 vss.n5859 vss.n5858 27.1064
R7327 vss.n5858 vss.n5683 27.1064
R7328 vss.n5852 vss.n5683 27.1064
R7329 vss.n5852 vss.n5851 27.1064
R7330 vss.n5851 vss.n5691 27.1064
R7331 vss.n5844 vss.n5691 27.1064
R7332 vss.n5844 vss.n5843 27.1064
R7333 vss.n5843 vss.n5705 27.1064
R7334 vss.n5721 vss.n5705 27.1064
R7335 vss.n5833 vss.n5721 27.1064
R7336 vss.n5833 vss.n5832 27.1064
R7337 vss.n5832 vss.n5722 27.1064
R7338 vss.n5826 vss.n5722 27.1064
R7339 vss.n5826 vss.n5825 27.1064
R7340 vss.n5825 vss.n5730 27.1064
R7341 vss.n5818 vss.n5730 27.1064
R7342 vss.n5818 vss.n5817 27.1064
R7343 vss.n5817 vss.n5744 27.1064
R7344 vss.n5758 vss.n5744 27.1064
R7345 vss.n5807 vss.n5758 27.1064
R7346 vss.n5807 vss.n5806 27.1064
R7347 vss.n5572 vss.n274 27.1064
R7348 vss.n5585 vss.n267 27.1064
R7349 vss.n5586 vss.n5585 27.1064
R7350 vss.n5586 vss.n263 27.1064
R7351 vss.n263 vss.n259 27.1064
R7352 vss.n5596 vss.n259 27.1064
R7353 vss.n5597 vss.n5596 27.1064
R7354 vss.n5597 vss.n253 27.1064
R7355 vss.n5605 vss.n253 27.1064
R7356 vss.n5606 vss.n5605 27.1064
R7357 vss.n5606 vss.n244 27.1064
R7358 vss.n5615 vss.n244 27.1064
R7359 vss.n5616 vss.n5615 27.1064
R7360 vss.n5617 vss.n5616 27.1064
R7361 vss.n5617 vss.n229 27.1064
R7362 vss.n234 vss.n229 27.1064
R7363 vss.n235 vss.n234 27.1064
R7364 vss.n238 vss.n235 27.1064
R7365 vss.n5627 vss.n238 27.1064
R7366 vss.n5628 vss.n5627 27.1064
R7367 vss.n5633 vss.n5628 27.1064
R7368 vss.n5636 vss.n5633 27.1064
R7369 vss.n5642 vss.n5636 27.1064
R7370 vss.n5643 vss.n5642 27.1064
R7371 vss.n5648 vss.n5643 27.1064
R7372 vss.n5652 vss.n5648 27.1064
R7373 vss.n5653 vss.n5652 27.1064
R7374 vss.n5656 vss.n5653 27.1064
R7375 vss.n5662 vss.n5656 27.1064
R7376 vss.n5663 vss.n5662 27.1064
R7377 vss.n5669 vss.n5663 27.1064
R7378 vss.n5672 vss.n5669 27.1064
R7379 vss.n5678 vss.n5672 27.1064
R7380 vss.n5679 vss.n5678 27.1064
R7381 vss.n5684 vss.n5679 27.1064
R7382 vss.n5688 vss.n5684 27.1064
R7383 vss.n5689 vss.n5688 27.1064
R7384 vss.n5692 vss.n5689 27.1064
R7385 vss.n5700 vss.n5692 27.1064
R7386 vss.n5701 vss.n5700 27.1064
R7387 vss.n5706 vss.n5701 27.1064
R7388 vss.n5709 vss.n5706 27.1064
R7389 vss.n5716 vss.n5709 27.1064
R7390 vss.n5717 vss.n5716 27.1064
R7391 vss.n5723 vss.n5717 27.1064
R7392 vss.n5727 vss.n5723 27.1064
R7393 vss.n5728 vss.n5727 27.1064
R7394 vss.n5731 vss.n5728 27.1064
R7395 vss.n5739 vss.n5731 27.1064
R7396 vss.n5740 vss.n5739 27.1064
R7397 vss.n5745 vss.n5740 27.1064
R7398 vss.n5748 vss.n5745 27.1064
R7399 vss.n5754 vss.n5748 27.1064
R7400 vss.n5755 vss.n5754 27.1064
R7401 vss.n5577 vss.n272 27.1064
R7402 vss.n5540 vss.n5539 27.1064
R7403 vss.n2974 vss.n2973 27.1064
R7404 vss.n4330 vss.n1110 27.1064
R7405 vss.n4333 vss.n1098 27.1064
R7406 vss.n4336 vss.n1086 27.1064
R7407 vss.n4339 vss.n1074 27.1064
R7408 vss.n4342 vss.n1062 27.1064
R7409 vss.n4345 vss.n1050 27.1064
R7410 vss.n4348 vss.n1038 27.1064
R7411 vss.n4327 vss.n1026 27.1064
R7412 vss.n4356 vss.n1013 27.1064
R7413 vss.n4387 vss.n314 27.1064
R7414 vss.n4319 vss.n328 27.1064
R7415 vss.n4316 vss.n342 27.1064
R7416 vss.n4403 vss.n356 27.1064
R7417 vss.n4410 vss.n370 27.1064
R7418 vss.n4416 vss.n384 27.1064
R7419 vss.n4308 vss.n398 27.1064
R7420 vss.n4304 vss.n412 27.1064
R7421 vss.n4433 vss.n426 27.1064
R7422 vss.n4441 vss.n440 27.1064
R7423 vss.n4299 vss.n454 27.1064
R7424 vss.n4453 vss.n468 27.1064
R7425 vss.n4461 vss.n482 27.1064
R7426 vss.n4294 vss.n496 27.1064
R7427 vss.n4473 vss.n510 27.1064
R7428 vss.n4481 vss.n524 27.1064
R7429 vss.n4486 vss.n538 27.1064
R7430 vss.n4493 vss.n552 27.1064
R7431 vss.n4497 vss.n566 27.1064
R7432 vss.n4503 vss.n580 27.1064
R7433 vss.n4284 vss.n594 27.1064
R7434 vss.n4515 vss.n608 27.1064
R7435 vss.n4523 vss.n622 27.1064
R7436 vss.n4279 vss.n636 27.1064
R7437 vss.n4535 vss.n650 27.1064
R7438 vss.n4543 vss.n664 27.1064
R7439 vss.n4274 vss.n678 27.1064
R7440 vss.n4555 vss.n692 27.1064
R7441 vss.n4563 vss.n706 27.1064
R7442 vss.n4269 vss.n720 27.1064
R7443 vss.n4571 vss.n734 27.1064
R7444 vss.n4266 vss.n755 27.1064
R7445 vss.n4582 vss.n765 27.1064
R7446 vss.n4578 vss.n781 27.1064
R7447 vss.n798 vss.n797 27.1064
R7448 vss.n822 vss.n813 27.1064
R7449 vss.n833 vss.n832 27.1064
R7450 vss.n854 vss.n846 27.1064
R7451 vss.n865 vss.n864 27.1064
R7452 vss.n1003 vss.n892 27.1064
R7453 vss.n5345 vss.n5344 27.1064
R7454 vss.n5347 vss.n5346 27.1064
R7455 vss.n2309 vss.n2216 27.0554
R7456 vss.n2292 vss.n2291 26.7299
R7457 vss.n5580 vss.n265 26.3319
R7458 vss.n5588 vss.n265 26.3319
R7459 vss.n5590 vss.n5588 26.3319
R7460 vss.n5590 vss.n5589 26.3319
R7461 vss.n5589 vss.n257 26.3319
R7462 vss.n5599 vss.n257 26.3319
R7463 vss.n5600 vss.n5599 26.3319
R7464 vss.n5600 vss.n251 26.3319
R7465 vss.n5608 vss.n251 26.3319
R7466 vss.n5609 vss.n5608 26.3319
R7467 vss.n5609 vss.n248 26.3319
R7468 vss.n248 vss.n247 26.3319
R7469 vss.n247 vss.n226 26.3319
R7470 vss.n5911 vss.n227 26.3319
R7471 vss.n5905 vss.n227 26.3319
R7472 vss.n5905 vss.n5904 26.3319
R7473 vss.n5904 vss.n237 26.3319
R7474 vss.n5630 vss.n237 26.3319
R7475 vss.n5894 vss.n5630 26.3319
R7476 vss.n5894 vss.n5893 26.3319
R7477 vss.n5893 vss.n5635 26.3319
R7478 vss.n5645 vss.n5635 26.3319
R7479 vss.n5882 vss.n5645 26.3319
R7480 vss.n5882 vss.n5881 26.3319
R7481 vss.n5881 vss.n5880 26.3319
R7482 vss.n5880 vss.n5650 26.3319
R7483 vss.n5667 vss.n5666 26.3319
R7484 vss.n5867 vss.n5667 26.3319
R7485 vss.n5867 vss.n5866 26.3319
R7486 vss.n5866 vss.n5671 26.3319
R7487 vss.n5681 vss.n5671 26.3319
R7488 vss.n5856 vss.n5681 26.3319
R7489 vss.n5856 vss.n5855 26.3319
R7490 vss.n5855 vss.n5854 26.3319
R7491 vss.n5854 vss.n5686 26.3319
R7492 vss.n5703 vss.n5686 26.3319
R7493 vss.n5704 vss.n5703 26.3319
R7494 vss.n5841 vss.n5704 26.3319
R7495 vss.n5841 vss.n5840 26.3319
R7496 vss.n5720 vss.n5719 26.3319
R7497 vss.n5830 vss.n5720 26.3319
R7498 vss.n5830 vss.n5829 26.3319
R7499 vss.n5829 vss.n5828 26.3319
R7500 vss.n5828 vss.n5725 26.3319
R7501 vss.n5742 vss.n5725 26.3319
R7502 vss.n5743 vss.n5742 26.3319
R7503 vss.n5815 vss.n5743 26.3319
R7504 vss.n5815 vss.n5814 26.3319
R7505 vss.n5814 vss.n5747 26.3319
R7506 vss.n5757 vss.n5747 26.3319
R7507 vss.n5804 vss.n5757 26.3319
R7508 vss.n5804 vss.n218 26.3319
R7509 vss.n4287 vss.n4286 26.038
R7510 vss.n4307 vss.n4306 26.038
R7511 vss.n4428 vss.n4427 26.038
R7512 vss.n4438 vss.n4437 26.038
R7513 vss.n4448 vss.n4447 26.038
R7514 vss.n4458 vss.n4457 26.038
R7515 vss.n4468 vss.n4467 26.038
R7516 vss.n4478 vss.n4477 26.038
R7517 vss.n4510 vss.n4509 26.038
R7518 vss.n4520 vss.n4519 26.038
R7519 vss.n4530 vss.n4529 26.038
R7520 vss.n4540 vss.n4539 26.038
R7521 vss.n4550 vss.n4549 26.038
R7522 vss.n4560 vss.n4559 26.038
R7523 vss.n5675 vss.n5674 25.8481
R7524 vss.n5751 vss.n5750 25.8481
R7525 vss.n5737 vss.n5733 25.8481
R7526 vss.n5715 vss.n5714 25.8481
R7527 vss.n5712 vss.n5711 25.8481
R7528 vss.n5698 vss.n5694 25.8481
R7529 vss.n5677 vss.n5676 25.8481
R7530 vss.n5889 vss.n5640 25.8481
R7531 vss.n5626 vss.n5625 25.8481
R7532 vss.n5623 vss.n240 25.8481
R7533 vss.n242 vss.n241 25.8481
R7534 vss.n5554 vss.n5550 25.8481
R7535 vss.n5558 vss.n5549 25.8481
R7536 vss.n5561 vss.n5548 25.8481
R7537 vss.t17 vss.n665 25.8269
R7538 vss.t2 vss.n2736 25.8269
R7539 vss.n2640 vss.n219 25.4353
R7540 vss.n2641 vss.n2640 25.4353
R7541 vss.n5919 vss.n5918 25.4353
R7542 vss.n5920 vss.n5919 25.4353
R7543 vss.n221 vss.n220 25.4353
R7544 vss.n2510 vss.n221 25.4353
R7545 vss.n2286 vss.n2247 24.6682
R7546 vss.n2434 vss.n1027 24.4676
R7547 vss.n2499 vss.n2498 24.4676
R7548 vss.n2564 vss.n2563 24.4676
R7549 vss.n2763 vss.n721 24.4676
R7550 vss.n5376 vss.n5375 24.4676
R7551 vss.n5579 vss.n5578 23.7047
R7552 vss.n4215 vss.n1314 23.3417
R7553 vss.n2435 vss.n2434 23.1083
R7554 vss.t25 vss.n679 23.1083
R7555 vss.n2746 vss.t296 23.1083
R7556 vss.n5146 vss.n1105 23.0776
R7557 vss.n5152 vss.n1093 23.0776
R7558 vss.n5158 vss.n1081 23.0776
R7559 vss.n5164 vss.n1069 23.0776
R7560 vss.n5170 vss.n1057 23.0776
R7561 vss.n5176 vss.n1045 23.0776
R7562 vss.n5182 vss.n1033 23.0776
R7563 vss.n5188 vss.n1021 23.0776
R7564 vss.n5201 vss.n1009 23.0776
R7565 vss.n5208 vss.n308 23.0776
R7566 vss.n5526 vss.n313 23.0776
R7567 vss.n5522 vss.n327 23.0776
R7568 vss.n5518 vss.n341 23.0776
R7569 vss.n5514 vss.n355 23.0776
R7570 vss.n5510 vss.n369 23.0776
R7571 vss.n5506 vss.n383 23.0776
R7572 vss.n5502 vss.n397 23.0776
R7573 vss.n5498 vss.n411 23.0776
R7574 vss.n5494 vss.n425 23.0776
R7575 vss.n5490 vss.n439 23.0776
R7576 vss.n5486 vss.n453 23.0776
R7577 vss.n5482 vss.n467 23.0776
R7578 vss.n5478 vss.n481 23.0776
R7579 vss.n5474 vss.n495 23.0776
R7580 vss.n5470 vss.n509 23.0776
R7581 vss.n5466 vss.n523 23.0776
R7582 vss.n5462 vss.n537 23.0776
R7583 vss.n5458 vss.n551 23.0776
R7584 vss.n5454 vss.n565 23.0776
R7585 vss.n5450 vss.n579 23.0776
R7586 vss.n5446 vss.n593 23.0776
R7587 vss.n5442 vss.n607 23.0776
R7588 vss.n5438 vss.n621 23.0776
R7589 vss.n5434 vss.n635 23.0776
R7590 vss.n5430 vss.n649 23.0776
R7591 vss.n5426 vss.n663 23.0776
R7592 vss.n5422 vss.n677 23.0776
R7593 vss.n5418 vss.n691 23.0776
R7594 vss.n5414 vss.n705 23.0776
R7595 vss.n5410 vss.n719 23.0776
R7596 vss.n2448 vss.n2447 22.9652
R7597 vss.n2294 vss.n2236 22.5887
R7598 vss.n2223 vss.n2222 22.5887
R7599 vss.n4223 vss.n4222 22.5887
R7600 vss.n2972 vss.n2971 22.5887
R7601 vss.n2404 vss.n2403 22.5887
R7602 vss.n2438 vss.n2437 22.5887
R7603 vss.n3013 vss.n3012 22.5887
R7604 vss.n5530 vss.n302 22.5887
R7605 vss.n746 vss.n733 22.3024
R7606 vss.n2303 vss.n2302 22.2123
R7607 vss.n2565 vss.n455 21.749
R7608 vss.n2641 vss.n553 21.749
R7609 vss.n2687 vss.n2686 21.749
R7610 vss.n2756 vss.n2755 21.749
R7611 vss.n5917 vss.n217 21.6672
R7612 vss.t10 vss.n217 21.6672
R7613 vss.n5915 vss.n5914 21.6672
R7614 vss.n5914 vss.t285 21.6672
R7615 vss.n5913 vss.n5912 21.6672
R7616 vss.t285 vss.n5913 21.6672
R7617 vss.n5708 vss.n216 21.6672
R7618 vss.t10 vss.n216 21.6672
R7619 vss.n5394 vss.n754 20.7108
R7620 vss.n5390 vss.n766 20.7108
R7621 vss.n5384 vss.n782 20.7108
R7622 vss.n5380 vss.n799 20.7108
R7623 vss.n5374 vss.n815 20.7108
R7624 vss.n5370 vss.n834 20.7108
R7625 vss.n5364 vss.n847 20.7108
R7626 vss.n5354 vss.n882 20.7108
R7627 vss.n4233 vss.n1293 20.6895
R7628 vss.n4227 vss.n4226 20.6895
R7629 vss.n3024 vss.n3021 20.6895
R7630 vss.n4206 vss.n4205 20.6895
R7631 vss.n3306 vss.t260 20.2931
R7632 vss.n5146 vss.n1115 20.2634
R7633 vss.n5152 vss.n1105 20.2634
R7634 vss.n5158 vss.n1093 20.2634
R7635 vss.n5164 vss.n1081 20.2634
R7636 vss.n5170 vss.n1069 20.2634
R7637 vss.n5176 vss.n1057 20.2634
R7638 vss.n5182 vss.n1045 20.2634
R7639 vss.n5188 vss.n1033 20.2634
R7640 vss.n5201 vss.n1021 20.2634
R7641 vss.n5208 vss.n1009 20.2634
R7642 vss.n5526 vss.n308 20.2634
R7643 vss.n5522 vss.n313 20.2634
R7644 vss.n5518 vss.n327 20.2634
R7645 vss.n5514 vss.n341 20.2634
R7646 vss.n5510 vss.n355 20.2634
R7647 vss.n5506 vss.n369 20.2634
R7648 vss.n5502 vss.n383 20.2634
R7649 vss.n5498 vss.n397 20.2634
R7650 vss.n5494 vss.n411 20.2634
R7651 vss.n5490 vss.n425 20.2634
R7652 vss.n5486 vss.n439 20.2634
R7653 vss.n5482 vss.n453 20.2634
R7654 vss.n5478 vss.n467 20.2634
R7655 vss.n5474 vss.n481 20.2634
R7656 vss.n5470 vss.n495 20.2634
R7657 vss.n5466 vss.n509 20.2634
R7658 vss.n5462 vss.n523 20.2634
R7659 vss.n5458 vss.n537 20.2634
R7660 vss.n5454 vss.n551 20.2634
R7661 vss.n5450 vss.n565 20.2634
R7662 vss.n5446 vss.n579 20.2634
R7663 vss.n5442 vss.n593 20.2634
R7664 vss.n5438 vss.n607 20.2634
R7665 vss.n5434 vss.n621 20.2634
R7666 vss.n5430 vss.n635 20.2634
R7667 vss.n5426 vss.n649 20.2634
R7668 vss.n5422 vss.n663 20.2634
R7669 vss.n5418 vss.n677 20.2634
R7670 vss.n5414 vss.n691 20.2634
R7671 vss.n5410 vss.n705 20.2634
R7672 vss.n5406 vss.n719 20.2634
R7673 vss.n5719 vss.n5708 20.1148
R7674 vss.n2990 vss.n2989 19.8938
R7675 vss.n3306 vss.t195 19.5844
R7676 vss.t42 vss.n2395 19.3956
R7677 vss.n2519 vss.n385 19.0305
R7678 vss.n2633 vss.n2632 19.0305
R7679 vss.n2688 vss.n623 19.0305
R7680 vss.n806 vss.n776 19.0305
R7681 vss.n2318 vss.n1313 18.824
R7682 vss.n2445 vss.n2444 18.4476
R7683 vss.n2227 vss.n2226 18.3023
R7684 vss.n2279 vss.n2278 18.2817
R7685 vss.n2280 vss.n2279 18.2817
R7686 vss.n2276 vss.n2275 18.2817
R7687 vss.n2275 vss.n2274 18.2817
R7688 vss.n5390 vss.n754 18.1851
R7689 vss.n5384 vss.n766 18.1851
R7690 vss.n5380 vss.n782 18.1851
R7691 vss.n5374 vss.n799 18.1851
R7692 vss.n5370 vss.n815 18.1851
R7693 vss.n5364 vss.n834 18.1851
R7694 vss.n5360 vss.n847 18.1851
R7695 vss.n2410 vss.n2396 18.0711
R7696 vss.n2315 vss.n2207 17.6946
R7697 vss.t271 vss.n441 17.6712
R7698 vss.t285 vss.n223 17.6712
R7699 vss.t291 vss.n497 17.6712
R7700 vss.n2609 vss.t27 17.6712
R7701 vss.n3007 vss.n3006 17.5066
R7702 vss.n5666 vss.n5665 16.8234
R7703 vss.n4234 vss.n1291 16.7109
R7704 vss.n2211 vss.n1111 16.7109
R7705 vss.n2194 vss.n1099 16.7109
R7706 vss.n2200 vss.n1087 16.7109
R7707 vss.n2979 vss.n1075 16.7109
R7708 vss.n2330 vss.n1063 16.7109
R7709 vss.n3189 vss.n3187 16.4264
R7710 vss.n3101 vss.n3099 16.4264
R7711 vss.n3106 vss.n3104 16.4264
R7712 vss.n3111 vss.n3109 16.4264
R7713 vss.n3117 vss.n3115 16.4264
R7714 vss.n3123 vss.n3121 16.4264
R7715 vss.n3127 vss.n3125 16.4264
R7716 vss.n3134 vss.n3132 16.4264
R7717 vss.n3140 vss.n3138 16.4264
R7718 vss.n3144 vss.n3142 16.4264
R7719 vss.n3151 vss.n3149 16.4264
R7720 vss.n3157 vss.n3155 16.4264
R7721 vss.n3161 vss.n3159 16.4264
R7722 vss.n3168 vss.n3166 16.4264
R7723 vss.n3174 vss.n3172 16.4264
R7724 vss.n3178 vss.n3176 16.4264
R7725 vss.n3185 vss.n3183 16.4264
R7726 vss.n3194 vss.n3192 16.4264
R7727 vss.n3201 vss.n3199 16.4264
R7728 vss.n3205 vss.n3203 16.4264
R7729 vss.n3212 vss.n3210 16.4264
R7730 vss.n3218 vss.n3216 16.4264
R7731 vss.n3222 vss.n3220 16.4264
R7732 vss.n3229 vss.n3227 16.4264
R7733 vss.n3235 vss.n3233 16.4264
R7734 vss.n3239 vss.n3237 16.4264
R7735 vss.n3246 vss.n3244 16.4264
R7736 vss.n3252 vss.n3250 16.4264
R7737 vss.n3256 vss.n3254 16.4264
R7738 vss.n3263 vss.n3261 16.4264
R7739 vss.n3269 vss.n3267 16.4264
R7740 vss.n3273 vss.n3271 16.4264
R7741 vss.n3280 vss.n3278 16.4264
R7742 vss.n3286 vss.n3284 16.4264
R7743 vss.n3290 vss.n3288 16.4264
R7744 vss.n3297 vss.n3295 16.4264
R7745 vss.n3301 vss.n3299 16.4264
R7746 vss.t284 vss.n2233 16.313
R7747 vss.n2395 vss.n1039 16.3119
R7748 vss.n2512 vss.n2511 16.3119
R7749 vss.n2556 vss.n2555 16.3119
R7750 vss.n5920 vss.n214 16.3119
R7751 vss.n5379 vss.n807 16.3119
R7752 vss.n3189 vss.n3188 15.7177
R7753 vss.n3101 vss.n3100 15.7177
R7754 vss.n3106 vss.n3105 15.7177
R7755 vss.n3111 vss.n3110 15.7177
R7756 vss.n3117 vss.n3116 15.7177
R7757 vss.n3123 vss.n3122 15.7177
R7758 vss.n3127 vss.n3126 15.7177
R7759 vss.n3134 vss.n3133 15.7177
R7760 vss.n3140 vss.n3139 15.7177
R7761 vss.n3144 vss.n3143 15.7177
R7762 vss.n3151 vss.n3150 15.7177
R7763 vss.n3157 vss.n3156 15.7177
R7764 vss.n3161 vss.n3160 15.7177
R7765 vss.n3168 vss.n3167 15.7177
R7766 vss.n3174 vss.n3173 15.7177
R7767 vss.n3178 vss.n3177 15.7177
R7768 vss.n3185 vss.n3184 15.7177
R7769 vss.n3194 vss.n3193 15.7177
R7770 vss.n3201 vss.n3200 15.7177
R7771 vss.n3205 vss.n3204 15.7177
R7772 vss.n3212 vss.n3211 15.7177
R7773 vss.n3218 vss.n3217 15.7177
R7774 vss.n3222 vss.n3221 15.7177
R7775 vss.n3229 vss.n3228 15.7177
R7776 vss.n3235 vss.n3234 15.7177
R7777 vss.n3239 vss.n3238 15.7177
R7778 vss.n3246 vss.n3245 15.7177
R7779 vss.n3252 vss.n3251 15.7177
R7780 vss.n3256 vss.n3255 15.7177
R7781 vss.n3263 vss.n3262 15.7177
R7782 vss.n3269 vss.n3268 15.7177
R7783 vss.n3273 vss.n3272 15.7177
R7784 vss.n3280 vss.n3279 15.7177
R7785 vss.n3286 vss.n3285 15.7177
R7786 vss.n3290 vss.n3289 15.7177
R7787 vss.n3297 vss.n3296 15.7177
R7788 vss.n3301 vss.n3300 15.7177
R7789 vss.n5394 vss.n746 15.1543
R7790 vss.t97 vss.n2270 15.1194
R7791 vss.t169 vss.n2102 15.1194
R7792 vss.t81 vss.n2100 15.1194
R7793 vss.t150 vss.n2098 15.1194
R7794 vss.t87 vss.n2096 15.1194
R7795 vss.t161 vss.n2094 15.1194
R7796 vss.t69 vss.n2092 15.1194
R7797 vss.t143 vss.n2047 15.1194
R7798 vss.t53 vss.n2045 15.1194
R7799 vss.t103 vss.n2043 15.1194
R7800 vss.t101 vss.n2041 15.1194
R7801 vss.t47 vss.n2039 15.1194
R7802 vss.t43 vss.n1994 15.1194
R7803 vss.t123 vss.n1992 15.1194
R7804 vss.t93 vss.n1990 15.1194
R7805 vss.t79 vss.n1988 15.1194
R7806 vss.t77 vss.n1986 15.1194
R7807 vss.t55 vss.n1984 15.1194
R7808 vss.t188 vss.n1935 15.1194
R7809 vss.t71 vss.n1933 15.1194
R7810 vss.t65 vss.n1931 15.1194
R7811 vss.t51 vss.n1929 15.1194
R7812 vss.t49 vss.n1927 15.1194
R7813 vss.t125 vss.n1925 15.1194
R7814 vss.t83 vss.n1880 15.1194
R7815 vss.t157 vss.n1878 15.1194
R7816 vss.t57 vss.n1876 15.1194
R7817 vss.t141 vss.n1874 15.1194
R7818 vss.t135 vss.n1872 15.1194
R7819 vss.t177 vss.n1827 15.1194
R7820 vss.t85 vss.n1825 15.1194
R7821 vss.t131 vss.n1823 15.1194
R7822 vss.t127 vss.n1821 15.1194
R7823 vss.t113 vss.n1819 15.1194
R7824 vss.t91 vss.n1817 15.1194
R7825 vss.t163 vss.n1768 15.1194
R7826 vss.n2252 vss.t73 15.1194
R7827 vss.t147 vss.n2260 15.1194
R7828 vss.t184 vss.n2258 15.1194
R7829 vss.t155 vss.n2256 15.1194
R7830 vss.t61 vss.n2254 15.1194
R7831 vss.t137 vss.n1723 15.1194
R7832 vss.t45 vss.n1721 15.1194
R7833 vss.t117 vss.n1719 15.1194
R7834 vss.t95 vss.n1717 15.1194
R7835 vss.t129 vss.n1715 15.1194
R7836 vss.t200 vss.n1713 15.1194
R7837 vss.t109 vss.n1664 15.1194
R7838 vss.t190 vss.n1662 15.1194
R7839 vss.t159 vss.n1660 15.1194
R7840 vss.t67 vss.n1658 15.1194
R7841 vss.t107 vss.n1656 15.1194
R7842 vss.t182 vss.n1611 15.1194
R7843 vss.t89 vss.n1609 15.1194
R7844 vss.t59 vss.n1607 15.1194
R7845 vss.t133 vss.n1605 15.1194
R7846 vss.t206 vss.n1603 15.1194
R7847 vss.t115 vss.n1601 15.1194
R7848 vss.t167 vss.n1556 15.1194
R7849 vss.t139 vss.n1554 15.1194
R7850 vss.t197 vss.n1552 15.1194
R7851 vss.t119 vss.n1550 15.1194
R7852 vss.t186 vss.n1548 15.1194
R7853 vss.t105 vss.n1546 15.1194
R7854 vss.t63 vss.n1497 15.1194
R7855 vss.t111 vss.n1495 15.1194
R7856 vss.t180 vss.n1493 15.1194
R7857 vss.t99 vss.n1491 15.1194
R7858 vss.t172 vss.n1489 15.1194
R7859 vss.t145 vss.n1444 15.1194
R7860 vss.t203 vss.n1442 15.1194
R7861 vss.t121 vss.n1440 15.1194
R7862 vss.t165 vss.n1438 15.1194
R7863 vss.t75 vss.n1436 15.1194
R7864 vss.t194 vss.n1434 15.1194
R7865 vss.n2421 vss.n2419 15.1194
R7866 vss.n2271 vss.t97 14.3237
R7867 vss.n2269 vss.t169 14.3237
R7868 vss.n2101 vss.t81 14.3237
R7869 vss.n2099 vss.t150 14.3237
R7870 vss.n2097 vss.t87 14.3237
R7871 vss.n2095 vss.t161 14.3237
R7872 vss.n2093 vss.t69 14.3237
R7873 vss.n2048 vss.t143 14.3237
R7874 vss.n2046 vss.t53 14.3237
R7875 vss.n2044 vss.t103 14.3237
R7876 vss.n2042 vss.t101 14.3237
R7877 vss.n2040 vss.t47 14.3237
R7878 vss.n2038 vss.t43 14.3237
R7879 vss.n1993 vss.t123 14.3237
R7880 vss.n1991 vss.t93 14.3237
R7881 vss.n1989 vss.t79 14.3237
R7882 vss.n1987 vss.t77 14.3237
R7883 vss.n1985 vss.t55 14.3237
R7884 vss.n1983 vss.t188 14.3237
R7885 vss.n1934 vss.t71 14.3237
R7886 vss.n1932 vss.t65 14.3237
R7887 vss.n1930 vss.t51 14.3237
R7888 vss.n1928 vss.t49 14.3237
R7889 vss.n1926 vss.t125 14.3237
R7890 vss.n1881 vss.t83 14.3237
R7891 vss.n1879 vss.t157 14.3237
R7892 vss.n1877 vss.t57 14.3237
R7893 vss.n1875 vss.t141 14.3237
R7894 vss.n1873 vss.t135 14.3237
R7895 vss.n1871 vss.t177 14.3237
R7896 vss.n1826 vss.t85 14.3237
R7897 vss.n1824 vss.t131 14.3237
R7898 vss.n1822 vss.t127 14.3237
R7899 vss.n1820 vss.t113 14.3237
R7900 vss.n1818 vss.t91 14.3237
R7901 vss.n1816 vss.t163 14.3237
R7902 vss.t73 vss.n2251 14.3237
R7903 vss.t147 vss.n2253 14.3237
R7904 vss.n2259 vss.t184 14.3237
R7905 vss.n2257 vss.t155 14.3237
R7906 vss.n2255 vss.t61 14.3237
R7907 vss.n1724 vss.t137 14.3237
R7908 vss.n1722 vss.t45 14.3237
R7909 vss.n1720 vss.t117 14.3237
R7910 vss.n1718 vss.t95 14.3237
R7911 vss.n1716 vss.t129 14.3237
R7912 vss.n1714 vss.t200 14.3237
R7913 vss.n1665 vss.t109 14.3237
R7914 vss.n1663 vss.t190 14.3237
R7915 vss.n1661 vss.t159 14.3237
R7916 vss.n1659 vss.t67 14.3237
R7917 vss.n1657 vss.t107 14.3237
R7918 vss.n1655 vss.t182 14.3237
R7919 vss.n1610 vss.t89 14.3237
R7920 vss.n1608 vss.t59 14.3237
R7921 vss.n1606 vss.t133 14.3237
R7922 vss.n1604 vss.t206 14.3237
R7923 vss.n1602 vss.t115 14.3237
R7924 vss.n1557 vss.t167 14.3237
R7925 vss.n1555 vss.t139 14.3237
R7926 vss.n1553 vss.t197 14.3237
R7927 vss.n1551 vss.t119 14.3237
R7928 vss.n1549 vss.t186 14.3237
R7929 vss.n1547 vss.t105 14.3237
R7930 vss.n1498 vss.t63 14.3237
R7931 vss.n1496 vss.t111 14.3237
R7932 vss.n1494 vss.t180 14.3237
R7933 vss.n1492 vss.t99 14.3237
R7934 vss.n1490 vss.t172 14.3237
R7935 vss.n1488 vss.t145 14.3237
R7936 vss.n1443 vss.t203 14.3237
R7937 vss.n1441 vss.t121 14.3237
R7938 vss.n1439 vss.t165 14.3237
R7939 vss.n1437 vss.t75 14.3237
R7940 vss.n1435 vss.t194 14.3237
R7941 vss.n2400 vss.n2399 14.3237
R7942 vss.n2321 vss.n2317 14.3064
R7943 vss.n2412 vss.n2411 13.9299
R7944 vss.n2557 vss.n441 13.5933
R7945 vss.n2653 vss.n567 13.5933
R7946 vss.n2762 vss.n2761 13.5933
R7947 vss.n2412 vss.n2379 13.5534
R7948 vss.n5912 vss.n5911 13.5319
R7949 vss.n2321 vss.n2320 13.177
R7950 vss.n2283 vss.n2282 13.1301
R7951 vss.n5912 vss.n226 12.8005
R7952 vss.n2282 vss.n2281 12.3343
R7953 vss.n2602 vss.t29 12.2341
R7954 vss.t0 vss.n2678 12.2341
R7955 vss.t14 vss.n623 12.2341
R7956 vss.t10 vss.n2706 12.2341
R7957 vss.n2737 vss.t2 12.2341
R7958 vss.n3027 vss.n841 12.2341
R7959 vss.n2223 vss.n2218 12.0952
R7960 vss.n4223 vss.n1308 12.0952
R7961 vss.n2971 vss.n2326 12.0952
R7962 vss.n2403 vss.n2398 12.0952
R7963 vss.n2437 vss.n2382 12.0952
R7964 vss.n5531 vss.n5530 12.0952
R7965 vss.n4234 vss.n4233 11.9365
R7966 vss.n3007 vss.n1063 11.9365
R7967 vss.n2421 vss.n1051 11.9365
R7968 vss.n2418 vss.n2417 11.9365
R7969 vss.n5406 vss.n733 11.5391
R7970 vss.t284 vss.n2234 11.5386
R7971 vss.n2401 vss.n2343 11.5386
R7972 vss.n2643 vss.n2642 10.8748
R7973 vss.n2680 vss.n609 10.8748
R7974 vss.n5388 vss.n5387 10.8748
R7975 vss.n5580 vss.n5579 10.2405
R7976 vss.n5360 vss.n866 10.176
R7977 vss.n895 vss.n879 10.176
R7978 vss.n895 vss.n881 10.176
R7979 vss.n5357 vss.n866 10.176
R7980 vss.n2292 vss.n2238 10.0534
R7981 vss.t41 vss.n2329 9.94715
R7982 vss.n2304 vss.n2207 9.78874
R7983 vss.n1303 vss.n1111 9.54928
R7984 vss.n2989 vss.n2966 9.54928
R7985 vss.n2435 vss.n2433 9.51548
R7986 vss.n2456 vss.t4 9.51548
R7987 vss.n2565 vss.t19 9.51548
R7988 vss.t269 vss.n2581 9.51548
R7989 vss.n2698 vss.t12 9.51548
R7990 vss.t302 vss.n2715 9.51548
R7991 vss.t39 vss.n721 9.51548
R7992 vss.n5665 vss.n5650 9.50907
R7993 vss.n2396 vss.n2334 9.41227
R7994 vss.n4383 vss.n4382 9.38072
R7995 vss.n941 vss.n938 9.3005
R7996 vss.n942 vss.n937 9.3005
R7997 vss.n943 vss.n936 9.3005
R7998 vss.n935 vss.n883 9.3005
R7999 vss.n934 vss.n860 9.3005
R8000 vss.n933 vss.n932 9.3005
R8001 vss.n931 vss.n842 9.3005
R8002 vss.n930 vss.n929 9.3005
R8003 vss.n928 vss.n828 9.3005
R8004 vss.n927 vss.n926 9.3005
R8005 vss.n925 vss.n809 9.3005
R8006 vss.n924 vss.n923 9.3005
R8007 vss.n922 vss.n793 9.3005
R8008 vss.n921 vss.n920 9.3005
R8009 vss.n919 vss.n777 9.3005
R8010 vss.n918 vss.n917 9.3005
R8011 vss.n916 vss.n762 9.3005
R8012 vss.n915 vss.n914 9.3005
R8013 vss.n913 vss.n740 9.3005
R8014 vss.n5404 vss.n739 9.3005
R8015 vss.n5405 vss.n738 9.3005
R8016 vss.n737 vss.n714 9.3005
R8017 vss.n5411 vss.n713 9.3005
R8018 vss.n5412 vss.n712 9.3005
R8019 vss.n5413 vss.n711 9.3005
R8020 vss.n710 vss.n686 9.3005
R8021 vss.n5419 vss.n685 9.3005
R8022 vss.n5420 vss.n684 9.3005
R8023 vss.n5421 vss.n683 9.3005
R8024 vss.n682 vss.n658 9.3005
R8025 vss.n5427 vss.n657 9.3005
R8026 vss.n5428 vss.n656 9.3005
R8027 vss.n5429 vss.n655 9.3005
R8028 vss.n654 vss.n630 9.3005
R8029 vss.n5435 vss.n629 9.3005
R8030 vss.n5436 vss.n628 9.3005
R8031 vss.n5437 vss.n627 9.3005
R8032 vss.n626 vss.n602 9.3005
R8033 vss.n5443 vss.n601 9.3005
R8034 vss.n5444 vss.n600 9.3005
R8035 vss.n5445 vss.n599 9.3005
R8036 vss.n598 vss.n574 9.3005
R8037 vss.n5451 vss.n573 9.3005
R8038 vss.n5452 vss.n572 9.3005
R8039 vss.n5453 vss.n571 9.3005
R8040 vss.n570 vss.n546 9.3005
R8041 vss.n5459 vss.n545 9.3005
R8042 vss.n5460 vss.n544 9.3005
R8043 vss.n5461 vss.n543 9.3005
R8044 vss.n542 vss.n518 9.3005
R8045 vss.n5467 vss.n517 9.3005
R8046 vss.n5468 vss.n516 9.3005
R8047 vss.n5469 vss.n515 9.3005
R8048 vss.n514 vss.n490 9.3005
R8049 vss.n5475 vss.n489 9.3005
R8050 vss.n5476 vss.n488 9.3005
R8051 vss.n5477 vss.n487 9.3005
R8052 vss.n486 vss.n462 9.3005
R8053 vss.n5483 vss.n461 9.3005
R8054 vss.n5484 vss.n460 9.3005
R8055 vss.n5485 vss.n459 9.3005
R8056 vss.n458 vss.n434 9.3005
R8057 vss.n5491 vss.n433 9.3005
R8058 vss.n5492 vss.n432 9.3005
R8059 vss.n5493 vss.n431 9.3005
R8060 vss.n430 vss.n406 9.3005
R8061 vss.n5499 vss.n405 9.3005
R8062 vss.n5500 vss.n404 9.3005
R8063 vss.n5501 vss.n403 9.3005
R8064 vss.n402 vss.n378 9.3005
R8065 vss.n5507 vss.n377 9.3005
R8066 vss.n5508 vss.n376 9.3005
R8067 vss.n5509 vss.n375 9.3005
R8068 vss.n374 vss.n350 9.3005
R8069 vss.n5515 vss.n349 9.3005
R8070 vss.n5516 vss.n348 9.3005
R8071 vss.n5517 vss.n347 9.3005
R8072 vss.n346 vss.n322 9.3005
R8073 vss.n5523 vss.n321 9.3005
R8074 vss.n5524 vss.n320 9.3005
R8075 vss.n5525 vss.n319 9.3005
R8076 vss.n5205 vss.n318 9.3005
R8077 vss.n5207 vss.n5206 9.3005
R8078 vss.n5204 vss.n1018 9.3005
R8079 vss.n5203 vss.n5202 9.3005
R8080 vss.n1020 vss.n1019 9.3005
R8081 vss.n5187 vss.n5186 9.3005
R8082 vss.n5185 vss.n1042 9.3005
R8083 vss.n5184 vss.n5183 9.3005
R8084 vss.n1044 vss.n1043 9.3005
R8085 vss.n5175 vss.n5174 9.3005
R8086 vss.n5173 vss.n1066 9.3005
R8087 vss.n5172 vss.n5171 9.3005
R8088 vss.n1068 vss.n1067 9.3005
R8089 vss.n5163 vss.n5162 9.3005
R8090 vss.n5161 vss.n1090 9.3005
R8091 vss.n5160 vss.n5159 9.3005
R8092 vss.n1092 vss.n1091 9.3005
R8093 vss.n5151 vss.n5150 9.3005
R8094 vss.n5149 vss.n1114 9.3005
R8095 vss.n909 vss.n906 9.3005
R8096 vss.n910 vss.n905 9.3005
R8097 vss.n5355 vss.n904 9.3005
R8098 vss.n5356 vss.n903 9.3005
R8099 vss.n1117 vss.n876 9.3005
R8100 vss.n1119 vss.n1118 9.3005
R8101 vss.n1120 vss.n852 9.3005
R8102 vss.n1122 vss.n1121 9.3005
R8103 vss.n1123 vss.n840 9.3005
R8104 vss.n1125 vss.n1124 9.3005
R8105 vss.n1126 vss.n820 9.3005
R8106 vss.n1128 vss.n1127 9.3005
R8107 vss.n1129 vss.n805 9.3005
R8108 vss.n1131 vss.n1130 9.3005
R8109 vss.n1132 vss.n787 9.3005
R8110 vss.n1134 vss.n1133 9.3005
R8111 vss.n1135 vss.n771 9.3005
R8112 vss.n1137 vss.n1136 9.3005
R8113 vss.n1138 vss.n747 9.3005
R8114 vss.n1139 vss.n741 9.3005
R8115 vss.n1140 vss.n729 9.3005
R8116 vss.n1142 vss.n1141 9.3005
R8117 vss.n1143 vss.n715 9.3005
R8118 vss.n1145 vss.n1144 9.3005
R8119 vss.n1146 vss.n701 9.3005
R8120 vss.n1148 vss.n1147 9.3005
R8121 vss.n1149 vss.n687 9.3005
R8122 vss.n1151 vss.n1150 9.3005
R8123 vss.n1152 vss.n673 9.3005
R8124 vss.n1154 vss.n1153 9.3005
R8125 vss.n1155 vss.n659 9.3005
R8126 vss.n1157 vss.n1156 9.3005
R8127 vss.n1158 vss.n645 9.3005
R8128 vss.n1160 vss.n1159 9.3005
R8129 vss.n1161 vss.n631 9.3005
R8130 vss.n1163 vss.n1162 9.3005
R8131 vss.n1164 vss.n617 9.3005
R8132 vss.n1166 vss.n1165 9.3005
R8133 vss.n1167 vss.n603 9.3005
R8134 vss.n1169 vss.n1168 9.3005
R8135 vss.n1170 vss.n589 9.3005
R8136 vss.n1172 vss.n1171 9.3005
R8137 vss.n1173 vss.n575 9.3005
R8138 vss.n1175 vss.n1174 9.3005
R8139 vss.n1176 vss.n561 9.3005
R8140 vss.n1178 vss.n1177 9.3005
R8141 vss.n1179 vss.n547 9.3005
R8142 vss.n1181 vss.n1180 9.3005
R8143 vss.n1182 vss.n533 9.3005
R8144 vss.n1184 vss.n1183 9.3005
R8145 vss.n1185 vss.n519 9.3005
R8146 vss.n1187 vss.n1186 9.3005
R8147 vss.n1188 vss.n505 9.3005
R8148 vss.n1190 vss.n1189 9.3005
R8149 vss.n1191 vss.n491 9.3005
R8150 vss.n1193 vss.n1192 9.3005
R8151 vss.n1194 vss.n477 9.3005
R8152 vss.n1196 vss.n1195 9.3005
R8153 vss.n1197 vss.n463 9.3005
R8154 vss.n1199 vss.n1198 9.3005
R8155 vss.n1200 vss.n449 9.3005
R8156 vss.n1202 vss.n1201 9.3005
R8157 vss.n1203 vss.n435 9.3005
R8158 vss.n1205 vss.n1204 9.3005
R8159 vss.n1206 vss.n421 9.3005
R8160 vss.n1208 vss.n1207 9.3005
R8161 vss.n1209 vss.n407 9.3005
R8162 vss.n1211 vss.n1210 9.3005
R8163 vss.n1212 vss.n393 9.3005
R8164 vss.n1214 vss.n1213 9.3005
R8165 vss.n1215 vss.n379 9.3005
R8166 vss.n1217 vss.n1216 9.3005
R8167 vss.n1218 vss.n365 9.3005
R8168 vss.n1220 vss.n1219 9.3005
R8169 vss.n1221 vss.n351 9.3005
R8170 vss.n1223 vss.n1222 9.3005
R8171 vss.n1224 vss.n337 9.3005
R8172 vss.n1226 vss.n1225 9.3005
R8173 vss.n1227 vss.n323 9.3005
R8174 vss.n1229 vss.n1228 9.3005
R8175 vss.n1230 vss.n309 9.3005
R8176 vss.n1232 vss.n1231 9.3005
R8177 vss.n1233 vss.n1010 9.3005
R8178 vss.n1235 vss.n1234 9.3005
R8179 vss.n1236 vss.n1022 9.3005
R8180 vss.n1238 vss.n1237 9.3005
R8181 vss.n1239 vss.n1034 9.3005
R8182 vss.n1241 vss.n1240 9.3005
R8183 vss.n1242 vss.n1046 9.3005
R8184 vss.n1244 vss.n1243 9.3005
R8185 vss.n1245 vss.n1058 9.3005
R8186 vss.n1247 vss.n1246 9.3005
R8187 vss.n1248 vss.n1070 9.3005
R8188 vss.n1250 vss.n1249 9.3005
R8189 vss.n1251 vss.n1082 9.3005
R8190 vss.n1253 vss.n1252 9.3005
R8191 vss.n1254 vss.n1094 9.3005
R8192 vss.n1256 vss.n1255 9.3005
R8193 vss.n1257 vss.n1106 9.3005
R8194 vss.n1259 vss.n1258 9.3005
R8195 vss.n967 vss.n964 9.3005
R8196 vss.n968 vss.n963 9.3005
R8197 vss.n969 vss.n962 9.3005
R8198 vss.n961 vss.n884 9.3005
R8199 vss.n960 vss.n861 9.3005
R8200 vss.n959 vss.n958 9.3005
R8201 vss.n957 vss.n843 9.3005
R8202 vss.n956 vss.n955 9.3005
R8203 vss.n954 vss.n829 9.3005
R8204 vss.n953 vss.n952 9.3005
R8205 vss.n951 vss.n810 9.3005
R8206 vss.n950 vss.n949 9.3005
R8207 vss.n948 vss.n794 9.3005
R8208 vss.n947 vss.n946 9.3005
R8209 vss.n945 vss.n778 9.3005
R8210 vss.n944 vss.n761 9.3005
R8211 vss.n5391 vss.n760 9.3005
R8212 vss.n5392 vss.n759 9.3005
R8213 vss.n5393 vss.n758 9.3005
R8214 vss.n757 vss.n728 9.3005
R8215 vss.n5407 vss.n727 9.3005
R8216 vss.n5408 vss.n726 9.3005
R8217 vss.n5409 vss.n725 9.3005
R8218 vss.n724 vss.n700 9.3005
R8219 vss.n5415 vss.n699 9.3005
R8220 vss.n5416 vss.n698 9.3005
R8221 vss.n5417 vss.n697 9.3005
R8222 vss.n696 vss.n672 9.3005
R8223 vss.n5423 vss.n671 9.3005
R8224 vss.n5424 vss.n670 9.3005
R8225 vss.n5425 vss.n669 9.3005
R8226 vss.n668 vss.n644 9.3005
R8227 vss.n5431 vss.n643 9.3005
R8228 vss.n5432 vss.n642 9.3005
R8229 vss.n5433 vss.n641 9.3005
R8230 vss.n640 vss.n616 9.3005
R8231 vss.n5439 vss.n615 9.3005
R8232 vss.n5440 vss.n614 9.3005
R8233 vss.n5441 vss.n613 9.3005
R8234 vss.n612 vss.n588 9.3005
R8235 vss.n5447 vss.n587 9.3005
R8236 vss.n5448 vss.n586 9.3005
R8237 vss.n5449 vss.n585 9.3005
R8238 vss.n584 vss.n560 9.3005
R8239 vss.n5455 vss.n559 9.3005
R8240 vss.n5456 vss.n558 9.3005
R8241 vss.n5457 vss.n557 9.3005
R8242 vss.n556 vss.n532 9.3005
R8243 vss.n5463 vss.n531 9.3005
R8244 vss.n5464 vss.n530 9.3005
R8245 vss.n5465 vss.n529 9.3005
R8246 vss.n528 vss.n504 9.3005
R8247 vss.n5471 vss.n503 9.3005
R8248 vss.n5472 vss.n502 9.3005
R8249 vss.n5473 vss.n501 9.3005
R8250 vss.n500 vss.n476 9.3005
R8251 vss.n5479 vss.n475 9.3005
R8252 vss.n5480 vss.n474 9.3005
R8253 vss.n5481 vss.n473 9.3005
R8254 vss.n472 vss.n448 9.3005
R8255 vss.n5487 vss.n447 9.3005
R8256 vss.n5488 vss.n446 9.3005
R8257 vss.n5489 vss.n445 9.3005
R8258 vss.n444 vss.n420 9.3005
R8259 vss.n5495 vss.n419 9.3005
R8260 vss.n5496 vss.n418 9.3005
R8261 vss.n5497 vss.n417 9.3005
R8262 vss.n416 vss.n392 9.3005
R8263 vss.n5503 vss.n391 9.3005
R8264 vss.n5504 vss.n390 9.3005
R8265 vss.n5505 vss.n389 9.3005
R8266 vss.n388 vss.n364 9.3005
R8267 vss.n5511 vss.n363 9.3005
R8268 vss.n5512 vss.n362 9.3005
R8269 vss.n5513 vss.n361 9.3005
R8270 vss.n360 vss.n336 9.3005
R8271 vss.n5519 vss.n335 9.3005
R8272 vss.n5520 vss.n334 9.3005
R8273 vss.n5521 vss.n333 9.3005
R8274 vss.n5193 vss.n332 9.3005
R8275 vss.n5194 vss.n317 9.3005
R8276 vss.n5196 vss.n5195 9.3005
R8277 vss.n5197 vss.n1017 9.3005
R8278 vss.n5199 vss.n5198 9.3005
R8279 vss.n5200 vss.n5192 9.3005
R8280 vss.n5191 vss.n1030 9.3005
R8281 vss.n5190 vss.n5189 9.3005
R8282 vss.n1032 vss.n1031 9.3005
R8283 vss.n5181 vss.n5180 9.3005
R8284 vss.n5179 vss.n1054 9.3005
R8285 vss.n5178 vss.n5177 9.3005
R8286 vss.n1056 vss.n1055 9.3005
R8287 vss.n5169 vss.n5168 9.3005
R8288 vss.n5167 vss.n1078 9.3005
R8289 vss.n5166 vss.n5165 9.3005
R8290 vss.n1080 vss.n1079 9.3005
R8291 vss.n5157 vss.n5156 9.3005
R8292 vss.n5155 vss.n1102 9.3005
R8293 vss.n5154 vss.n5153 9.3005
R8294 vss.n1104 vss.n1103 9.3005
R8295 vss.n5332 vss.n5329 9.3005
R8296 vss.n5333 vss.n5328 9.3005
R8297 vss.n5334 vss.n5327 9.3005
R8298 vss.n5326 vss.n901 9.3005
R8299 vss.n5325 vss.n874 9.3005
R8300 vss.n5324 vss.n5323 9.3005
R8301 vss.n5322 vss.n851 9.3005
R8302 vss.n5321 vss.n5320 9.3005
R8303 vss.n5319 vss.n839 9.3005
R8304 vss.n5318 vss.n5317 9.3005
R8305 vss.n5316 vss.n819 9.3005
R8306 vss.n5315 vss.n5314 9.3005
R8307 vss.n5313 vss.n804 9.3005
R8308 vss.n5312 vss.n5311 9.3005
R8309 vss.n5310 vss.n786 9.3005
R8310 vss.n5309 vss.n5308 9.3005
R8311 vss.n5307 vss.n770 9.3005
R8312 vss.n5306 vss.n5305 9.3005
R8313 vss.n5304 vss.n748 9.3005
R8314 vss.n5303 vss.n742 9.3005
R8315 vss.n5302 vss.n730 9.3005
R8316 vss.n5301 vss.n5300 9.3005
R8317 vss.n5299 vss.n716 9.3005
R8318 vss.n5298 vss.n5297 9.3005
R8319 vss.n5296 vss.n702 9.3005
R8320 vss.n5295 vss.n5294 9.3005
R8321 vss.n5293 vss.n688 9.3005
R8322 vss.n5292 vss.n5291 9.3005
R8323 vss.n5290 vss.n674 9.3005
R8324 vss.n5289 vss.n5288 9.3005
R8325 vss.n5287 vss.n660 9.3005
R8326 vss.n5286 vss.n5285 9.3005
R8327 vss.n5284 vss.n646 9.3005
R8328 vss.n5283 vss.n5282 9.3005
R8329 vss.n5281 vss.n632 9.3005
R8330 vss.n5280 vss.n5279 9.3005
R8331 vss.n5278 vss.n618 9.3005
R8332 vss.n5277 vss.n5276 9.3005
R8333 vss.n5275 vss.n604 9.3005
R8334 vss.n5274 vss.n5273 9.3005
R8335 vss.n5272 vss.n590 9.3005
R8336 vss.n5271 vss.n5270 9.3005
R8337 vss.n5269 vss.n576 9.3005
R8338 vss.n5268 vss.n5267 9.3005
R8339 vss.n5266 vss.n562 9.3005
R8340 vss.n5265 vss.n5264 9.3005
R8341 vss.n5263 vss.n548 9.3005
R8342 vss.n5262 vss.n5261 9.3005
R8343 vss.n5260 vss.n534 9.3005
R8344 vss.n5259 vss.n5258 9.3005
R8345 vss.n5257 vss.n520 9.3005
R8346 vss.n5256 vss.n5255 9.3005
R8347 vss.n5254 vss.n506 9.3005
R8348 vss.n5253 vss.n5252 9.3005
R8349 vss.n5251 vss.n492 9.3005
R8350 vss.n5250 vss.n5249 9.3005
R8351 vss.n5248 vss.n478 9.3005
R8352 vss.n5247 vss.n5246 9.3005
R8353 vss.n5245 vss.n464 9.3005
R8354 vss.n5244 vss.n5243 9.3005
R8355 vss.n5242 vss.n450 9.3005
R8356 vss.n5241 vss.n5240 9.3005
R8357 vss.n5239 vss.n436 9.3005
R8358 vss.n5238 vss.n5237 9.3005
R8359 vss.n5236 vss.n422 9.3005
R8360 vss.n5235 vss.n5234 9.3005
R8361 vss.n5233 vss.n408 9.3005
R8362 vss.n5232 vss.n5231 9.3005
R8363 vss.n5230 vss.n394 9.3005
R8364 vss.n5229 vss.n5228 9.3005
R8365 vss.n5227 vss.n380 9.3005
R8366 vss.n5226 vss.n5225 9.3005
R8367 vss.n5224 vss.n366 9.3005
R8368 vss.n5223 vss.n5222 9.3005
R8369 vss.n5221 vss.n352 9.3005
R8370 vss.n5220 vss.n5219 9.3005
R8371 vss.n5218 vss.n338 9.3005
R8372 vss.n5217 vss.n5216 9.3005
R8373 vss.n5215 vss.n324 9.3005
R8374 vss.n5214 vss.n5213 9.3005
R8375 vss.n5212 vss.n310 9.3005
R8376 vss.n5211 vss.n5210 9.3005
R8377 vss.n5209 vss.n1007 9.3005
R8378 vss.n1262 vss.n1008 9.3005
R8379 vss.n1263 vss.n1023 9.3005
R8380 vss.n1265 vss.n1264 9.3005
R8381 vss.n1266 vss.n1035 9.3005
R8382 vss.n1268 vss.n1267 9.3005
R8383 vss.n1269 vss.n1047 9.3005
R8384 vss.n1271 vss.n1270 9.3005
R8385 vss.n1272 vss.n1059 9.3005
R8386 vss.n1274 vss.n1273 9.3005
R8387 vss.n1275 vss.n1071 9.3005
R8388 vss.n1277 vss.n1276 9.3005
R8389 vss.n1278 vss.n1083 9.3005
R8390 vss.n1280 vss.n1279 9.3005
R8391 vss.n1281 vss.n1095 9.3005
R8392 vss.n1283 vss.n1282 9.3005
R8393 vss.n1284 vss.n1107 9.3005
R8394 vss.n1286 vss.n1285 9.3005
R8395 vss.n997 vss.n994 9.3005
R8396 vss.n998 vss.n993 9.3005
R8397 vss.n999 vss.n992 9.3005
R8398 vss.n991 vss.n886 9.3005
R8399 vss.n990 vss.n862 9.3005
R8400 vss.n989 vss.n988 9.3005
R8401 vss.n987 vss.n844 9.3005
R8402 vss.n986 vss.n985 9.3005
R8403 vss.n984 vss.n830 9.3005
R8404 vss.n983 vss.n982 9.3005
R8405 vss.n981 vss.n811 9.3005
R8406 vss.n980 vss.n979 9.3005
R8407 vss.n978 vss.n795 9.3005
R8408 vss.n977 vss.n976 9.3005
R8409 vss.n975 vss.n779 9.3005
R8410 vss.n974 vss.n973 9.3005
R8411 vss.n972 vss.n763 9.3005
R8412 vss.n971 vss.n745 9.3005
R8413 vss.n5395 vss.n744 9.3005
R8414 vss.n5396 vss.n743 9.3005
R8415 vss.n5023 vss.n736 9.3005
R8416 vss.n5025 vss.n5024 9.3005
R8417 vss.n5026 vss.n723 9.3005
R8418 vss.n5028 vss.n5027 9.3005
R8419 vss.n5029 vss.n709 9.3005
R8420 vss.n5031 vss.n5030 9.3005
R8421 vss.n5032 vss.n695 9.3005
R8422 vss.n5034 vss.n5033 9.3005
R8423 vss.n5035 vss.n681 9.3005
R8424 vss.n5037 vss.n5036 9.3005
R8425 vss.n5038 vss.n667 9.3005
R8426 vss.n5040 vss.n5039 9.3005
R8427 vss.n5041 vss.n653 9.3005
R8428 vss.n5043 vss.n5042 9.3005
R8429 vss.n5044 vss.n639 9.3005
R8430 vss.n5046 vss.n5045 9.3005
R8431 vss.n5047 vss.n625 9.3005
R8432 vss.n5049 vss.n5048 9.3005
R8433 vss.n5050 vss.n611 9.3005
R8434 vss.n5052 vss.n5051 9.3005
R8435 vss.n5053 vss.n597 9.3005
R8436 vss.n5055 vss.n5054 9.3005
R8437 vss.n5056 vss.n583 9.3005
R8438 vss.n5058 vss.n5057 9.3005
R8439 vss.n5059 vss.n569 9.3005
R8440 vss.n5061 vss.n5060 9.3005
R8441 vss.n5062 vss.n555 9.3005
R8442 vss.n5064 vss.n5063 9.3005
R8443 vss.n5065 vss.n541 9.3005
R8444 vss.n5067 vss.n5066 9.3005
R8445 vss.n5068 vss.n527 9.3005
R8446 vss.n5070 vss.n5069 9.3005
R8447 vss.n5071 vss.n513 9.3005
R8448 vss.n5073 vss.n5072 9.3005
R8449 vss.n5074 vss.n499 9.3005
R8450 vss.n5076 vss.n5075 9.3005
R8451 vss.n5077 vss.n485 9.3005
R8452 vss.n5079 vss.n5078 9.3005
R8453 vss.n5080 vss.n471 9.3005
R8454 vss.n5082 vss.n5081 9.3005
R8455 vss.n5083 vss.n457 9.3005
R8456 vss.n5085 vss.n5084 9.3005
R8457 vss.n5086 vss.n443 9.3005
R8458 vss.n5088 vss.n5087 9.3005
R8459 vss.n5089 vss.n429 9.3005
R8460 vss.n5091 vss.n5090 9.3005
R8461 vss.n5092 vss.n415 9.3005
R8462 vss.n5094 vss.n5093 9.3005
R8463 vss.n5095 vss.n401 9.3005
R8464 vss.n5097 vss.n5096 9.3005
R8465 vss.n5098 vss.n387 9.3005
R8466 vss.n5100 vss.n5099 9.3005
R8467 vss.n5101 vss.n373 9.3005
R8468 vss.n5103 vss.n5102 9.3005
R8469 vss.n5104 vss.n359 9.3005
R8470 vss.n5106 vss.n5105 9.3005
R8471 vss.n5107 vss.n345 9.3005
R8472 vss.n5109 vss.n5108 9.3005
R8473 vss.n5110 vss.n331 9.3005
R8474 vss.n5112 vss.n5111 9.3005
R8475 vss.n5113 vss.n316 9.3005
R8476 vss.n5115 vss.n5114 9.3005
R8477 vss.n5116 vss.n1016 9.3005
R8478 vss.n5118 vss.n5117 9.3005
R8479 vss.n5119 vss.n1029 9.3005
R8480 vss.n5121 vss.n5120 9.3005
R8481 vss.n5122 vss.n1041 9.3005
R8482 vss.n5124 vss.n5123 9.3005
R8483 vss.n5125 vss.n1053 9.3005
R8484 vss.n5127 vss.n5126 9.3005
R8485 vss.n5128 vss.n1065 9.3005
R8486 vss.n5130 vss.n5129 9.3005
R8487 vss.n5131 vss.n1077 9.3005
R8488 vss.n5133 vss.n5132 9.3005
R8489 vss.n5134 vss.n1089 9.3005
R8490 vss.n5136 vss.n5135 9.3005
R8491 vss.n5137 vss.n1101 9.3005
R8492 vss.n5139 vss.n5138 9.3005
R8493 vss.n5140 vss.n1113 9.3005
R8494 vss.n5142 vss.n5141 9.3005
R8495 vss.n4867 vss.n4864 9.3005
R8496 vss.n4869 vss.n4868 9.3005
R8497 vss.n4870 vss.n1006 9.3005
R8498 vss.n4871 vss.n899 9.3005
R8499 vss.n4872 vss.n872 9.3005
R8500 vss.n4874 vss.n4873 9.3005
R8501 vss.n4875 vss.n850 9.3005
R8502 vss.n4877 vss.n4876 9.3005
R8503 vss.n4878 vss.n838 9.3005
R8504 vss.n4880 vss.n4879 9.3005
R8505 vss.n4881 vss.n818 9.3005
R8506 vss.n4883 vss.n4882 9.3005
R8507 vss.n4884 vss.n803 9.3005
R8508 vss.n4886 vss.n4885 9.3005
R8509 vss.n4887 vss.n785 9.3005
R8510 vss.n4889 vss.n4888 9.3005
R8511 vss.n4890 vss.n769 9.3005
R8512 vss.n4892 vss.n4891 9.3005
R8513 vss.n4893 vss.n749 9.3005
R8514 vss.n4895 vss.n4894 9.3005
R8515 vss.n4863 vss.n731 9.3005
R8516 vss.n4862 vss.n4861 9.3005
R8517 vss.n4860 vss.n717 9.3005
R8518 vss.n4859 vss.n4858 9.3005
R8519 vss.n4857 vss.n703 9.3005
R8520 vss.n4856 vss.n4855 9.3005
R8521 vss.n4854 vss.n689 9.3005
R8522 vss.n4853 vss.n4852 9.3005
R8523 vss.n4851 vss.n675 9.3005
R8524 vss.n4850 vss.n4849 9.3005
R8525 vss.n4848 vss.n661 9.3005
R8526 vss.n4847 vss.n4846 9.3005
R8527 vss.n4845 vss.n647 9.3005
R8528 vss.n4844 vss.n4843 9.3005
R8529 vss.n4842 vss.n633 9.3005
R8530 vss.n4841 vss.n4840 9.3005
R8531 vss.n4839 vss.n619 9.3005
R8532 vss.n4838 vss.n4837 9.3005
R8533 vss.n4836 vss.n605 9.3005
R8534 vss.n4835 vss.n4834 9.3005
R8535 vss.n4833 vss.n591 9.3005
R8536 vss.n4832 vss.n4831 9.3005
R8537 vss.n4830 vss.n577 9.3005
R8538 vss.n4829 vss.n4828 9.3005
R8539 vss.n4827 vss.n563 9.3005
R8540 vss.n4826 vss.n4825 9.3005
R8541 vss.n4824 vss.n549 9.3005
R8542 vss.n4823 vss.n4822 9.3005
R8543 vss.n4821 vss.n535 9.3005
R8544 vss.n4820 vss.n4819 9.3005
R8545 vss.n4818 vss.n521 9.3005
R8546 vss.n4817 vss.n4816 9.3005
R8547 vss.n4815 vss.n507 9.3005
R8548 vss.n4814 vss.n4813 9.3005
R8549 vss.n4812 vss.n493 9.3005
R8550 vss.n4811 vss.n4810 9.3005
R8551 vss.n4809 vss.n479 9.3005
R8552 vss.n4808 vss.n4807 9.3005
R8553 vss.n4806 vss.n465 9.3005
R8554 vss.n4805 vss.n4804 9.3005
R8555 vss.n4803 vss.n451 9.3005
R8556 vss.n4802 vss.n4801 9.3005
R8557 vss.n4800 vss.n437 9.3005
R8558 vss.n4799 vss.n4798 9.3005
R8559 vss.n4797 vss.n423 9.3005
R8560 vss.n4796 vss.n4795 9.3005
R8561 vss.n4794 vss.n409 9.3005
R8562 vss.n4793 vss.n4792 9.3005
R8563 vss.n4791 vss.n395 9.3005
R8564 vss.n4790 vss.n4789 9.3005
R8565 vss.n4788 vss.n381 9.3005
R8566 vss.n4787 vss.n4786 9.3005
R8567 vss.n4785 vss.n367 9.3005
R8568 vss.n4784 vss.n4783 9.3005
R8569 vss.n4782 vss.n353 9.3005
R8570 vss.n4781 vss.n4780 9.3005
R8571 vss.n4779 vss.n339 9.3005
R8572 vss.n4778 vss.n4777 9.3005
R8573 vss.n4776 vss.n325 9.3005
R8574 vss.n4775 vss.n4774 9.3005
R8575 vss.n4773 vss.n311 9.3005
R8576 vss.n4772 vss.n4771 9.3005
R8577 vss.n4770 vss.n1011 9.3005
R8578 vss.n4769 vss.n4768 9.3005
R8579 vss.n4767 vss.n1024 9.3005
R8580 vss.n4766 vss.n4765 9.3005
R8581 vss.n4764 vss.n1036 9.3005
R8582 vss.n4763 vss.n4762 9.3005
R8583 vss.n4761 vss.n1048 9.3005
R8584 vss.n4760 vss.n4759 9.3005
R8585 vss.n4758 vss.n1060 9.3005
R8586 vss.n4757 vss.n4756 9.3005
R8587 vss.n4755 vss.n1072 9.3005
R8588 vss.n4754 vss.n4753 9.3005
R8589 vss.n4752 vss.n1084 9.3005
R8590 vss.n4751 vss.n4750 9.3005
R8591 vss.n4749 vss.n1096 9.3005
R8592 vss.n4748 vss.n4747 9.3005
R8593 vss.n4746 vss.n1108 9.3005
R8594 vss.n4745 vss.n4744 9.3005
R8595 vss.n4239 vss.n4236 9.3005
R8596 vss.n4241 vss.n4240 9.3005
R8597 vss.n4242 vss.n1001 9.3005
R8598 vss.n4243 vss.n888 9.3005
R8599 vss.n4244 vss.n863 9.3005
R8600 vss.n4246 vss.n4245 9.3005
R8601 vss.n4247 vss.n845 9.3005
R8602 vss.n4249 vss.n4248 9.3005
R8603 vss.n4250 vss.n831 9.3005
R8604 vss.n4252 vss.n4251 9.3005
R8605 vss.n4253 vss.n812 9.3005
R8606 vss.n4255 vss.n4254 9.3005
R8607 vss.n4256 vss.n796 9.3005
R8608 vss.n4258 vss.n4257 9.3005
R8609 vss.n4259 vss.n780 9.3005
R8610 vss.n4261 vss.n4260 9.3005
R8611 vss.n4262 vss.n764 9.3005
R8612 vss.n4264 vss.n4263 9.3005
R8613 vss.n4265 vss.n756 9.3005
R8614 vss.n4900 vss.n4899 9.3005
R8615 vss.n4901 vss.n735 9.3005
R8616 vss.n4903 vss.n4902 9.3005
R8617 vss.n4904 vss.n722 9.3005
R8618 vss.n4906 vss.n4905 9.3005
R8619 vss.n4907 vss.n708 9.3005
R8620 vss.n4909 vss.n4908 9.3005
R8621 vss.n4910 vss.n694 9.3005
R8622 vss.n4912 vss.n4911 9.3005
R8623 vss.n4913 vss.n680 9.3005
R8624 vss.n4915 vss.n4914 9.3005
R8625 vss.n4916 vss.n666 9.3005
R8626 vss.n4918 vss.n4917 9.3005
R8627 vss.n4919 vss.n652 9.3005
R8628 vss.n4921 vss.n4920 9.3005
R8629 vss.n4922 vss.n638 9.3005
R8630 vss.n4924 vss.n4923 9.3005
R8631 vss.n4925 vss.n624 9.3005
R8632 vss.n4927 vss.n4926 9.3005
R8633 vss.n4928 vss.n610 9.3005
R8634 vss.n4930 vss.n4929 9.3005
R8635 vss.n4931 vss.n596 9.3005
R8636 vss.n4933 vss.n4932 9.3005
R8637 vss.n4934 vss.n582 9.3005
R8638 vss.n4936 vss.n4935 9.3005
R8639 vss.n4937 vss.n568 9.3005
R8640 vss.n4939 vss.n4938 9.3005
R8641 vss.n4940 vss.n554 9.3005
R8642 vss.n4942 vss.n4941 9.3005
R8643 vss.n4943 vss.n540 9.3005
R8644 vss.n4945 vss.n4944 9.3005
R8645 vss.n4946 vss.n526 9.3005
R8646 vss.n4948 vss.n4947 9.3005
R8647 vss.n4949 vss.n512 9.3005
R8648 vss.n4951 vss.n4950 9.3005
R8649 vss.n4952 vss.n498 9.3005
R8650 vss.n4954 vss.n4953 9.3005
R8651 vss.n4955 vss.n484 9.3005
R8652 vss.n4957 vss.n4956 9.3005
R8653 vss.n4958 vss.n470 9.3005
R8654 vss.n4960 vss.n4959 9.3005
R8655 vss.n4961 vss.n456 9.3005
R8656 vss.n4963 vss.n4962 9.3005
R8657 vss.n4964 vss.n442 9.3005
R8658 vss.n4966 vss.n4965 9.3005
R8659 vss.n4967 vss.n428 9.3005
R8660 vss.n4969 vss.n4968 9.3005
R8661 vss.n4970 vss.n414 9.3005
R8662 vss.n4972 vss.n4971 9.3005
R8663 vss.n4973 vss.n400 9.3005
R8664 vss.n4975 vss.n4974 9.3005
R8665 vss.n4976 vss.n386 9.3005
R8666 vss.n4978 vss.n4977 9.3005
R8667 vss.n4979 vss.n372 9.3005
R8668 vss.n4981 vss.n4980 9.3005
R8669 vss.n4982 vss.n358 9.3005
R8670 vss.n4984 vss.n4983 9.3005
R8671 vss.n4985 vss.n344 9.3005
R8672 vss.n4987 vss.n4986 9.3005
R8673 vss.n4988 vss.n330 9.3005
R8674 vss.n4990 vss.n4989 9.3005
R8675 vss.n4991 vss.n315 9.3005
R8676 vss.n4993 vss.n4992 9.3005
R8677 vss.n4994 vss.n1015 9.3005
R8678 vss.n4996 vss.n4995 9.3005
R8679 vss.n4997 vss.n1028 9.3005
R8680 vss.n4999 vss.n4998 9.3005
R8681 vss.n5000 vss.n1040 9.3005
R8682 vss.n5002 vss.n5001 9.3005
R8683 vss.n5003 vss.n1052 9.3005
R8684 vss.n5005 vss.n5004 9.3005
R8685 vss.n5006 vss.n1064 9.3005
R8686 vss.n5008 vss.n5007 9.3005
R8687 vss.n5009 vss.n1076 9.3005
R8688 vss.n5011 vss.n5010 9.3005
R8689 vss.n5012 vss.n1088 9.3005
R8690 vss.n5014 vss.n5013 9.3005
R8691 vss.n5015 vss.n1100 9.3005
R8692 vss.n5017 vss.n5016 9.3005
R8693 vss.n5018 vss.n1112 9.3005
R8694 vss.n5020 vss.n5019 9.3005
R8695 vss.n4713 vss.n4710 9.3005
R8696 vss.n4715 vss.n4714 9.3005
R8697 vss.n4716 vss.n1005 9.3005
R8698 vss.n4717 vss.n897 9.3005
R8699 vss.n4718 vss.n870 9.3005
R8700 vss.n4720 vss.n4719 9.3005
R8701 vss.n4721 vss.n849 9.3005
R8702 vss.n4723 vss.n4722 9.3005
R8703 vss.n4724 vss.n837 9.3005
R8704 vss.n4726 vss.n4725 9.3005
R8705 vss.n4727 vss.n817 9.3005
R8706 vss.n4729 vss.n4728 9.3005
R8707 vss.n4730 vss.n802 9.3005
R8708 vss.n4732 vss.n4731 9.3005
R8709 vss.n4733 vss.n784 9.3005
R8710 vss.n4735 vss.n4734 9.3005
R8711 vss.n4736 vss.n768 9.3005
R8712 vss.n4738 vss.n4737 9.3005
R8713 vss.n4739 vss.n750 9.3005
R8714 vss.n4741 vss.n4740 9.3005
R8715 vss.n4709 vss.n732 9.3005
R8716 vss.n4708 vss.n4707 9.3005
R8717 vss.n4706 vss.n718 9.3005
R8718 vss.n4705 vss.n4704 9.3005
R8719 vss.n4703 vss.n704 9.3005
R8720 vss.n4702 vss.n4701 9.3005
R8721 vss.n4700 vss.n690 9.3005
R8722 vss.n4699 vss.n4698 9.3005
R8723 vss.n4697 vss.n676 9.3005
R8724 vss.n4696 vss.n4695 9.3005
R8725 vss.n4694 vss.n662 9.3005
R8726 vss.n4693 vss.n4692 9.3005
R8727 vss.n4691 vss.n648 9.3005
R8728 vss.n4690 vss.n4689 9.3005
R8729 vss.n4688 vss.n634 9.3005
R8730 vss.n4687 vss.n4686 9.3005
R8731 vss.n4685 vss.n620 9.3005
R8732 vss.n4684 vss.n4683 9.3005
R8733 vss.n4682 vss.n606 9.3005
R8734 vss.n4681 vss.n4680 9.3005
R8735 vss.n4679 vss.n592 9.3005
R8736 vss.n4678 vss.n4677 9.3005
R8737 vss.n4676 vss.n578 9.3005
R8738 vss.n4675 vss.n4674 9.3005
R8739 vss.n4673 vss.n564 9.3005
R8740 vss.n4672 vss.n4671 9.3005
R8741 vss.n4670 vss.n550 9.3005
R8742 vss.n4669 vss.n4668 9.3005
R8743 vss.n4667 vss.n536 9.3005
R8744 vss.n4666 vss.n4665 9.3005
R8745 vss.n4664 vss.n522 9.3005
R8746 vss.n4663 vss.n4662 9.3005
R8747 vss.n4661 vss.n508 9.3005
R8748 vss.n4660 vss.n4659 9.3005
R8749 vss.n4658 vss.n494 9.3005
R8750 vss.n4657 vss.n4656 9.3005
R8751 vss.n4655 vss.n480 9.3005
R8752 vss.n4654 vss.n4653 9.3005
R8753 vss.n4652 vss.n466 9.3005
R8754 vss.n4651 vss.n4650 9.3005
R8755 vss.n4649 vss.n452 9.3005
R8756 vss.n4648 vss.n4647 9.3005
R8757 vss.n4646 vss.n438 9.3005
R8758 vss.n4645 vss.n4644 9.3005
R8759 vss.n4643 vss.n424 9.3005
R8760 vss.n4642 vss.n4641 9.3005
R8761 vss.n4640 vss.n410 9.3005
R8762 vss.n4639 vss.n4638 9.3005
R8763 vss.n4637 vss.n396 9.3005
R8764 vss.n4636 vss.n4635 9.3005
R8765 vss.n4634 vss.n382 9.3005
R8766 vss.n4633 vss.n4632 9.3005
R8767 vss.n4631 vss.n368 9.3005
R8768 vss.n4630 vss.n4629 9.3005
R8769 vss.n4628 vss.n354 9.3005
R8770 vss.n4627 vss.n4626 9.3005
R8771 vss.n4625 vss.n340 9.3005
R8772 vss.n4624 vss.n4623 9.3005
R8773 vss.n4622 vss.n326 9.3005
R8774 vss.n4621 vss.n4620 9.3005
R8775 vss.n4619 vss.n312 9.3005
R8776 vss.n4618 vss.n4617 9.3005
R8777 vss.n4616 vss.n1012 9.3005
R8778 vss.n4615 vss.n4614 9.3005
R8779 vss.n4613 vss.n1025 9.3005
R8780 vss.n4612 vss.n4611 9.3005
R8781 vss.n4610 vss.n1037 9.3005
R8782 vss.n4609 vss.n4608 9.3005
R8783 vss.n4607 vss.n1049 9.3005
R8784 vss.n4606 vss.n4605 9.3005
R8785 vss.n4604 vss.n1061 9.3005
R8786 vss.n4603 vss.n4602 9.3005
R8787 vss.n4601 vss.n1073 9.3005
R8788 vss.n4600 vss.n4599 9.3005
R8789 vss.n4598 vss.n1085 9.3005
R8790 vss.n4597 vss.n4596 9.3005
R8791 vss.n4595 vss.n1097 9.3005
R8792 vss.n4594 vss.n4593 9.3005
R8793 vss.n4592 vss.n1109 9.3005
R8794 vss.n4591 vss.n4590 9.3005
R8795 vss.n5581 vss.n5580 9.3005
R8796 vss.n5584 vss.n265 9.3005
R8797 vss.n5588 vss.n5587 9.3005
R8798 vss.n5591 vss.n5590 9.3005
R8799 vss.n5589 vss.n260 9.3005
R8800 vss.n5595 vss.n257 9.3005
R8801 vss.n5599 vss.n5598 9.3005
R8802 vss.n5601 vss.n5600 9.3005
R8803 vss.n5604 vss.n251 9.3005
R8804 vss.n5608 vss.n5607 9.3005
R8805 vss.n5610 vss.n5609 9.3005
R8806 vss.n5614 vss.n248 9.3005
R8807 vss.n247 vss.n243 9.3005
R8808 vss.n5618 vss.n226 9.3005
R8809 vss.n5911 vss.n5910 9.3005
R8810 vss.n230 vss.n227 9.3005
R8811 vss.n5906 vss.n5905 9.3005
R8812 vss.n5904 vss.n5903 9.3005
R8813 vss.n239 vss.n237 9.3005
R8814 vss.n5898 vss.n5630 9.3005
R8815 vss.n5895 vss.n5894 9.3005
R8816 vss.n5893 vss.n5892 9.3005
R8817 vss.n5637 vss.n5635 9.3005
R8818 vss.n5886 vss.n5645 9.3005
R8819 vss.n5883 vss.n5882 9.3005
R8820 vss.n5881 vss.n5649 9.3005
R8821 vss.n5880 vss.n5879 9.3005
R8822 vss.n5876 vss.n5650 9.3005
R8823 vss.n5666 vss.n5657 9.3005
R8824 vss.n5871 vss.n5667 9.3005
R8825 vss.n5868 vss.n5867 9.3005
R8826 vss.n5866 vss.n5865 9.3005
R8827 vss.n5673 vss.n5671 9.3005
R8828 vss.n5860 vss.n5681 9.3005
R8829 vss.n5857 vss.n5856 9.3005
R8830 vss.n5855 vss.n5685 9.3005
R8831 vss.n5854 vss.n5853 9.3005
R8832 vss.n5850 vss.n5686 9.3005
R8833 vss.n5703 vss.n5693 9.3005
R8834 vss.n5845 vss.n5704 9.3005
R8835 vss.n5842 vss.n5841 9.3005
R8836 vss.n5840 vss.n5839 9.3005
R8837 vss.n5719 vss.n5710 9.3005
R8838 vss.n5834 vss.n5720 9.3005
R8839 vss.n5831 vss.n5830 9.3005
R8840 vss.n5829 vss.n5724 9.3005
R8841 vss.n5828 vss.n5827 9.3005
R8842 vss.n5824 vss.n5725 9.3005
R8843 vss.n5742 vss.n5732 9.3005
R8844 vss.n5819 vss.n5743 9.3005
R8845 vss.n5816 vss.n5815 9.3005
R8846 vss.n5814 vss.n5813 9.3005
R8847 vss.n5749 vss.n5747 9.3005
R8848 vss.n5808 vss.n5757 9.3005
R8849 vss.n5805 vss.n5804 9.3005
R8850 vss.n5802 vss.n218 9.3005
R8851 vss.n5581 vss.n267 9.3005
R8852 vss.n5585 vss.n5584 9.3005
R8853 vss.n5587 vss.n5586 9.3005
R8854 vss.n5591 vss.n263 9.3005
R8855 vss.n260 vss.n259 9.3005
R8856 vss.n5596 vss.n5595 9.3005
R8857 vss.n5598 vss.n5597 9.3005
R8858 vss.n5601 vss.n253 9.3005
R8859 vss.n5605 vss.n5604 9.3005
R8860 vss.n5607 vss.n5606 9.3005
R8861 vss.n5610 vss.n244 9.3005
R8862 vss.n5615 vss.n5614 9.3005
R8863 vss.n5616 vss.n243 9.3005
R8864 vss.n5618 vss.n5617 9.3005
R8865 vss.n5910 vss.n229 9.3005
R8866 vss.n234 vss.n230 9.3005
R8867 vss.n5906 vss.n235 9.3005
R8868 vss.n5903 vss.n238 9.3005
R8869 vss.n5627 vss.n239 9.3005
R8870 vss.n5898 vss.n5628 9.3005
R8871 vss.n5895 vss.n5633 9.3005
R8872 vss.n5892 vss.n5636 9.3005
R8873 vss.n5642 vss.n5637 9.3005
R8874 vss.n5886 vss.n5643 9.3005
R8875 vss.n5883 vss.n5648 9.3005
R8876 vss.n5652 vss.n5649 9.3005
R8877 vss.n5879 vss.n5653 9.3005
R8878 vss.n5876 vss.n5656 9.3005
R8879 vss.n5662 vss.n5657 9.3005
R8880 vss.n5871 vss.n5663 9.3005
R8881 vss.n5868 vss.n5669 9.3005
R8882 vss.n5865 vss.n5672 9.3005
R8883 vss.n5678 vss.n5673 9.3005
R8884 vss.n5860 vss.n5679 9.3005
R8885 vss.n5857 vss.n5684 9.3005
R8886 vss.n5688 vss.n5685 9.3005
R8887 vss.n5853 vss.n5689 9.3005
R8888 vss.n5850 vss.n5692 9.3005
R8889 vss.n5700 vss.n5693 9.3005
R8890 vss.n5845 vss.n5701 9.3005
R8891 vss.n5842 vss.n5706 9.3005
R8892 vss.n5839 vss.n5709 9.3005
R8893 vss.n5716 vss.n5710 9.3005
R8894 vss.n5834 vss.n5717 9.3005
R8895 vss.n5831 vss.n5723 9.3005
R8896 vss.n5727 vss.n5724 9.3005
R8897 vss.n5827 vss.n5728 9.3005
R8898 vss.n5824 vss.n5731 9.3005
R8899 vss.n5739 vss.n5732 9.3005
R8900 vss.n5819 vss.n5740 9.3005
R8901 vss.n5816 vss.n5745 9.3005
R8902 vss.n5813 vss.n5748 9.3005
R8903 vss.n5754 vss.n5749 9.3005
R8904 vss.n5808 vss.n5755 9.3005
R8905 vss.n5582 vss.n5581 9.3005
R8906 vss.n5584 vss.n5583 9.3005
R8907 vss.n5587 vss.n261 9.3005
R8908 vss.n5592 vss.n5591 9.3005
R8909 vss.n5593 vss.n260 9.3005
R8910 vss.n5595 vss.n5594 9.3005
R8911 vss.n5598 vss.n255 9.3005
R8912 vss.n5602 vss.n5601 9.3005
R8913 vss.n5604 vss.n5603 9.3005
R8914 vss.n5607 vss.n249 9.3005
R8915 vss.n5611 vss.n5610 9.3005
R8916 vss.n5614 vss.n5613 9.3005
R8917 vss.n5612 vss.n243 9.3005
R8918 vss.n5618 vss.n231 9.3005
R8919 vss.n5910 vss.n5909 9.3005
R8920 vss.n5908 vss.n230 9.3005
R8921 vss.n5907 vss.n5906 9.3005
R8922 vss.n5903 vss.n232 9.3005
R8923 vss.n5631 vss.n239 9.3005
R8924 vss.n5898 vss.n5897 9.3005
R8925 vss.n5896 vss.n5895 9.3005
R8926 vss.n5892 vss.n5632 9.3005
R8927 vss.n5646 vss.n5637 9.3005
R8928 vss.n5886 vss.n5885 9.3005
R8929 vss.n5884 vss.n5883 9.3005
R8930 vss.n5649 vss.n5647 9.3005
R8931 vss.n5879 vss.n5878 9.3005
R8932 vss.n5877 vss.n5876 9.3005
R8933 vss.n5657 vss.n5655 9.3005
R8934 vss.n5871 vss.n5870 9.3005
R8935 vss.n5869 vss.n5868 9.3005
R8936 vss.n5865 vss.n5668 9.3005
R8937 vss.n5682 vss.n5673 9.3005
R8938 vss.n5860 vss.n5859 9.3005
R8939 vss.n5858 vss.n5857 9.3005
R8940 vss.n5685 vss.n5683 9.3005
R8941 vss.n5853 vss.n5852 9.3005
R8942 vss.n5851 vss.n5850 9.3005
R8943 vss.n5693 vss.n5691 9.3005
R8944 vss.n5845 vss.n5844 9.3005
R8945 vss.n5843 vss.n5842 9.3005
R8946 vss.n5839 vss.n5705 9.3005
R8947 vss.n5721 vss.n5710 9.3005
R8948 vss.n5834 vss.n5833 9.3005
R8949 vss.n5832 vss.n5831 9.3005
R8950 vss.n5724 vss.n5722 9.3005
R8951 vss.n5827 vss.n5826 9.3005
R8952 vss.n5825 vss.n5824 9.3005
R8953 vss.n5732 vss.n5730 9.3005
R8954 vss.n5819 vss.n5818 9.3005
R8955 vss.n5817 vss.n5816 9.3005
R8956 vss.n5813 vss.n5744 9.3005
R8957 vss.n5758 vss.n5749 9.3005
R8958 vss.n5808 vss.n5807 9.3005
R8959 vss.n5806 vss.n5805 9.3005
R8960 vss.n5573 vss.n272 9.3005
R8961 vss.n5577 vss.n5576 9.3005
R8962 vss.n5573 vss.n5572 9.3005
R8963 vss.n5576 vss.n274 9.3005
R8964 vss.n5574 vss.n5573 9.3005
R8965 vss.n5576 vss.n5575 9.3005
R8966 vss.n2220 vss.n2219 9.3005
R8967 vss.n2222 vss.n2221 9.3005
R8968 vss.n4220 vss.n1309 9.3005
R8969 vss.n4222 vss.n4221 9.3005
R8970 vss.n2976 vss.n2975 9.3005
R8971 vss.n2972 vss.n2969 9.3005
R8972 vss.n2406 vss.n2405 9.3005
R8973 vss.n2404 vss.n2397 9.3005
R8974 vss.n5539 vss.n5538 9.3005
R8975 vss.n5538 vss.n296 9.3005
R8976 vss.n2248 vss.n2240 9.3005
R8977 vss.n2289 vss.n2241 9.3005
R8978 vss.n2243 vss.n2242 9.3005
R8979 vss.n2306 vss.n2209 9.3005
R8980 vss.n2313 vss.n2312 9.3005
R8981 vss.n2214 vss.n1298 9.3005
R8982 vss.n2213 vss.n1299 9.3005
R8983 vss.n2210 vss.n1300 9.3005
R8984 vss.n4218 vss.n1311 9.3005
R8985 vss.n2197 vss.n1312 9.3005
R8986 vss.n2198 vss.n1315 9.3005
R8987 vss.n4209 vss.n1317 9.3005
R8988 vss.n2981 vss.n2978 9.3005
R8989 vss.n2986 vss.n2984 9.3005
R8990 vss.n2983 vss.n2335 9.3005
R8991 vss.n3010 vss.n2336 9.3005
R8992 vss.n2408 vss.n2392 9.3005
R8993 vss.n2423 vss.n2393 9.3005
R8994 vss.n2426 vss.n2424 9.3005
R8995 vss.n2387 vss.n2380 9.3005
R8996 vss.n2442 vss.n2381 9.3005
R8997 vss.n2450 vss.n2376 9.3005
R8998 vss.n2245 vss.n2240 9.3005
R8999 vss.n2289 vss.n2288 9.3005
R9000 vss.n2243 vss.n2229 9.3005
R9001 vss.n2307 vss.n2306 9.3005
R9002 vss.n2313 vss.n1297 9.3005
R9003 vss.n4231 vss.n1298 9.3005
R9004 vss.n4230 vss.n1299 9.3005
R9005 vss.n4229 vss.n1300 9.3005
R9006 vss.n4218 vss.n1301 9.3005
R9007 vss.n3022 vss.n1312 9.3005
R9008 vss.n1319 vss.n1315 9.3005
R9009 vss.n4209 vss.n4208 9.3005
R9010 vss.n2978 vss.n1320 9.3005
R9011 vss.n2987 vss.n2986 9.3005
R9012 vss.n2338 vss.n2335 9.3005
R9013 vss.n3010 vss.n3009 9.3005
R9014 vss.n2408 vss.n2339 9.3005
R9015 vss.n2393 vss.n2390 9.3005
R9016 vss.n2427 vss.n2426 9.3005
R9017 vss.n2428 vss.n2380 9.3005
R9018 vss.n2442 vss.n2374 9.3005
R9019 vss.n2451 vss.n2450 9.3005
R9020 vss.n2293 vss.n2237 9.3005
R9021 vss.n2295 vss.n2294 9.3005
R9022 vss.n2297 vss.n2296 9.3005
R9023 vss.n2440 vss.n2378 9.3005
R9024 vss.n2439 vss.n2438 9.3005
R9025 vss.n2244 vss.n2231 9.3005
R9026 vss.n2303 vss.n2230 9.3005
R9027 vss.n2317 vss.n2316 9.3005
R9028 vss.n2320 vss.n2319 9.3005
R9029 vss.n4213 vss.n4212 9.3005
R9030 vss.n2985 vss.n2333 9.3005
R9031 vss.n3012 vss.n3011 9.3005
R9032 vss.n2411 vss.n2391 9.3005
R9033 vss.n2425 vss.n2379 9.3005
R9034 vss.n2449 vss.n2448 9.3005
R9035 vss.n2377 vss.n300 9.3005
R9036 vss.n2291 vss.n2290 9.3005
R9037 vss.n2315 vss.n2314 9.3005
R9038 vss.n2305 vss.n2304 9.3005
R9039 vss.n4215 vss.n4214 9.3005
R9040 vss.n4217 vss.n4216 9.3005
R9041 vss.n2318 vss.n1310 9.3005
R9042 vss.n2410 vss.n2409 9.3005
R9043 vss.n2337 vss.n2334 9.3005
R9044 vss.n2446 vss.n2375 9.3005
R9045 vss.n2444 vss.n2443 9.3005
R9046 vss.n5537 vss.n5536 9.3005
R9047 vss.n2973 vss.n2968 9.3005
R9048 vss.n1318 vss.n1316 9.3005
R9049 vss.n4211 vss.n4210 9.3005
R9050 vss.n5534 vss.n5533 9.3005
R9051 vss.n5532 vss.n302 9.3005
R9052 vss.n4381 vss.n4380 9.3005
R9053 vss.n4377 vss.n4376 9.3005
R9054 vss.n4373 vss.n4372 9.3005
R9055 vss.n4371 vss.n4370 9.3005
R9056 vss.n4368 vss.n4365 9.3005
R9057 vss.n5541 vss.n5540 9.3005
R9058 vss.n5543 vss.n5542 9.3005
R9059 vss.n5535 vss.n301 9.3005
R9060 vss.n4584 vss.n753 9.3005
R9061 vss.n4586 vss.n4585 9.3005
R9062 vss.n5348 vss.n5343 9.3005
R9063 vss.n5342 vss.n5339 9.3005
R9064 vss.n5341 vss.n5338 9.3005
R9065 vss.n5340 vss.n5337 9.3005
R9066 vss.n5336 vss.n1004 9.3005
R9067 vss.n5335 vss.n894 9.3005
R9068 vss.n868 vss.n858 9.3005
R9069 vss.n867 vss.n857 9.3005
R9070 vss.n856 vss.n848 9.3005
R9071 vss.n855 vss.n853 9.3005
R9072 vss.n836 vss.n826 9.3005
R9073 vss.n835 vss.n825 9.3005
R9074 vss.n824 vss.n816 9.3005
R9075 vss.n823 vss.n821 9.3005
R9076 vss.n801 vss.n791 9.3005
R9077 vss.n800 vss.n790 9.3005
R9078 vss.n789 vss.n783 9.3005
R9079 vss.n4579 vss.n4577 9.3005
R9080 vss.n4580 vss.n767 9.3005
R9081 vss.n4583 vss.n4581 9.3005
R9082 vss.n4583 vss.n4576 9.3005
R9083 vss.n4580 vss.n772 9.3005
R9084 vss.n4579 vss.n788 9.3005
R9085 vss.n5383 vss.n789 9.3005
R9086 vss.n5382 vss.n790 9.3005
R9087 vss.n5381 vss.n791 9.3005
R9088 vss.n823 vss.n792 9.3005
R9089 vss.n5373 vss.n824 9.3005
R9090 vss.n5372 vss.n825 9.3005
R9091 vss.n5371 vss.n826 9.3005
R9092 vss.n855 vss.n827 9.3005
R9093 vss.n5363 vss.n856 9.3005
R9094 vss.n5362 vss.n857 9.3005
R9095 vss.n5361 vss.n858 9.3005
R9096 vss.n5335 vss.n859 9.3005
R9097 vss.n5353 vss.n5336 9.3005
R9098 vss.n5352 vss.n5337 9.3005
R9099 vss.n5351 vss.n5338 9.3005
R9100 vss.n5350 vss.n5339 9.3005
R9101 vss.n5349 vss.n5348 9.3005
R9102 vss.n5348 vss.n5347 9.3005
R9103 vss.n5346 vss.n5339 9.3005
R9104 vss.n5345 vss.n5338 9.3005
R9105 vss.n5344 vss.n5337 9.3005
R9106 vss.n5336 vss.n1003 9.3005
R9107 vss.n5335 vss.n892 9.3005
R9108 vss.n865 vss.n858 9.3005
R9109 vss.n864 vss.n857 9.3005
R9110 vss.n856 vss.n846 9.3005
R9111 vss.n855 vss.n854 9.3005
R9112 vss.n833 vss.n826 9.3005
R9113 vss.n832 vss.n825 9.3005
R9114 vss.n824 vss.n813 9.3005
R9115 vss.n823 vss.n822 9.3005
R9116 vss.n798 vss.n791 9.3005
R9117 vss.n797 vss.n790 9.3005
R9118 vss.n789 vss.n781 9.3005
R9119 vss.n4579 vss.n4578 9.3005
R9120 vss.n4580 vss.n765 9.3005
R9121 vss.n4583 vss.n4582 9.3005
R9122 vss.n4584 vss.n755 9.3005
R9123 vss.n4585 vss.n4266 9.3005
R9124 vss.n4267 vss.n734 9.3005
R9125 vss.n4572 vss.n4571 9.3005
R9126 vss.n4570 vss.n720 9.3005
R9127 vss.n4270 vss.n4269 9.3005
R9128 vss.n4566 vss.n706 9.3005
R9129 vss.n4564 vss.n4563 9.3005
R9130 vss.n4272 vss.n692 9.3005
R9131 vss.n4556 vss.n4555 9.3005
R9132 vss.n4553 vss.n678 9.3005
R9133 vss.n4275 vss.n4274 9.3005
R9134 vss.n4546 vss.n664 9.3005
R9135 vss.n4544 vss.n4543 9.3005
R9136 vss.n4277 vss.n650 9.3005
R9137 vss.n4536 vss.n4535 9.3005
R9138 vss.n4533 vss.n636 9.3005
R9139 vss.n4280 vss.n4279 9.3005
R9140 vss.n4526 vss.n622 9.3005
R9141 vss.n4524 vss.n4523 9.3005
R9142 vss.n4282 vss.n608 9.3005
R9143 vss.n4516 vss.n4515 9.3005
R9144 vss.n4513 vss.n594 9.3005
R9145 vss.n4285 vss.n4284 9.3005
R9146 vss.n4506 vss.n580 9.3005
R9147 vss.n4504 vss.n4503 9.3005
R9148 vss.n4288 vss.n566 9.3005
R9149 vss.n4498 vss.n4497 9.3005
R9150 vss.n4495 vss.n552 9.3005
R9151 vss.n4494 vss.n4493 9.3005
R9152 vss.n4485 vss.n538 9.3005
R9153 vss.n4487 vss.n4486 9.3005
R9154 vss.n4484 vss.n524 9.3005
R9155 vss.n4482 vss.n4481 9.3005
R9156 vss.n4292 vss.n510 9.3005
R9157 vss.n4474 vss.n4473 9.3005
R9158 vss.n4471 vss.n496 9.3005
R9159 vss.n4295 vss.n4294 9.3005
R9160 vss.n4464 vss.n482 9.3005
R9161 vss.n4462 vss.n4461 9.3005
R9162 vss.n4297 vss.n468 9.3005
R9163 vss.n4454 vss.n4453 9.3005
R9164 vss.n4451 vss.n454 9.3005
R9165 vss.n4300 vss.n4299 9.3005
R9166 vss.n4444 vss.n440 9.3005
R9167 vss.n4442 vss.n4441 9.3005
R9168 vss.n4302 vss.n426 9.3005
R9169 vss.n4434 vss.n4433 9.3005
R9170 vss.n4431 vss.n412 9.3005
R9171 vss.n4305 vss.n4304 9.3005
R9172 vss.n4424 vss.n398 9.3005
R9173 vss.n4309 vss.n4308 9.3005
R9174 vss.n4419 vss.n384 9.3005
R9175 vss.n4417 vss.n4416 9.3005
R9176 vss.n4311 vss.n370 9.3005
R9177 vss.n4411 vss.n4410 9.3005
R9178 vss.n4314 vss.n356 9.3005
R9179 vss.n4404 vss.n4403 9.3005
R9180 vss.n4402 vss.n342 9.3005
R9181 vss.n4317 vss.n4316 9.3005
R9182 vss.n4396 vss.n328 9.3005
R9183 vss.n4320 vss.n4319 9.3005
R9184 vss.n4390 vss.n314 9.3005
R9185 vss.n4388 vss.n4387 9.3005
R9186 vss.n4323 vss.n1013 9.3005
R9187 vss.n4357 vss.n4356 9.3005
R9188 vss.n4354 vss.n1026 9.3005
R9189 vss.n4328 vss.n4327 9.3005
R9190 vss.n4350 vss.n1038 9.3005
R9191 vss.n4349 vss.n4348 9.3005
R9192 vss.n4347 vss.n1050 9.3005
R9193 vss.n4346 vss.n4345 9.3005
R9194 vss.n4344 vss.n1062 9.3005
R9195 vss.n4343 vss.n4342 9.3005
R9196 vss.n4341 vss.n1074 9.3005
R9197 vss.n4340 vss.n4339 9.3005
R9198 vss.n4338 vss.n1086 9.3005
R9199 vss.n4337 vss.n4336 9.3005
R9200 vss.n4335 vss.n1098 9.3005
R9201 vss.n4334 vss.n4333 9.3005
R9202 vss.n4332 vss.n1110 9.3005
R9203 vss.n4331 vss.n4330 9.3005
R9204 vss.n6011 vss.n132 9.3005
R9205 vss.n5983 vss.n130 9.3005
R9206 vss.n5987 vss.n5984 9.3005
R9207 vss.n5990 vss.n5979 9.3005
R9208 vss.n5992 vss.n5977 9.3005
R9209 vss.n5995 vss.n5973 9.3005
R9210 vss.n5998 vss.n153 9.3005
R9211 vss.n6001 vss.n6000 9.3005
R9212 vss.n5966 vss.n152 9.3005
R9213 vss.n5963 vss.n161 9.3005
R9214 vss.n5960 vss.n5959 9.3005
R9215 vss.n5958 vss.n164 9.3005
R9216 vss.n5954 vss.n166 9.3005
R9217 vss.n5951 vss.n177 9.3005
R9218 vss.n5948 vss.n5947 9.3005
R9219 vss.n5946 vss.n5945 9.3005
R9220 vss.n5942 vss.n182 9.3005
R9221 vss.n5939 vss.n5938 9.3005
R9222 vss.n5937 vss.n5936 9.3005
R9223 vss.n5933 vss.n193 9.3005
R9224 vss.n5930 vss.n5929 9.3005
R9225 vss.n5928 vss.n5927 9.3005
R9226 vss.n5924 vss.n203 9.3005
R9227 vss.n213 vss.n208 9.3005
R9228 vss.n2769 vss.n2768 9.3005
R9229 vss.n2771 vss.n2770 9.3005
R9230 vss.n2774 vss.n2752 9.3005
R9231 vss.n2778 vss.n2777 9.3005
R9232 vss.n2780 vss.n2779 9.3005
R9233 vss.n2783 vss.n2739 9.3005
R9234 vss.n2787 vss.n2786 9.3005
R9235 vss.n2789 vss.n2788 9.3005
R9236 vss.n2792 vss.n2731 9.3005
R9237 vss.n2795 vss.n2723 9.3005
R9238 vss.n2796 vss.n2721 9.3005
R9239 vss.n2799 vss.n2709 9.3005
R9240 vss.n2803 vss.n2802 9.3005
R9241 vss.n2805 vss.n2804 9.3005
R9242 vss.n2808 vss.n2693 9.3005
R9243 vss.n2812 vss.n2811 9.3005
R9244 vss.n2814 vss.n2813 9.3005
R9245 vss.n2817 vss.n2685 9.3005
R9246 vss.n2820 vss.n2677 9.3005
R9247 vss.n2822 vss.n2675 9.3005
R9248 vss.n2825 vss.n2671 9.3005
R9249 vss.n2670 vss.n65 9.3005
R9250 vss.n2829 vss.n2660 9.3005
R9251 vss.n2832 vss.n2652 9.3005
R9252 vss.n2834 vss.n2650 9.3005
R9253 vss.n2837 vss.n2638 9.3005
R9254 vss.n2841 vss.n2840 9.3005
R9255 vss.n2843 vss.n2842 9.3005
R9256 vss.n2846 vss.n2625 9.3005
R9257 vss.n2850 vss.n2849 9.3005
R9258 vss.n2852 vss.n2851 9.3005
R9259 vss.n2855 vss.n2617 9.3005
R9260 vss.n2616 vss.n2606 9.3005
R9261 vss.n2859 vss.n2598 9.3005
R9262 vss.n2863 vss.n2862 9.3005
R9263 vss.n2865 vss.n2864 9.3005
R9264 vss.n2868 vss.n2585 9.3005
R9265 vss.n2872 vss.n2871 9.3005
R9266 vss.n2874 vss.n2873 9.3005
R9267 vss.n2877 vss.n2577 9.3005
R9268 vss.n2880 vss.n2571 9.3005
R9269 vss.n2882 vss.n2569 9.3005
R9270 vss.n2885 vss.n2562 9.3005
R9271 vss.n2888 vss.n2554 9.3005
R9272 vss.n2889 vss.n2552 9.3005
R9273 vss.n2892 vss.n2539 9.3005
R9274 vss.n2896 vss.n2895 9.3005
R9275 vss.n2898 vss.n2897 9.3005
R9276 vss.n2901 vss.n2534 9.3005
R9277 vss.n2904 vss.n2527 9.3005
R9278 vss.n2906 vss.n2525 9.3005
R9279 vss.n2909 vss.n2514 9.3005
R9280 vss.n2913 vss.n2912 9.3005
R9281 vss.n2915 vss.n2914 9.3005
R9282 vss.n2918 vss.n2505 9.3005
R9283 vss.n2504 vss.n26 9.3005
R9284 vss.n2922 vss.n2488 9.3005
R9285 vss.n2926 vss.n2925 9.3005
R9286 vss.n2928 vss.n2927 9.3005
R9287 vss.n2931 vss.n2475 9.3005
R9288 vss.n2935 vss.n2934 9.3005
R9289 vss.n2937 vss.n2936 9.3005
R9290 vss.n2940 vss.n2463 9.3005
R9291 vss.n2944 vss.n2943 9.3005
R9292 vss.n2946 vss.n2945 9.3005
R9293 vss.n2949 vss.n2370 9.3005
R9294 vss.n2369 vss.n2362 9.3005
R9295 vss.n2953 vss.n2361 9.3005
R9296 vss.n2955 vss.n2359 9.3005
R9297 vss.n2958 vss.n2350 9.3005
R9298 vss.n2962 vss.n2961 9.3005
R9299 vss.n3004 vss.n3003 9.3005
R9300 vss.n3001 vss.n2349 9.3005
R9301 vss.n2998 vss.n2993 9.3005
R9302 vss.n2995 vss.n1332 9.3005
R9303 vss.n4202 vss.n4201 9.3005
R9304 vss.n4199 vss.n1331 9.3005
R9305 vss.n4196 vss.n1340 9.3005
R9306 vss.n4192 vss.n1338 9.3005
R9307 vss.n4191 vss.n4190 9.3005
R9308 vss.n4187 vss.n1345 9.3005
R9309 vss.n4184 vss.n4183 9.3005
R9310 vss.n4182 vss.n4181 9.3005
R9311 vss.n4178 vss.n1357 9.3005
R9312 vss.n4175 vss.n4174 9.3005
R9313 vss.n4173 vss.n4172 9.3005
R9314 vss.n4169 vss.n1368 9.3005
R9315 vss.n4166 vss.n4165 9.3005
R9316 vss.n4164 vss.n4163 9.3005
R9317 vss.n4160 vss.n1380 9.3005
R9318 vss.n4156 vss.n1386 9.3005
R9319 vss.n4155 vss.n4154 9.3005
R9320 vss.n4151 vss.n1392 9.3005
R9321 vss.n4148 vss.n4147 9.3005
R9322 vss.n4146 vss.n4145 9.3005
R9323 vss.n4142 vss.n1404 9.3005
R9324 vss.n4139 vss.n4138 9.3005
R9325 vss.n4137 vss.n4136 9.3005
R9326 vss.n4133 vss.n1416 9.3005
R9327 vss.n4130 vss.n4129 9.3005
R9328 vss.n4128 vss.n4127 9.3005
R9329 vss.n1430 vss.n1428 9.3005
R9330 vss.n4121 vss.n1448 9.3005
R9331 vss.n4118 vss.n1453 9.3005
R9332 vss.n4115 vss.n4114 9.3005
R9333 vss.n4113 vss.n4112 9.3005
R9334 vss.n4109 vss.n1458 9.3005
R9335 vss.n4106 vss.n4105 9.3005
R9336 vss.n4104 vss.n4103 9.3005
R9337 vss.n4100 vss.n1470 9.3005
R9338 vss.n4097 vss.n4096 9.3005
R9339 vss.n4095 vss.n4094 9.3005
R9340 vss.n1484 vss.n1482 9.3005
R9341 vss.n4088 vss.n1502 9.3005
R9342 vss.n4085 vss.n1507 9.3005
R9343 vss.n4082 vss.n4081 9.3005
R9344 vss.n4080 vss.n4079 9.3005
R9345 vss.n4076 vss.n1512 9.3005
R9346 vss.n4073 vss.n4072 9.3005
R9347 vss.n4071 vss.n4070 9.3005
R9348 vss.n4067 vss.n1524 9.3005
R9349 vss.n4064 vss.n4063 9.3005
R9350 vss.n4062 vss.n4061 9.3005
R9351 vss.n4058 vss.n1536 9.3005
R9352 vss.n4054 vss.n1542 9.3005
R9353 vss.n4053 vss.n4052 9.3005
R9354 vss.n4049 vss.n1559 9.3005
R9355 vss.n4046 vss.n4045 9.3005
R9356 vss.n4044 vss.n4043 9.3005
R9357 vss.n4040 vss.n1571 9.3005
R9358 vss.n4037 vss.n4036 9.3005
R9359 vss.n4035 vss.n4034 9.3005
R9360 vss.n4031 vss.n1583 9.3005
R9361 vss.n4028 vss.n4027 9.3005
R9362 vss.n4026 vss.n4025 9.3005
R9363 vss.n1597 vss.n1595 9.3005
R9364 vss.n4019 vss.n1615 9.3005
R9365 vss.n4016 vss.n1620 9.3005
R9366 vss.n4013 vss.n4012 9.3005
R9367 vss.n4011 vss.n4010 9.3005
R9368 vss.n4007 vss.n1625 9.3005
R9369 vss.n4004 vss.n4003 9.3005
R9370 vss.n4002 vss.n4001 9.3005
R9371 vss.n3998 vss.n1637 9.3005
R9372 vss.n3995 vss.n3994 9.3005
R9373 vss.n3993 vss.n3992 9.3005
R9374 vss.n1651 vss.n1649 9.3005
R9375 vss.n3986 vss.n1669 9.3005
R9376 vss.n3983 vss.n1674 9.3005
R9377 vss.n3980 vss.n3979 9.3005
R9378 vss.n3978 vss.n3977 9.3005
R9379 vss.n3974 vss.n1679 9.3005
R9380 vss.n3971 vss.n3970 9.3005
R9381 vss.n3969 vss.n3968 9.3005
R9382 vss.n3965 vss.n1691 9.3005
R9383 vss.n3962 vss.n3961 9.3005
R9384 vss.n3960 vss.n3959 9.3005
R9385 vss.n3956 vss.n1703 9.3005
R9386 vss.n3952 vss.n1709 9.3005
R9387 vss.n3951 vss.n3950 9.3005
R9388 vss.n3947 vss.n1726 9.3005
R9389 vss.n3944 vss.n3943 9.3005
R9390 vss.n3942 vss.n3941 9.3005
R9391 vss.n3938 vss.n1738 9.3005
R9392 vss.n3935 vss.n3934 9.3005
R9393 vss.n3933 vss.n3932 9.3005
R9394 vss.n3929 vss.n1750 9.3005
R9395 vss.n3926 vss.n3925 9.3005
R9396 vss.n3924 vss.n3923 9.3005
R9397 vss.n1764 vss.n1762 9.3005
R9398 vss.n3917 vss.n1772 9.3005
R9399 vss.n3914 vss.n1777 9.3005
R9400 vss.n3911 vss.n3910 9.3005
R9401 vss.n3909 vss.n3908 9.3005
R9402 vss.n3905 vss.n1782 9.3005
R9403 vss.n3902 vss.n3901 9.3005
R9404 vss.n3900 vss.n3899 9.3005
R9405 vss.n3896 vss.n1794 9.3005
R9406 vss.n3893 vss.n3892 9.3005
R9407 vss.n3891 vss.n3890 9.3005
R9408 vss.n3887 vss.n1806 9.3005
R9409 vss.n3883 vss.n1812 9.3005
R9410 vss.n3882 vss.n3881 9.3005
R9411 vss.n3878 vss.n1829 9.3005
R9412 vss.n3875 vss.n3874 9.3005
R9413 vss.n3873 vss.n3872 9.3005
R9414 vss.n3869 vss.n1841 9.3005
R9415 vss.n3866 vss.n3865 9.3005
R9416 vss.n3864 vss.n3863 9.3005
R9417 vss.n3860 vss.n1853 9.3005
R9418 vss.n3857 vss.n3856 9.3005
R9419 vss.n3855 vss.n3854 9.3005
R9420 vss.n1867 vss.n1865 9.3005
R9421 vss.n3848 vss.n1885 9.3005
R9422 vss.n3845 vss.n1890 9.3005
R9423 vss.n3842 vss.n3841 9.3005
R9424 vss.n3840 vss.n3839 9.3005
R9425 vss.n3836 vss.n1895 9.3005
R9426 vss.n3833 vss.n3832 9.3005
R9427 vss.n3831 vss.n3830 9.3005
R9428 vss.n3827 vss.n1907 9.3005
R9429 vss.n3824 vss.n3823 9.3005
R9430 vss.n3822 vss.n3821 9.3005
R9431 vss.n1921 vss.n1919 9.3005
R9432 vss.n3815 vss.n1939 9.3005
R9433 vss.n3812 vss.n1944 9.3005
R9434 vss.n3809 vss.n3808 9.3005
R9435 vss.n3807 vss.n3806 9.3005
R9436 vss.n3803 vss.n1949 9.3005
R9437 vss.n3800 vss.n3799 9.3005
R9438 vss.n3798 vss.n3797 9.3005
R9439 vss.n3794 vss.n1961 9.3005
R9440 vss.n3791 vss.n3790 9.3005
R9441 vss.n3789 vss.n3788 9.3005
R9442 vss.n3785 vss.n1973 9.3005
R9443 vss.n3781 vss.n1979 9.3005
R9444 vss.n3780 vss.n3779 9.3005
R9445 vss.n3776 vss.n1996 9.3005
R9446 vss.n3773 vss.n3772 9.3005
R9447 vss.n3771 vss.n3770 9.3005
R9448 vss.n3767 vss.n2008 9.3005
R9449 vss.n3764 vss.n3763 9.3005
R9450 vss.n3762 vss.n3761 9.3005
R9451 vss.n3758 vss.n2020 9.3005
R9452 vss.n3755 vss.n3754 9.3005
R9453 vss.n3753 vss.n3752 9.3005
R9454 vss.n2034 vss.n2032 9.3005
R9455 vss.n3746 vss.n2052 9.3005
R9456 vss.n3743 vss.n2057 9.3005
R9457 vss.n3740 vss.n3739 9.3005
R9458 vss.n3738 vss.n3737 9.3005
R9459 vss.n3734 vss.n2062 9.3005
R9460 vss.n3731 vss.n3730 9.3005
R9461 vss.n3729 vss.n3728 9.3005
R9462 vss.n3725 vss.n2074 9.3005
R9463 vss.n3722 vss.n3721 9.3005
R9464 vss.n3720 vss.n3719 9.3005
R9465 vss.n2088 vss.n2086 9.3005
R9466 vss.n3713 vss.n2106 9.3005
R9467 vss.n3710 vss.n2111 9.3005
R9468 vss.n3707 vss.n3706 9.3005
R9469 vss.n3705 vss.n3704 9.3005
R9470 vss.n3701 vss.n2116 9.3005
R9471 vss.n3698 vss.n3697 9.3005
R9472 vss.n3696 vss.n3695 9.3005
R9473 vss.n3692 vss.n2128 9.3005
R9474 vss.n3689 vss.n3688 9.3005
R9475 vss.n3687 vss.n3686 9.3005
R9476 vss.n3683 vss.n2140 9.3005
R9477 vss.n3679 vss.n2146 9.3005
R9478 vss.n3678 vss.n3677 9.3005
R9479 vss.n3674 vss.n2152 9.3005
R9480 vss.n3671 vss.n3670 9.3005
R9481 vss.n3669 vss.n3668 9.3005
R9482 vss.n3665 vss.n2164 9.3005
R9483 vss.n3662 vss.n3661 9.3005
R9484 vss.n3660 vss.n3659 9.3005
R9485 vss.n3656 vss.n2176 9.3005
R9486 vss.n3653 vss.n3652 9.3005
R9487 vss.n3651 vss.n3650 9.3005
R9488 vss.n2190 vss.n2188 9.3005
R9489 vss.n3607 vss.n3606 9.3005
R9490 vss.n3609 vss.n3608 9.3005
R9491 vss.n3613 vss.n3077 9.3005
R9492 vss.n3071 vss.n3070 9.3005
R9493 vss.n3618 vss.n3617 9.3005
R9494 vss.n3620 vss.n3619 9.3005
R9495 vss.n3623 vss.n3061 9.3005
R9496 vss.n3627 vss.n3626 9.3005
R9497 vss.n3629 vss.n3628 9.3005
R9498 vss.n3632 vss.n3052 9.3005
R9499 vss.n3636 vss.n3635 9.3005
R9500 vss.n3638 vss.n3637 9.3005
R9501 vss.n3641 vss.n3048 9.3005
R9502 vss.n3644 vss.n3044 9.3005
R9503 vss.n6011 vss.n133 9.3005
R9504 vss.n5985 vss.n130 9.3005
R9505 vss.n5987 vss.n5986 9.3005
R9506 vss.n5990 vss.n5975 9.3005
R9507 vss.n5993 vss.n5992 9.3005
R9508 vss.n5995 vss.n5994 9.3005
R9509 vss.n5998 vss.n5970 9.3005
R9510 vss.n6000 vss.n146 9.3005
R9511 vss.n5966 vss.n156 9.3005
R9512 vss.n5963 vss.n5962 9.3005
R9513 vss.n5961 vss.n5960 9.3005
R9514 vss.n164 vss.n162 9.3005
R9515 vss.n5954 vss.n173 9.3005
R9516 vss.n5951 vss.n5950 9.3005
R9517 vss.n5949 vss.n5948 9.3005
R9518 vss.n5945 vss.n178 9.3005
R9519 vss.n5942 vss.n5941 9.3005
R9520 vss.n5940 vss.n5939 9.3005
R9521 vss.n5936 vss.n189 9.3005
R9522 vss.n5933 vss.n5932 9.3005
R9523 vss.n5931 vss.n5930 9.3005
R9524 vss.n5927 vss.n199 9.3005
R9525 vss.n5924 vss.n5923 9.3005
R9526 vss.n5922 vss.n208 9.3005
R9527 vss.n2768 vss.n210 9.3005
R9528 vss.n2771 vss.n2758 9.3005
R9529 vss.n2775 vss.n2774 9.3005
R9530 vss.n2777 vss.n2776 9.3005
R9531 vss.n2780 vss.n2743 9.3005
R9532 vss.n2784 vss.n2783 9.3005
R9533 vss.n2786 vss.n2785 9.3005
R9534 vss.n2789 vss.n2729 9.3005
R9535 vss.n2793 vss.n2792 9.3005
R9536 vss.n2795 vss.n2794 9.3005
R9537 vss.n2796 vss.n2712 9.3005
R9538 vss.n2800 vss.n2799 9.3005
R9539 vss.n2802 vss.n2801 9.3005
R9540 vss.n2805 vss.n2700 9.3005
R9541 vss.n2809 vss.n2808 9.3005
R9542 vss.n2811 vss.n2810 9.3005
R9543 vss.n2814 vss.n2683 9.3005
R9544 vss.n2818 vss.n2817 9.3005
R9545 vss.n2820 vss.n2819 9.3005
R9546 vss.n2822 vss.n2667 9.3005
R9547 vss.n2826 vss.n2825 9.3005
R9548 vss.n2827 vss.n65 9.3005
R9549 vss.n2829 vss.n2828 9.3005
R9550 vss.n2832 vss.n2648 9.3005
R9551 vss.n2835 vss.n2834 9.3005
R9552 vss.n2837 vss.n2836 9.3005
R9553 vss.n2840 vss.n2635 9.3005
R9554 vss.n2844 vss.n2843 9.3005
R9555 vss.n2846 vss.n2845 9.3005
R9556 vss.n2849 vss.n2619 9.3005
R9557 vss.n2853 vss.n2852 9.3005
R9558 vss.n2855 vss.n2854 9.3005
R9559 vss.n2606 vss.n2604 9.3005
R9560 vss.n2860 vss.n2859 9.3005
R9561 vss.n2862 vss.n2861 9.3005
R9562 vss.n2865 vss.n2589 9.3005
R9563 vss.n2869 vss.n2868 9.3005
R9564 vss.n2871 vss.n2870 9.3005
R9565 vss.n2874 vss.n2575 9.3005
R9566 vss.n2878 vss.n2877 9.3005
R9567 vss.n2880 vss.n2879 9.3005
R9568 vss.n2882 vss.n2560 9.3005
R9569 vss.n2886 vss.n2885 9.3005
R9570 vss.n2888 vss.n2887 9.3005
R9571 vss.n2889 vss.n2547 9.3005
R9572 vss.n2893 vss.n2892 9.3005
R9573 vss.n2895 vss.n2894 9.3005
R9574 vss.n2898 vss.n2532 9.3005
R9575 vss.n2902 vss.n2901 9.3005
R9576 vss.n2904 vss.n2903 9.3005
R9577 vss.n2906 vss.n2517 9.3005
R9578 vss.n2910 vss.n2909 9.3005
R9579 vss.n2912 vss.n2911 9.3005
R9580 vss.n2915 vss.n2501 9.3005
R9581 vss.n2919 vss.n2918 9.3005
R9582 vss.n2920 vss.n26 9.3005
R9583 vss.n2922 vss.n2921 9.3005
R9584 vss.n2925 vss.n2485 9.3005
R9585 vss.n2929 vss.n2928 9.3005
R9586 vss.n2931 vss.n2930 9.3005
R9587 vss.n2934 vss.n2470 9.3005
R9588 vss.n2938 vss.n2937 9.3005
R9589 vss.n2940 vss.n2939 9.3005
R9590 vss.n2943 vss.n2458 9.3005
R9591 vss.n2947 vss.n2946 9.3005
R9592 vss.n2949 vss.n2948 9.3005
R9593 vss.n2371 vss.n2362 9.3005
R9594 vss.n2953 vss.n2357 9.3005
R9595 vss.n2956 vss.n2955 9.3005
R9596 vss.n2958 vss.n2957 9.3005
R9597 vss.n2961 vss.n2352 9.3005
R9598 vss.n3003 vss.n2346 9.3005
R9599 vss.n3001 vss.n2964 9.3005
R9600 vss.n2998 vss.n2997 9.3005
R9601 vss.n2996 vss.n2995 9.3005
R9602 vss.n4201 vss.n1328 9.3005
R9603 vss.n4199 vss.n1335 9.3005
R9604 vss.n4196 vss.n4195 9.3005
R9605 vss.n4194 vss.n1338 9.3005
R9606 vss.n4190 vss.n1341 9.3005
R9607 vss.n4187 vss.n4186 9.3005
R9608 vss.n4185 vss.n4184 9.3005
R9609 vss.n4181 vss.n1353 9.3005
R9610 vss.n4178 vss.n4177 9.3005
R9611 vss.n4176 vss.n4175 9.3005
R9612 vss.n4172 vss.n1364 9.3005
R9613 vss.n4169 vss.n4168 9.3005
R9614 vss.n4167 vss.n4166 9.3005
R9615 vss.n4163 vss.n1376 9.3005
R9616 vss.n4160 vss.n4159 9.3005
R9617 vss.n4158 vss.n1386 9.3005
R9618 vss.n4154 vss.n1388 9.3005
R9619 vss.n4151 vss.n4150 9.3005
R9620 vss.n4149 vss.n4148 9.3005
R9621 vss.n4145 vss.n1400 9.3005
R9622 vss.n4142 vss.n4141 9.3005
R9623 vss.n4140 vss.n4139 9.3005
R9624 vss.n4136 vss.n1412 9.3005
R9625 vss.n4133 vss.n4132 9.3005
R9626 vss.n4131 vss.n4130 9.3005
R9627 vss.n4127 vss.n1424 9.3005
R9628 vss.n1445 vss.n1430 9.3005
R9629 vss.n4121 vss.n4120 9.3005
R9630 vss.n4119 vss.n4118 9.3005
R9631 vss.n4115 vss.n1450 9.3005
R9632 vss.n4112 vss.n4111 9.3005
R9633 vss.n4110 vss.n4109 9.3005
R9634 vss.n4106 vss.n1462 9.3005
R9635 vss.n4103 vss.n4102 9.3005
R9636 vss.n4101 vss.n4100 9.3005
R9637 vss.n4097 vss.n1474 9.3005
R9638 vss.n4094 vss.n4093 9.3005
R9639 vss.n4092 vss.n1484 9.3005
R9640 vss.n4088 vss.n1486 9.3005
R9641 vss.n4085 vss.n4084 9.3005
R9642 vss.n4083 vss.n4082 9.3005
R9643 vss.n4079 vss.n1508 9.3005
R9644 vss.n4076 vss.n4075 9.3005
R9645 vss.n4074 vss.n4073 9.3005
R9646 vss.n4070 vss.n1520 9.3005
R9647 vss.n4067 vss.n4066 9.3005
R9648 vss.n4065 vss.n4064 9.3005
R9649 vss.n4061 vss.n1532 9.3005
R9650 vss.n4058 vss.n4057 9.3005
R9651 vss.n4056 vss.n1542 9.3005
R9652 vss.n4052 vss.n1544 9.3005
R9653 vss.n4049 vss.n4048 9.3005
R9654 vss.n4047 vss.n4046 9.3005
R9655 vss.n4043 vss.n1567 9.3005
R9656 vss.n4040 vss.n4039 9.3005
R9657 vss.n4038 vss.n4037 9.3005
R9658 vss.n4034 vss.n1579 9.3005
R9659 vss.n4031 vss.n4030 9.3005
R9660 vss.n4029 vss.n4028 9.3005
R9661 vss.n4025 vss.n1591 9.3005
R9662 vss.n1612 vss.n1597 9.3005
R9663 vss.n4019 vss.n4018 9.3005
R9664 vss.n4017 vss.n4016 9.3005
R9665 vss.n4013 vss.n1617 9.3005
R9666 vss.n4010 vss.n4009 9.3005
R9667 vss.n4008 vss.n4007 9.3005
R9668 vss.n4004 vss.n1629 9.3005
R9669 vss.n4001 vss.n4000 9.3005
R9670 vss.n3999 vss.n3998 9.3005
R9671 vss.n3995 vss.n1641 9.3005
R9672 vss.n3992 vss.n3991 9.3005
R9673 vss.n3990 vss.n1651 9.3005
R9674 vss.n3986 vss.n1653 9.3005
R9675 vss.n3983 vss.n3982 9.3005
R9676 vss.n3981 vss.n3980 9.3005
R9677 vss.n3977 vss.n1675 9.3005
R9678 vss.n3974 vss.n3973 9.3005
R9679 vss.n3972 vss.n3971 9.3005
R9680 vss.n3968 vss.n1687 9.3005
R9681 vss.n3965 vss.n3964 9.3005
R9682 vss.n3963 vss.n3962 9.3005
R9683 vss.n3959 vss.n1699 9.3005
R9684 vss.n3956 vss.n3955 9.3005
R9685 vss.n3954 vss.n1709 9.3005
R9686 vss.n3950 vss.n1711 9.3005
R9687 vss.n3947 vss.n3946 9.3005
R9688 vss.n3945 vss.n3944 9.3005
R9689 vss.n3941 vss.n1734 9.3005
R9690 vss.n3938 vss.n3937 9.3005
R9691 vss.n3936 vss.n3935 9.3005
R9692 vss.n3932 vss.n1746 9.3005
R9693 vss.n3929 vss.n3928 9.3005
R9694 vss.n3927 vss.n3926 9.3005
R9695 vss.n3923 vss.n1758 9.3005
R9696 vss.n1769 vss.n1764 9.3005
R9697 vss.n3917 vss.n3916 9.3005
R9698 vss.n3915 vss.n3914 9.3005
R9699 vss.n3911 vss.n1774 9.3005
R9700 vss.n3908 vss.n3907 9.3005
R9701 vss.n3906 vss.n3905 9.3005
R9702 vss.n3902 vss.n1786 9.3005
R9703 vss.n3899 vss.n3898 9.3005
R9704 vss.n3897 vss.n3896 9.3005
R9705 vss.n3893 vss.n1798 9.3005
R9706 vss.n3890 vss.n3889 9.3005
R9707 vss.n3888 vss.n3887 9.3005
R9708 vss.n1812 vss.n1810 9.3005
R9709 vss.n3881 vss.n3880 9.3005
R9710 vss.n3879 vss.n3878 9.3005
R9711 vss.n3875 vss.n1833 9.3005
R9712 vss.n3872 vss.n3871 9.3005
R9713 vss.n3870 vss.n3869 9.3005
R9714 vss.n3866 vss.n1845 9.3005
R9715 vss.n3863 vss.n3862 9.3005
R9716 vss.n3861 vss.n3860 9.3005
R9717 vss.n3857 vss.n1857 9.3005
R9718 vss.n3854 vss.n3853 9.3005
R9719 vss.n3852 vss.n1867 9.3005
R9720 vss.n3848 vss.n1869 9.3005
R9721 vss.n3845 vss.n3844 9.3005
R9722 vss.n3843 vss.n3842 9.3005
R9723 vss.n3839 vss.n1891 9.3005
R9724 vss.n3836 vss.n3835 9.3005
R9725 vss.n3834 vss.n3833 9.3005
R9726 vss.n3830 vss.n1903 9.3005
R9727 vss.n3827 vss.n3826 9.3005
R9728 vss.n3825 vss.n3824 9.3005
R9729 vss.n3821 vss.n1915 9.3005
R9730 vss.n1936 vss.n1921 9.3005
R9731 vss.n3815 vss.n3814 9.3005
R9732 vss.n3813 vss.n3812 9.3005
R9733 vss.n3809 vss.n1941 9.3005
R9734 vss.n3806 vss.n3805 9.3005
R9735 vss.n3804 vss.n3803 9.3005
R9736 vss.n3800 vss.n1953 9.3005
R9737 vss.n3797 vss.n3796 9.3005
R9738 vss.n3795 vss.n3794 9.3005
R9739 vss.n3791 vss.n1965 9.3005
R9740 vss.n3788 vss.n3787 9.3005
R9741 vss.n3786 vss.n3785 9.3005
R9742 vss.n1979 vss.n1977 9.3005
R9743 vss.n3779 vss.n3778 9.3005
R9744 vss.n3777 vss.n3776 9.3005
R9745 vss.n3773 vss.n2000 9.3005
R9746 vss.n3770 vss.n3769 9.3005
R9747 vss.n3768 vss.n3767 9.3005
R9748 vss.n3764 vss.n2012 9.3005
R9749 vss.n3761 vss.n3760 9.3005
R9750 vss.n3759 vss.n3758 9.3005
R9751 vss.n3755 vss.n2024 9.3005
R9752 vss.n3752 vss.n3751 9.3005
R9753 vss.n3750 vss.n2034 9.3005
R9754 vss.n3746 vss.n2036 9.3005
R9755 vss.n3743 vss.n3742 9.3005
R9756 vss.n3741 vss.n3740 9.3005
R9757 vss.n3737 vss.n2058 9.3005
R9758 vss.n3734 vss.n3733 9.3005
R9759 vss.n3732 vss.n3731 9.3005
R9760 vss.n3728 vss.n2070 9.3005
R9761 vss.n3725 vss.n3724 9.3005
R9762 vss.n3723 vss.n3722 9.3005
R9763 vss.n3719 vss.n2082 9.3005
R9764 vss.n2103 vss.n2088 9.3005
R9765 vss.n3713 vss.n3712 9.3005
R9766 vss.n3711 vss.n3710 9.3005
R9767 vss.n3707 vss.n2108 9.3005
R9768 vss.n3704 vss.n3703 9.3005
R9769 vss.n3702 vss.n3701 9.3005
R9770 vss.n3698 vss.n2120 9.3005
R9771 vss.n3695 vss.n3694 9.3005
R9772 vss.n3693 vss.n3692 9.3005
R9773 vss.n3689 vss.n2132 9.3005
R9774 vss.n3686 vss.n3685 9.3005
R9775 vss.n3684 vss.n3683 9.3005
R9776 vss.n2146 vss.n2144 9.3005
R9777 vss.n3677 vss.n3676 9.3005
R9778 vss.n3675 vss.n3674 9.3005
R9779 vss.n3671 vss.n2156 9.3005
R9780 vss.n3668 vss.n3667 9.3005
R9781 vss.n3666 vss.n3665 9.3005
R9782 vss.n3662 vss.n2168 9.3005
R9783 vss.n3659 vss.n3658 9.3005
R9784 vss.n3657 vss.n3656 9.3005
R9785 vss.n3653 vss.n2180 9.3005
R9786 vss.n3650 vss.n3649 9.3005
R9787 vss.n3648 vss.n2190 9.3005
R9788 vss.n3606 vss.n3078 9.3005
R9789 vss.n3610 vss.n3609 9.3005
R9790 vss.n3613 vss.n3612 9.3005
R9791 vss.n3611 vss.n3071 9.3005
R9792 vss.n3617 vss.n3067 9.3005
R9793 vss.n3621 vss.n3620 9.3005
R9794 vss.n3623 vss.n3622 9.3005
R9795 vss.n3626 vss.n3058 9.3005
R9796 vss.n3630 vss.n3629 9.3005
R9797 vss.n3632 vss.n3631 9.3005
R9798 vss.n3635 vss.n3049 9.3005
R9799 vss.n3639 vss.n3638 9.3005
R9800 vss.n3641 vss.n3640 9.3005
R9801 vss.n3644 vss.n2192 9.3005
R9802 vss.n6011 vss.n131 9.3005
R9803 vss.n5981 vss.n130 9.3005
R9804 vss.n5987 vss.n5982 9.3005
R9805 vss.n5990 vss.n5978 9.3005
R9806 vss.n5992 vss.n5976 9.3005
R9807 vss.n5995 vss.n5972 9.3005
R9808 vss.n5998 vss.n5968 9.3005
R9809 vss.n6000 vss.n147 9.3005
R9810 vss.n5966 vss.n155 9.3005
R9811 vss.n5963 vss.n160 9.3005
R9812 vss.n5960 vss.n165 9.3005
R9813 vss.n5956 vss.n164 9.3005
R9814 vss.n5955 vss.n5954 9.3005
R9815 vss.n5951 vss.n170 9.3005
R9816 vss.n5948 vss.n181 9.3005
R9817 vss.n5945 vss.n185 9.3005
R9818 vss.n5942 vss.n188 9.3005
R9819 vss.n5939 vss.n192 9.3005
R9820 vss.n5936 vss.n195 9.3005
R9821 vss.n5933 vss.n198 9.3005
R9822 vss.n5930 vss.n202 9.3005
R9823 vss.n5927 vss.n205 9.3005
R9824 vss.n5924 vss.n209 9.3005
R9825 vss.n212 vss.n208 9.3005
R9826 vss.n2768 vss.n2767 9.3005
R9827 vss.n2771 vss.n2766 9.3005
R9828 vss.n2774 vss.n2759 9.3005
R9829 vss.n2777 vss.n2753 9.3005
R9830 vss.n2780 vss.n2750 9.3005
R9831 vss.n2783 vss.n2744 9.3005
R9832 vss.n2786 vss.n2740 9.3005
R9833 vss.n2789 vss.n2734 9.3005
R9834 vss.n2792 vss.n2730 9.3005
R9835 vss.n2795 vss.n2722 9.3005
R9836 vss.n2796 vss.n2720 9.3005
R9837 vss.n2799 vss.n2713 9.3005
R9838 vss.n2802 vss.n2710 9.3005
R9839 vss.n2805 vss.n2704 9.3005
R9840 vss.n2808 vss.n2701 9.3005
R9841 vss.n2811 vss.n2694 9.3005
R9842 vss.n2814 vss.n2691 9.3005
R9843 vss.n2817 vss.n2684 9.3005
R9844 vss.n2820 vss.n2676 9.3005
R9845 vss.n2822 vss.n2674 9.3005
R9846 vss.n2825 vss.n2669 9.3005
R9847 vss.n2668 vss.n65 9.3005
R9848 vss.n2829 vss.n2659 9.3005
R9849 vss.n2832 vss.n2651 9.3005
R9850 vss.n2834 vss.n2649 9.3005
R9851 vss.n2837 vss.n2646 9.3005
R9852 vss.n2840 vss.n2639 9.3005
R9853 vss.n2843 vss.n2636 9.3005
R9854 vss.n2846 vss.n2629 9.3005
R9855 vss.n2849 vss.n2626 9.3005
R9856 vss.n2852 vss.n2620 9.3005
R9857 vss.n2855 vss.n2615 9.3005
R9858 vss.n2614 vss.n2606 9.3005
R9859 vss.n2859 vss.n2605 9.3005
R9860 vss.n2862 vss.n2599 9.3005
R9861 vss.n2865 vss.n2596 9.3005
R9862 vss.n2868 vss.n2590 9.3005
R9863 vss.n2871 vss.n2586 9.3005
R9864 vss.n2874 vss.n2580 9.3005
R9865 vss.n2877 vss.n2576 9.3005
R9866 vss.n2880 vss.n2570 9.3005
R9867 vss.n2882 vss.n2568 9.3005
R9868 vss.n2885 vss.n2561 9.3005
R9869 vss.n2888 vss.n2553 9.3005
R9870 vss.n2889 vss.n2551 9.3005
R9871 vss.n2892 vss.n2548 9.3005
R9872 vss.n2895 vss.n2540 9.3005
R9873 vss.n2898 vss.n2537 9.3005
R9874 vss.n2901 vss.n2533 9.3005
R9875 vss.n2904 vss.n2526 9.3005
R9876 vss.n2906 vss.n2524 9.3005
R9877 vss.n2909 vss.n2518 9.3005
R9878 vss.n2912 vss.n2515 9.3005
R9879 vss.n2915 vss.n2509 9.3005
R9880 vss.n2918 vss.n2503 9.3005
R9881 vss.n2502 vss.n26 9.3005
R9882 vss.n2922 vss.n2495 9.3005
R9883 vss.n2925 vss.n2489 9.3005
R9884 vss.n2928 vss.n2486 9.3005
R9885 vss.n2931 vss.n2479 9.3005
R9886 vss.n2934 vss.n2476 9.3005
R9887 vss.n2937 vss.n2471 9.3005
R9888 vss.n2940 vss.n2468 9.3005
R9889 vss.n2943 vss.n2464 9.3005
R9890 vss.n2946 vss.n2459 9.3005
R9891 vss.n2949 vss.n2368 9.3005
R9892 vss.n2367 vss.n2362 9.3005
R9893 vss.n2953 vss.n2360 9.3005
R9894 vss.n2955 vss.n2358 9.3005
R9895 vss.n2958 vss.n2355 9.3005
R9896 vss.n2961 vss.n2351 9.3005
R9897 vss.n3003 vss.n2348 9.3005
R9898 vss.n3001 vss.n2963 9.3005
R9899 vss.n2998 vss.n2992 9.3005
R9900 vss.n2995 vss.n2994 9.3005
R9901 vss.n4201 vss.n1330 9.3005
R9902 vss.n4199 vss.n1334 9.3005
R9903 vss.n4196 vss.n1339 9.3005
R9904 vss.n1344 vss.n1338 9.3005
R9905 vss.n4190 vss.n1347 9.3005
R9906 vss.n4187 vss.n1352 9.3005
R9907 vss.n4184 vss.n1356 9.3005
R9908 vss.n4181 vss.n1359 9.3005
R9909 vss.n4178 vss.n1363 9.3005
R9910 vss.n4175 vss.n1367 9.3005
R9911 vss.n4172 vss.n1371 9.3005
R9912 vss.n4169 vss.n1375 9.3005
R9913 vss.n4166 vss.n1379 9.3005
R9914 vss.n4163 vss.n1383 9.3005
R9915 vss.n4160 vss.n1387 9.3005
R9916 vss.n1391 vss.n1386 9.3005
R9917 vss.n4154 vss.n1394 9.3005
R9918 vss.n4151 vss.n1399 9.3005
R9919 vss.n4148 vss.n1403 9.3005
R9920 vss.n4145 vss.n1407 9.3005
R9921 vss.n4142 vss.n1411 9.3005
R9922 vss.n4139 vss.n1415 9.3005
R9923 vss.n4136 vss.n1419 9.3005
R9924 vss.n4133 vss.n1423 9.3005
R9925 vss.n4130 vss.n1427 9.3005
R9926 vss.n4127 vss.n1431 9.3005
R9927 vss.n4123 vss.n1430 9.3005
R9928 vss.n4122 vss.n4121 9.3005
R9929 vss.n4118 vss.n1446 9.3005
R9930 vss.n4115 vss.n1457 9.3005
R9931 vss.n4112 vss.n1461 9.3005
R9932 vss.n4109 vss.n1465 9.3005
R9933 vss.n4106 vss.n1469 9.3005
R9934 vss.n4103 vss.n1473 9.3005
R9935 vss.n4100 vss.n1477 9.3005
R9936 vss.n4097 vss.n1481 9.3005
R9937 vss.n4094 vss.n1485 9.3005
R9938 vss.n4090 vss.n1484 9.3005
R9939 vss.n4089 vss.n4088 9.3005
R9940 vss.n4085 vss.n1500 9.3005
R9941 vss.n4082 vss.n1511 9.3005
R9942 vss.n4079 vss.n1515 9.3005
R9943 vss.n4076 vss.n1519 9.3005
R9944 vss.n4073 vss.n1523 9.3005
R9945 vss.n4070 vss.n1527 9.3005
R9946 vss.n4067 vss.n1531 9.3005
R9947 vss.n4064 vss.n1535 9.3005
R9948 vss.n4061 vss.n1539 9.3005
R9949 vss.n4058 vss.n1543 9.3005
R9950 vss.n1558 vss.n1542 9.3005
R9951 vss.n4052 vss.n1561 9.3005
R9952 vss.n4049 vss.n1566 9.3005
R9953 vss.n4046 vss.n1570 9.3005
R9954 vss.n4043 vss.n1574 9.3005
R9955 vss.n4040 vss.n1578 9.3005
R9956 vss.n4037 vss.n1582 9.3005
R9957 vss.n4034 vss.n1586 9.3005
R9958 vss.n4031 vss.n1590 9.3005
R9959 vss.n4028 vss.n1594 9.3005
R9960 vss.n4025 vss.n1598 9.3005
R9961 vss.n4021 vss.n1597 9.3005
R9962 vss.n4020 vss.n4019 9.3005
R9963 vss.n4016 vss.n1613 9.3005
R9964 vss.n4013 vss.n1624 9.3005
R9965 vss.n4010 vss.n1628 9.3005
R9966 vss.n4007 vss.n1632 9.3005
R9967 vss.n4004 vss.n1636 9.3005
R9968 vss.n4001 vss.n1640 9.3005
R9969 vss.n3998 vss.n1644 9.3005
R9970 vss.n3995 vss.n1648 9.3005
R9971 vss.n3992 vss.n1652 9.3005
R9972 vss.n3988 vss.n1651 9.3005
R9973 vss.n3987 vss.n3986 9.3005
R9974 vss.n3983 vss.n1667 9.3005
R9975 vss.n3980 vss.n1678 9.3005
R9976 vss.n3977 vss.n1682 9.3005
R9977 vss.n3974 vss.n1686 9.3005
R9978 vss.n3971 vss.n1690 9.3005
R9979 vss.n3968 vss.n1694 9.3005
R9980 vss.n3965 vss.n1698 9.3005
R9981 vss.n3962 vss.n1702 9.3005
R9982 vss.n3959 vss.n1706 9.3005
R9983 vss.n3956 vss.n1710 9.3005
R9984 vss.n1725 vss.n1709 9.3005
R9985 vss.n3950 vss.n1728 9.3005
R9986 vss.n3947 vss.n1733 9.3005
R9987 vss.n3944 vss.n1737 9.3005
R9988 vss.n3941 vss.n1741 9.3005
R9989 vss.n3938 vss.n1745 9.3005
R9990 vss.n3935 vss.n1749 9.3005
R9991 vss.n3932 vss.n1753 9.3005
R9992 vss.n3929 vss.n1757 9.3005
R9993 vss.n3926 vss.n1761 9.3005
R9994 vss.n3923 vss.n1765 9.3005
R9995 vss.n3919 vss.n1764 9.3005
R9996 vss.n3918 vss.n3917 9.3005
R9997 vss.n3914 vss.n1770 9.3005
R9998 vss.n3911 vss.n1781 9.3005
R9999 vss.n3908 vss.n1785 9.3005
R10000 vss.n3905 vss.n1789 9.3005
R10001 vss.n3902 vss.n1793 9.3005
R10002 vss.n3899 vss.n1797 9.3005
R10003 vss.n3896 vss.n1801 9.3005
R10004 vss.n3893 vss.n1805 9.3005
R10005 vss.n3890 vss.n1809 9.3005
R10006 vss.n3887 vss.n1813 9.3005
R10007 vss.n1828 vss.n1812 9.3005
R10008 vss.n3881 vss.n1831 9.3005
R10009 vss.n3878 vss.n1836 9.3005
R10010 vss.n3875 vss.n1840 9.3005
R10011 vss.n3872 vss.n1844 9.3005
R10012 vss.n3869 vss.n1848 9.3005
R10013 vss.n3866 vss.n1852 9.3005
R10014 vss.n3863 vss.n1856 9.3005
R10015 vss.n3860 vss.n1860 9.3005
R10016 vss.n3857 vss.n1864 9.3005
R10017 vss.n3854 vss.n1868 9.3005
R10018 vss.n3850 vss.n1867 9.3005
R10019 vss.n3849 vss.n3848 9.3005
R10020 vss.n3845 vss.n1883 9.3005
R10021 vss.n3842 vss.n1894 9.3005
R10022 vss.n3839 vss.n1898 9.3005
R10023 vss.n3836 vss.n1902 9.3005
R10024 vss.n3833 vss.n1906 9.3005
R10025 vss.n3830 vss.n1910 9.3005
R10026 vss.n3827 vss.n1914 9.3005
R10027 vss.n3824 vss.n1918 9.3005
R10028 vss.n3821 vss.n1922 9.3005
R10029 vss.n3817 vss.n1921 9.3005
R10030 vss.n3816 vss.n3815 9.3005
R10031 vss.n3812 vss.n1937 9.3005
R10032 vss.n3809 vss.n1948 9.3005
R10033 vss.n3806 vss.n1952 9.3005
R10034 vss.n3803 vss.n1956 9.3005
R10035 vss.n3800 vss.n1960 9.3005
R10036 vss.n3797 vss.n1964 9.3005
R10037 vss.n3794 vss.n1968 9.3005
R10038 vss.n3791 vss.n1972 9.3005
R10039 vss.n3788 vss.n1976 9.3005
R10040 vss.n3785 vss.n1980 9.3005
R10041 vss.n1995 vss.n1979 9.3005
R10042 vss.n3779 vss.n1998 9.3005
R10043 vss.n3776 vss.n2003 9.3005
R10044 vss.n3773 vss.n2007 9.3005
R10045 vss.n3770 vss.n2011 9.3005
R10046 vss.n3767 vss.n2015 9.3005
R10047 vss.n3764 vss.n2019 9.3005
R10048 vss.n3761 vss.n2023 9.3005
R10049 vss.n3758 vss.n2027 9.3005
R10050 vss.n3755 vss.n2031 9.3005
R10051 vss.n3752 vss.n2035 9.3005
R10052 vss.n3748 vss.n2034 9.3005
R10053 vss.n3747 vss.n3746 9.3005
R10054 vss.n3743 vss.n2050 9.3005
R10055 vss.n3740 vss.n2061 9.3005
R10056 vss.n3737 vss.n2065 9.3005
R10057 vss.n3734 vss.n2069 9.3005
R10058 vss.n3731 vss.n2073 9.3005
R10059 vss.n3728 vss.n2077 9.3005
R10060 vss.n3725 vss.n2081 9.3005
R10061 vss.n3722 vss.n2085 9.3005
R10062 vss.n3719 vss.n2089 9.3005
R10063 vss.n3715 vss.n2088 9.3005
R10064 vss.n3714 vss.n3713 9.3005
R10065 vss.n3710 vss.n2104 9.3005
R10066 vss.n3707 vss.n2115 9.3005
R10067 vss.n3704 vss.n2119 9.3005
R10068 vss.n3701 vss.n2123 9.3005
R10069 vss.n3698 vss.n2127 9.3005
R10070 vss.n3695 vss.n2131 9.3005
R10071 vss.n3692 vss.n2135 9.3005
R10072 vss.n3689 vss.n2139 9.3005
R10073 vss.n3686 vss.n2143 9.3005
R10074 vss.n3683 vss.n2147 9.3005
R10075 vss.n2151 vss.n2146 9.3005
R10076 vss.n3677 vss.n2154 9.3005
R10077 vss.n3674 vss.n2159 9.3005
R10078 vss.n3671 vss.n2163 9.3005
R10079 vss.n3668 vss.n2167 9.3005
R10080 vss.n3665 vss.n2171 9.3005
R10081 vss.n3662 vss.n2175 9.3005
R10082 vss.n3659 vss.n2179 9.3005
R10083 vss.n3656 vss.n2183 9.3005
R10084 vss.n3653 vss.n2187 9.3005
R10085 vss.n3650 vss.n2191 9.3005
R10086 vss.n3646 vss.n2190 9.3005
R10087 vss.n3606 vss.n3604 9.3005
R10088 vss.n3609 vss.n3080 9.3005
R10089 vss.n3613 vss.n3076 9.3005
R10090 vss.n3075 vss.n3071 9.3005
R10091 vss.n3617 vss.n3072 9.3005
R10092 vss.n3620 vss.n3069 9.3005
R10093 vss.n3623 vss.n3066 9.3005
R10094 vss.n3626 vss.n3063 9.3005
R10095 vss.n3629 vss.n3060 9.3005
R10096 vss.n3632 vss.n3057 9.3005
R10097 vss.n3635 vss.n3054 9.3005
R10098 vss.n3638 vss.n3051 9.3005
R10099 vss.n3641 vss.n3042 9.3005
R10100 vss.n3645 vss.n3644 9.3005
R10101 vss.n3606 vss.n3605 9.3005
R10102 vss.n3609 vss.n3073 9.3005
R10103 vss.n3614 vss.n3613 9.3005
R10104 vss.n3615 vss.n3071 9.3005
R10105 vss.n3617 vss.n3616 9.3005
R10106 vss.n3620 vss.n3064 9.3005
R10107 vss.n3624 vss.n3623 9.3005
R10108 vss.n3626 vss.n3625 9.3005
R10109 vss.n3629 vss.n3055 9.3005
R10110 vss.n3633 vss.n3632 9.3005
R10111 vss.n3635 vss.n3634 9.3005
R10112 vss.n3638 vss.n3046 9.3005
R10113 vss.n3642 vss.n3641 9.3005
R10114 vss.n3644 vss.n3643 9.3005
R10115 vss.n3041 vss.n2190 9.3005
R10116 vss.n3650 vss.n2184 9.3005
R10117 vss.n3654 vss.n3653 9.3005
R10118 vss.n3656 vss.n3655 9.3005
R10119 vss.n3659 vss.n2172 9.3005
R10120 vss.n3663 vss.n3662 9.3005
R10121 vss.n3665 vss.n3664 9.3005
R10122 vss.n3668 vss.n2160 9.3005
R10123 vss.n3672 vss.n3671 9.3005
R10124 vss.n3674 vss.n3673 9.3005
R10125 vss.n3677 vss.n2148 9.3005
R10126 vss.n3681 vss.n2146 9.3005
R10127 vss.n3683 vss.n3682 9.3005
R10128 vss.n3686 vss.n2136 9.3005
R10129 vss.n3690 vss.n3689 9.3005
R10130 vss.n3692 vss.n3691 9.3005
R10131 vss.n3695 vss.n2124 9.3005
R10132 vss.n3699 vss.n3698 9.3005
R10133 vss.n3701 vss.n3700 9.3005
R10134 vss.n3704 vss.n2112 9.3005
R10135 vss.n3708 vss.n3707 9.3005
R10136 vss.n3710 vss.n3709 9.3005
R10137 vss.n3713 vss.n2090 9.3005
R10138 vss.n3717 vss.n2088 9.3005
R10139 vss.n3719 vss.n3718 9.3005
R10140 vss.n3722 vss.n2078 9.3005
R10141 vss.n3726 vss.n3725 9.3005
R10142 vss.n3728 vss.n3727 9.3005
R10143 vss.n3731 vss.n2066 9.3005
R10144 vss.n3735 vss.n3734 9.3005
R10145 vss.n3737 vss.n3736 9.3005
R10146 vss.n3740 vss.n2054 9.3005
R10147 vss.n3744 vss.n3743 9.3005
R10148 vss.n3746 vss.n3745 9.3005
R10149 vss.n2049 vss.n2034 9.3005
R10150 vss.n3752 vss.n2028 9.3005
R10151 vss.n3756 vss.n3755 9.3005
R10152 vss.n3758 vss.n3757 9.3005
R10153 vss.n3761 vss.n2016 9.3005
R10154 vss.n3765 vss.n3764 9.3005
R10155 vss.n3767 vss.n3766 9.3005
R10156 vss.n3770 vss.n2004 9.3005
R10157 vss.n3774 vss.n3773 9.3005
R10158 vss.n3776 vss.n3775 9.3005
R10159 vss.n3779 vss.n1981 9.3005
R10160 vss.n3783 vss.n1979 9.3005
R10161 vss.n3785 vss.n3784 9.3005
R10162 vss.n3788 vss.n1969 9.3005
R10163 vss.n3792 vss.n3791 9.3005
R10164 vss.n3794 vss.n3793 9.3005
R10165 vss.n3797 vss.n1957 9.3005
R10166 vss.n3801 vss.n3800 9.3005
R10167 vss.n3803 vss.n3802 9.3005
R10168 vss.n3806 vss.n1945 9.3005
R10169 vss.n3810 vss.n3809 9.3005
R10170 vss.n3812 vss.n3811 9.3005
R10171 vss.n3815 vss.n1923 9.3005
R10172 vss.n3819 vss.n1921 9.3005
R10173 vss.n3821 vss.n3820 9.3005
R10174 vss.n3824 vss.n1911 9.3005
R10175 vss.n3828 vss.n3827 9.3005
R10176 vss.n3830 vss.n3829 9.3005
R10177 vss.n3833 vss.n1899 9.3005
R10178 vss.n3837 vss.n3836 9.3005
R10179 vss.n3839 vss.n3838 9.3005
R10180 vss.n3842 vss.n1887 9.3005
R10181 vss.n3846 vss.n3845 9.3005
R10182 vss.n3848 vss.n3847 9.3005
R10183 vss.n1882 vss.n1867 9.3005
R10184 vss.n3854 vss.n1861 9.3005
R10185 vss.n3858 vss.n3857 9.3005
R10186 vss.n3860 vss.n3859 9.3005
R10187 vss.n3863 vss.n1849 9.3005
R10188 vss.n3867 vss.n3866 9.3005
R10189 vss.n3869 vss.n3868 9.3005
R10190 vss.n3872 vss.n1837 9.3005
R10191 vss.n3876 vss.n3875 9.3005
R10192 vss.n3878 vss.n3877 9.3005
R10193 vss.n3881 vss.n1814 9.3005
R10194 vss.n3885 vss.n1812 9.3005
R10195 vss.n3887 vss.n3886 9.3005
R10196 vss.n3890 vss.n1802 9.3005
R10197 vss.n3894 vss.n3893 9.3005
R10198 vss.n3896 vss.n3895 9.3005
R10199 vss.n3899 vss.n1790 9.3005
R10200 vss.n3903 vss.n3902 9.3005
R10201 vss.n3905 vss.n3904 9.3005
R10202 vss.n3908 vss.n1778 9.3005
R10203 vss.n3912 vss.n3911 9.3005
R10204 vss.n3914 vss.n3913 9.3005
R10205 vss.n3917 vss.n1766 9.3005
R10206 vss.n3921 vss.n1764 9.3005
R10207 vss.n3923 vss.n3922 9.3005
R10208 vss.n3926 vss.n1754 9.3005
R10209 vss.n3930 vss.n3929 9.3005
R10210 vss.n3932 vss.n3931 9.3005
R10211 vss.n3935 vss.n1742 9.3005
R10212 vss.n3939 vss.n3938 9.3005
R10213 vss.n3941 vss.n3940 9.3005
R10214 vss.n3944 vss.n1730 9.3005
R10215 vss.n3948 vss.n3947 9.3005
R10216 vss.n3950 vss.n3949 9.3005
R10217 vss.n1709 vss.n1707 9.3005
R10218 vss.n3957 vss.n3956 9.3005
R10219 vss.n3959 vss.n3958 9.3005
R10220 vss.n3962 vss.n1695 9.3005
R10221 vss.n3966 vss.n3965 9.3005
R10222 vss.n3968 vss.n3967 9.3005
R10223 vss.n3971 vss.n1683 9.3005
R10224 vss.n3975 vss.n3974 9.3005
R10225 vss.n3977 vss.n3976 9.3005
R10226 vss.n3980 vss.n1671 9.3005
R10227 vss.n3984 vss.n3983 9.3005
R10228 vss.n3986 vss.n3985 9.3005
R10229 vss.n1666 vss.n1651 9.3005
R10230 vss.n3992 vss.n1645 9.3005
R10231 vss.n3996 vss.n3995 9.3005
R10232 vss.n3998 vss.n3997 9.3005
R10233 vss.n4001 vss.n1633 9.3005
R10234 vss.n4005 vss.n4004 9.3005
R10235 vss.n4007 vss.n4006 9.3005
R10236 vss.n4010 vss.n1621 9.3005
R10237 vss.n4014 vss.n4013 9.3005
R10238 vss.n4016 vss.n4015 9.3005
R10239 vss.n4019 vss.n1599 9.3005
R10240 vss.n4023 vss.n1597 9.3005
R10241 vss.n4025 vss.n4024 9.3005
R10242 vss.n4028 vss.n1587 9.3005
R10243 vss.n4032 vss.n4031 9.3005
R10244 vss.n4034 vss.n4033 9.3005
R10245 vss.n4037 vss.n1575 9.3005
R10246 vss.n4041 vss.n4040 9.3005
R10247 vss.n4043 vss.n4042 9.3005
R10248 vss.n4046 vss.n1563 9.3005
R10249 vss.n4050 vss.n4049 9.3005
R10250 vss.n4052 vss.n4051 9.3005
R10251 vss.n1542 vss.n1540 9.3005
R10252 vss.n4059 vss.n4058 9.3005
R10253 vss.n4061 vss.n4060 9.3005
R10254 vss.n4064 vss.n1528 9.3005
R10255 vss.n4068 vss.n4067 9.3005
R10256 vss.n4070 vss.n4069 9.3005
R10257 vss.n4073 vss.n1516 9.3005
R10258 vss.n4077 vss.n4076 9.3005
R10259 vss.n4079 vss.n4078 9.3005
R10260 vss.n4082 vss.n1504 9.3005
R10261 vss.n4086 vss.n4085 9.3005
R10262 vss.n4088 vss.n4087 9.3005
R10263 vss.n1499 vss.n1484 9.3005
R10264 vss.n4094 vss.n1478 9.3005
R10265 vss.n4098 vss.n4097 9.3005
R10266 vss.n4100 vss.n4099 9.3005
R10267 vss.n4103 vss.n1466 9.3005
R10268 vss.n4107 vss.n4106 9.3005
R10269 vss.n4109 vss.n4108 9.3005
R10270 vss.n4112 vss.n1454 9.3005
R10271 vss.n4116 vss.n4115 9.3005
R10272 vss.n4118 vss.n4117 9.3005
R10273 vss.n4121 vss.n1432 9.3005
R10274 vss.n4125 vss.n1430 9.3005
R10275 vss.n4127 vss.n4126 9.3005
R10276 vss.n4130 vss.n1420 9.3005
R10277 vss.n4134 vss.n4133 9.3005
R10278 vss.n4136 vss.n4135 9.3005
R10279 vss.n4139 vss.n1408 9.3005
R10280 vss.n4143 vss.n4142 9.3005
R10281 vss.n4145 vss.n4144 9.3005
R10282 vss.n4148 vss.n1396 9.3005
R10283 vss.n4152 vss.n4151 9.3005
R10284 vss.n4154 vss.n4153 9.3005
R10285 vss.n1386 vss.n1384 9.3005
R10286 vss.n4161 vss.n4160 9.3005
R10287 vss.n4163 vss.n4162 9.3005
R10288 vss.n4166 vss.n1372 9.3005
R10289 vss.n4170 vss.n4169 9.3005
R10290 vss.n4172 vss.n4171 9.3005
R10291 vss.n4175 vss.n1360 9.3005
R10292 vss.n4179 vss.n4178 9.3005
R10293 vss.n4181 vss.n4180 9.3005
R10294 vss.n4184 vss.n1349 9.3005
R10295 vss.n4188 vss.n4187 9.3005
R10296 vss.n4190 vss.n4189 9.3005
R10297 vss.n1338 vss.n1336 9.3005
R10298 vss.n4197 vss.n4196 9.3005
R10299 vss.n4199 vss.n4198 9.3005
R10300 vss.n4201 vss.n1327 9.3005
R10301 vss.n2995 vss.n2965 9.3005
R10302 vss.n2999 vss.n2998 9.3005
R10303 vss.n3001 vss.n3000 9.3005
R10304 vss.n3003 vss.n2345 9.3005
R10305 vss.n2961 vss.n2960 9.3005
R10306 vss.n2959 vss.n2958 9.3005
R10307 vss.n2955 vss.n2354 9.3005
R10308 vss.n2953 vss.n2952 9.3005
R10309 vss.n2951 vss.n2362 9.3005
R10310 vss.n2950 vss.n2949 9.3005
R10311 vss.n2946 vss.n2366 9.3005
R10312 vss.n2943 vss.n2942 9.3005
R10313 vss.n2941 vss.n2940 9.3005
R10314 vss.n2937 vss.n2467 9.3005
R10315 vss.n2934 vss.n2933 9.3005
R10316 vss.n2932 vss.n2931 9.3005
R10317 vss.n2928 vss.n2478 9.3005
R10318 vss.n2925 vss.n2924 9.3005
R10319 vss.n2923 vss.n2922 9.3005
R10320 vss.n2494 vss.n26 9.3005
R10321 vss.n2918 vss.n2917 9.3005
R10322 vss.n2916 vss.n2915 9.3005
R10323 vss.n2912 vss.n2508 9.3005
R10324 vss.n2909 vss.n2908 9.3005
R10325 vss.n2907 vss.n2906 9.3005
R10326 vss.n2904 vss.n2523 9.3005
R10327 vss.n2901 vss.n2900 9.3005
R10328 vss.n2899 vss.n2898 9.3005
R10329 vss.n2895 vss.n2536 9.3005
R10330 vss.n2892 vss.n2891 9.3005
R10331 vss.n2890 vss.n2889 9.3005
R10332 vss.n2888 vss.n2550 9.3005
R10333 vss.n2885 vss.n2884 9.3005
R10334 vss.n2883 vss.n2882 9.3005
R10335 vss.n2880 vss.n2567 9.3005
R10336 vss.n2877 vss.n2876 9.3005
R10337 vss.n2875 vss.n2874 9.3005
R10338 vss.n2871 vss.n2579 9.3005
R10339 vss.n2868 vss.n2867 9.3005
R10340 vss.n2866 vss.n2865 9.3005
R10341 vss.n2862 vss.n2595 9.3005
R10342 vss.n2859 vss.n2858 9.3005
R10343 vss.n2857 vss.n2606 9.3005
R10344 vss.n2856 vss.n2855 9.3005
R10345 vss.n2852 vss.n2612 9.3005
R10346 vss.n2849 vss.n2848 9.3005
R10347 vss.n2847 vss.n2846 9.3005
R10348 vss.n2843 vss.n2628 9.3005
R10349 vss.n2840 vss.n2839 9.3005
R10350 vss.n2838 vss.n2837 9.3005
R10351 vss.n2834 vss.n2645 9.3005
R10352 vss.n2832 vss.n2831 9.3005
R10353 vss.n2830 vss.n2829 9.3005
R10354 vss.n2658 vss.n65 9.3005
R10355 vss.n2825 vss.n2824 9.3005
R10356 vss.n2823 vss.n2822 9.3005
R10357 vss.n2820 vss.n2673 9.3005
R10358 vss.n2817 vss.n2816 9.3005
R10359 vss.n2815 vss.n2814 9.3005
R10360 vss.n2811 vss.n2690 9.3005
R10361 vss.n2808 vss.n2807 9.3005
R10362 vss.n2806 vss.n2805 9.3005
R10363 vss.n2802 vss.n2703 9.3005
R10364 vss.n2799 vss.n2798 9.3005
R10365 vss.n2797 vss.n2796 9.3005
R10366 vss.n2795 vss.n2719 9.3005
R10367 vss.n2792 vss.n2791 9.3005
R10368 vss.n2790 vss.n2789 9.3005
R10369 vss.n2786 vss.n2733 9.3005
R10370 vss.n2783 vss.n2782 9.3005
R10371 vss.n2781 vss.n2780 9.3005
R10372 vss.n2777 vss.n2749 9.3005
R10373 vss.n2774 vss.n2773 9.3005
R10374 vss.n2772 vss.n2771 9.3005
R10375 vss.n2768 vss.n2765 9.3005
R10376 vss.n208 vss.n206 9.3005
R10377 vss.n5925 vss.n5924 9.3005
R10378 vss.n5927 vss.n5926 9.3005
R10379 vss.n5930 vss.n196 9.3005
R10380 vss.n5934 vss.n5933 9.3005
R10381 vss.n5936 vss.n5935 9.3005
R10382 vss.n5939 vss.n186 9.3005
R10383 vss.n5943 vss.n5942 9.3005
R10384 vss.n5945 vss.n5944 9.3005
R10385 vss.n5948 vss.n174 9.3005
R10386 vss.n5952 vss.n5951 9.3005
R10387 vss.n5954 vss.n5953 9.3005
R10388 vss.n169 vss.n164 9.3005
R10389 vss.n5960 vss.n157 9.3005
R10390 vss.n5964 vss.n5963 9.3005
R10391 vss.n5966 vss.n5965 9.3005
R10392 vss.n6000 vss.n145 9.3005
R10393 vss.n5998 vss.n5997 9.3005
R10394 vss.n5996 vss.n5995 9.3005
R10395 vss.n5992 vss.n5971 9.3005
R10396 vss.n5990 vss.n5989 9.3005
R10397 vss.n5988 vss.n5987 9.3005
R10398 vss.n134 vss.n130 9.3005
R10399 vss.n6011 vss.n6010 9.3005
R10400 vss.n2225 vss.n2217 9.15142
R10401 vss.n2446 vss.n2445 9.03579
R10402 vss.n5357 vss.n893 8.95415
R10403 vss.n889 vss.n879 8.95415
R10404 vss.n890 vss.n880 8.95415
R10405 vss.n890 vss.n881 8.95415
R10406 vss.n889 vss.n882 8.95415
R10407 vss.n5354 vss.n893 8.95415
R10408 vss.n4216 vss.n1313 8.65932
R10409 vss.n2521 vss.n2520 8.1562
R10410 vss.n2544 vss.n2543 8.1562
R10411 vss.n773 vss.n752 8.1562
R10412 vss.n5386 vss.n5385 8.1562
R10413 vss.n2218 vss.n2203 7.34399
R10414 vss.n2325 vss.n1308 7.34399
R10415 vss.n3017 vss.n2326 7.34399
R10416 vss.n2398 vss.n2327 7.34399
R10417 vss.n2414 vss.n2382 7.34399
R10418 vss.n1343 vss.n1099 7.16209
R10419 vss.n4206 vss.n1323 7.16209
R10420 vss.n2529 vss.t5 6.79692
R10421 vss.t275 vss.n2621 6.79692
R10422 vss.t273 vss.n2754 6.79692
R10423 vss.n4204 vss.n1325 6.76422
R10424 vss.n5840 vss.n5708 6.21764
R10425 vss.n4286 vss.t9 5.8005
R10426 vss.n4286 vss.t36 5.8005
R10427 vss.n5674 vss.t304 5.8005
R10428 vss.n5674 vss.t24 5.8005
R10429 vss.n5750 vss.t298 5.8005
R10430 vss.n5750 vss.t274 5.8005
R10431 vss.n5733 vss.t301 5.8005
R10432 vss.n5733 vss.t3 5.8005
R10433 vss.n5714 vss.t306 5.8005
R10434 vss.n5714 vss.t268 5.8005
R10435 vss.n5711 vss.t282 5.8005
R10436 vss.n5711 vss.t281 5.8005
R10437 vss.n5694 vss.t308 5.8005
R10438 vss.n5694 vss.t37 5.8005
R10439 vss.n5676 vss.t300 5.8005
R10440 vss.n5676 vss.t1 5.8005
R10441 vss.n5640 vss.t290 5.8005
R10442 vss.n5640 vss.t277 5.8005
R10443 vss.n5625 vss.t314 5.8005
R10444 vss.n5625 vss.t30 5.8005
R10445 vss.n240 vss.t270 5.8005
R10446 vss.n240 vss.t34 5.8005
R10447 vss.n241 vss.t20 5.8005
R10448 vss.n241 vss.t286 5.8005
R10449 vss.n5550 vss.t315 5.8005
R10450 vss.n5550 vss.t289 5.8005
R10451 vss.n5549 vss.t318 5.8005
R10452 vss.n5549 vss.t312 5.8005
R10453 vss.n5548 vss.t22 5.8005
R10454 vss.n5548 vss.t6 5.8005
R10455 vss.n4306 vss.t305 5.8005
R10456 vss.n4306 vss.t311 5.8005
R10457 vss.n4427 vss.t310 5.8005
R10458 vss.n4427 vss.t288 5.8005
R10459 vss.n4437 vss.t279 5.8005
R10460 vss.n4437 vss.t272 5.8005
R10461 vss.n4447 vss.t294 5.8005
R10462 vss.n4447 vss.t313 5.8005
R10463 vss.n4457 vss.t280 5.8005
R10464 vss.n4457 vss.t317 5.8005
R10465 vss.n4467 vss.t292 5.8005
R10466 vss.n4467 vss.t293 5.8005
R10467 vss.n4477 vss.t28 5.8005
R10468 vss.n4477 vss.t276 5.8005
R10469 vss.n4509 vss.t320 5.8005
R10470 vss.n4509 vss.t38 5.8005
R10471 vss.n4519 vss.t316 5.8005
R10472 vss.n4519 vss.t15 5.8005
R10473 vss.n4529 vss.t13 5.8005
R10474 vss.n4529 vss.t11 5.8005
R10475 vss.n4539 vss.t303 5.8005
R10476 vss.n4539 vss.t18 5.8005
R10477 vss.n4549 vss.t26 5.8005
R10478 vss.n4549 vss.t16 5.8005
R10479 vss.n4559 vss.t297 5.8005
R10480 vss.n4559 vss.t295 5.8005
R10481 vss.n2194 vss.n1305 5.57062
R10482 vss.n2419 vss.n2418 5.57062
R10483 vss.n940 vss.n939 5.49286
R10484 vss.n5148 vss.n5147 5.49286
R10485 vss.n908 vss.n907 5.49286
R10486 vss.n1260 vss.n1116 5.49286
R10487 vss.n966 vss.n965 5.49286
R10488 vss.n5145 vss.n5144 5.49286
R10489 vss.n5331 vss.n5330 5.49286
R10490 vss.n1287 vss.n1261 5.49286
R10491 vss.n996 vss.n995 5.49286
R10492 vss.n5143 vss.n5022 5.49286
R10493 vss.n4866 vss.n4865 5.49286
R10494 vss.n4743 vss.n1288 5.49286
R10495 vss.n4238 vss.n4237 5.49286
R10496 vss.n5021 vss.n4235 5.49286
R10497 vss.n4712 vss.n4711 5.49286
R10498 vss.n4589 vss.n1289 5.49286
R10499 vss.n4329 vss.n1290 5.49286
R10500 vss.n2545 vss.n427 5.43763
R10501 vss.n2662 vss.n581 5.43763
R10502 vss.n2664 vss.n2663 5.43763
R10503 vss.n751 vss.n215 5.43763
R10504 vss.n2302 vss.n2231 5.27109
R10505 vss.t7 vss.n2205 5.17276
R10506 vss.n4226 vss.n4225 5.17276
R10507 vss.t283 vss.n2200 5.17276
R10508 vss.n279 vss.n270 4.94293
R10509 vss.n2297 vss.n2236 4.89462
R10510 vss.n3013 vss.n2333 4.89462
R10511 vss.n2286 vss.n2233 4.77489
R10512 vss.n1323 vss.n1087 4.77489
R10513 vss.n2447 vss.n300 4.51815
R10514 vss.n5569 vss.n280 4.5005
R10515 vss.n285 vss.n277 4.5005
R10516 vss.n289 vss.n277 4.5005
R10517 vss.n284 vss.n277 4.5005
R10518 vss.n292 vss.n277 4.5005
R10519 vss.n283 vss.n277 4.5005
R10520 vss.n285 vss.n278 4.5005
R10521 vss.n289 vss.n278 4.5005
R10522 vss.n284 vss.n278 4.5005
R10523 vss.n283 vss.n278 4.5005
R10524 vss.n285 vss.n282 4.5005
R10525 vss.n289 vss.n282 4.5005
R10526 vss.n284 vss.n282 4.5005
R10527 vss.n283 vss.n282 4.5005
R10528 vss.n5569 vss.n278 4.5005
R10529 vss.n5569 vss.n282 4.5005
R10530 vss.n5569 vss.n277 4.5005
R10531 vss.n5569 vss.n5568 4.5005
R10532 vss.n5568 vss.n285 4.5005
R10533 vss.n5568 vss.n289 4.5005
R10534 vss.n5568 vss.n284 4.5005
R10535 vss.n5568 vss.n292 4.5005
R10536 vss.n5568 vss.n283 4.5005
R10537 vss.n5568 vss.n5567 4.5005
R10538 vss.n4378 vss.n4321 4.5005
R10539 vss.n4413 vss.n4312 4.5005
R10540 vss.n4384 vss.n4359 4.5005
R10541 vss.n4385 vss.n4384 4.5005
R10542 vss.n4382 vss.n4321 4.5005
R10543 vss.n4392 vss.n4322 4.5005
R10544 vss.n4212 vss.n1314 4.14168
R10545 vss.n5528 vss.n306 4.07835
R10546 vss.t5 vss.n399 4.07835
R10547 vss.t287 vss.n2544 4.07835
R10548 vss.t31 vss.n539 4.07835
R10549 vss.n2283 vss.n2247 3.97916
R10550 vss.n3021 vss.n3020 3.97916
R10551 vss.n3187 vss.t128 3.86717
R10552 vss.n3187 vss.t199 3.86717
R10553 vss.n3188 vss.t259 3.86717
R10554 vss.n3188 vss.t114 3.86717
R10555 vss.n3099 vss.t98 3.86717
R10556 vss.n3099 vss.t240 3.86717
R10557 vss.n3100 vss.t243 3.86717
R10558 vss.n3100 vss.t170 3.86717
R10559 vss.n3104 vss.t82 3.86717
R10560 vss.n3104 vss.t228 3.86717
R10561 vss.n3105 vss.t229 3.86717
R10562 vss.n3105 vss.t151 3.86717
R10563 vss.n3109 vss.t88 3.86717
R10564 vss.n3109 vss.t233 3.86717
R10565 vss.n3110 vss.t236 3.86717
R10566 vss.n3110 vss.t162 3.86717
R10567 vss.n3115 vss.t70 3.86717
R10568 vss.n3115 vss.t221 3.86717
R10569 vss.n3116 vss.t224 3.86717
R10570 vss.n3116 vss.t144 3.86717
R10571 vss.n3121 vss.t54 3.86717
R10572 vss.n3121 vss.t192 3.86717
R10573 vss.n3122 vss.t211 3.86717
R10574 vss.n3122 vss.t104 3.86717
R10575 vss.n3125 vss.t102 3.86717
R10576 vss.n3125 vss.t149 3.86717
R10577 vss.n3126 vss.t245 3.86717
R10578 vss.n3126 vss.t48 3.86717
R10579 vss.n3132 vss.t44 3.86717
R10580 vss.n3132 vss.t124 3.86717
R10581 vss.n3133 vss.t208 3.86717
R10582 vss.n3133 vss.t257 3.86717
R10583 vss.n3138 vss.t94 3.86717
R10584 vss.n3138 vss.t174 3.86717
R10585 vss.n3139 vss.t239 3.86717
R10586 vss.n3139 vss.t80 3.86717
R10587 vss.n3142 vss.t78 3.86717
R10588 vss.n3142 vss.t153 3.86717
R10589 vss.n3143 vss.t227 3.86717
R10590 vss.n3143 vss.t56 3.86717
R10591 vss.n3149 vss.t253 3.86717
R10592 vss.n3149 vss.t171 3.86717
R10593 vss.n3150 vss.t189 3.86717
R10594 vss.n3150 vss.t72 3.86717
R10595 vss.n3155 vss.t66 3.86717
R10596 vss.n3155 vss.t152 3.86717
R10597 vss.n3156 vss.t220 3.86717
R10598 vss.n3156 vss.t52 3.86717
R10599 vss.n3159 vss.t50 3.86717
R10600 vss.n3159 vss.t126 3.86717
R10601 vss.n3160 vss.t210 3.86717
R10602 vss.n3160 vss.t258 3.86717
R10603 vss.n3166 vss.t175 3.86717
R10604 vss.n3166 vss.t231 3.86717
R10605 vss.n3167 vss.t84 3.86717
R10606 vss.n3167 vss.t158 3.86717
R10607 vss.n3172 vss.t154 3.86717
R10608 vss.n3172 vss.t217 3.86717
R10609 vss.n3173 vss.t58 3.86717
R10610 vss.n3173 vss.t142 3.86717
R10611 vss.n3176 vss.t136 3.86717
R10612 vss.n3176 vss.t247 3.86717
R10613 vss.n3177 vss.t262 3.86717
R10614 vss.n3177 vss.t178 3.86717
R10615 vss.n3183 vss.t176 3.86717
R10616 vss.n3183 vss.t213 3.86717
R10617 vss.n3184 vss.t86 3.86717
R10618 vss.n3184 vss.t132 3.86717
R10619 vss.n3192 vss.t92 3.86717
R10620 vss.n3192 vss.t234 3.86717
R10621 vss.n3193 vss.t237 3.86717
R10622 vss.n3193 vss.t164 3.86717
R10623 vss.n3199 vss.t74 3.86717
R10624 vss.n3199 vss.t222 3.86717
R10625 vss.n3200 vss.t225 3.86717
R10626 vss.n3200 vss.t148 3.86717
R10627 vss.n3203 vss.t251 3.86717
R10628 vss.n3203 vss.t230 3.86717
R10629 vss.n3204 vss.t185 3.86717
R10630 vss.n3204 vss.t156 3.86717
R10631 vss.n3210 vss.t62 3.86717
R10632 vss.n3210 vss.t215 3.86717
R10633 vss.n3211 vss.t218 3.86717
R10634 vss.n3211 vss.t138 3.86717
R10635 vss.n3216 vss.t46 3.86717
R10636 vss.n3216 vss.t205 3.86717
R10637 vss.n3217 vss.t209 3.86717
R10638 vss.n3217 vss.t118 3.86717
R10639 vss.n3220 vss.t96 3.86717
R10640 vss.n3220 vss.t212 3.86717
R10641 vss.n3221 vss.t241 3.86717
R10642 vss.n3221 vss.t130 3.86717
R10643 vss.n3227 vss.t263 3.86717
R10644 vss.n3227 vss.t196 3.86717
R10645 vss.n3228 vss.t201 3.86717
R10646 vss.n3228 vss.t110 3.86717
R10647 vss.n3233 vss.t254 3.86717
R10648 vss.n3233 vss.t232 3.86717
R10649 vss.n3234 vss.t191 3.86717
R10650 vss.n3234 vss.t160 3.86717
R10651 vss.n3237 vss.t68 3.86717
R10652 vss.n3237 vss.t193 3.86717
R10653 vss.n3238 vss.t223 3.86717
R10654 vss.n3238 vss.t108 3.86717
R10655 vss.n3244 vss.t249 3.86717
R10656 vss.n3244 vss.t179 3.86717
R10657 vss.n3245 vss.t183 3.86717
R10658 vss.n3245 vss.t90 3.86717
R10659 vss.n3250 vss.t60 3.86717
R10660 vss.n3250 vss.t214 3.86717
R10661 vss.n3251 vss.t216 3.86717
R10662 vss.n3251 vss.t134 3.86717
R10663 vss.n3254 vss.t266 3.86717
R10664 vss.n3254 vss.t202 3.86717
R10665 vss.n3255 vss.t207 3.86717
R10666 vss.n3255 vss.t116 3.86717
R10667 vss.n3261 vss.t238 3.86717
R10668 vss.n3261 vss.t140 3.86717
R10669 vss.n3262 vss.t168 3.86717
R10670 vss.n3262 vss.t264 3.86717
R10671 vss.n3267 vss.t261 3.86717
R10672 vss.n3267 vss.t120 3.86717
R10673 vss.n3268 vss.t198 3.86717
R10674 vss.n3268 vss.t255 3.86717
R10675 vss.n3271 vss.t252 3.86717
R10676 vss.n3271 vss.t106 3.86717
R10677 vss.n3272 vss.t187 3.86717
R10678 vss.n3272 vss.t246 3.86717
R10679 vss.n3278 vss.t64 3.86717
R10680 vss.n3278 vss.t112 3.86717
R10681 vss.n3279 vss.t219 3.86717
R10682 vss.n3279 vss.t250 3.86717
R10683 vss.n3284 vss.t248 3.86717
R10684 vss.n3284 vss.t100 3.86717
R10685 vss.n3285 vss.t181 3.86717
R10686 vss.n3285 vss.t244 3.86717
R10687 vss.n3288 vss.t242 3.86717
R10688 vss.n3288 vss.t146 3.86717
R10689 vss.n3289 vss.t173 3.86717
R10690 vss.n3289 vss.t267 3.86717
R10691 vss.n3295 vss.t265 3.86717
R10692 vss.n3295 vss.t122 3.86717
R10693 vss.n3296 vss.t204 3.86717
R10694 vss.n3296 vss.t256 3.86717
R10695 vss.n3299 vss.t235 3.86717
R10696 vss.n3299 vss.t76 3.86717
R10697 vss.n3300 vss.t166 3.86717
R10698 vss.n3300 vss.t226 3.86717
R10699 vss.t7 vss.n1293 3.58129
R10700 vss.n3025 vss.n3024 3.58129
R10701 vss.n2979 vss.n1325 3.58129
R10702 vss.n2277 vss.n2261 3.56757
R10703 vss.n2261 vss.t147 3.56757
R10704 vss.n2262 vss.n2250 3.56757
R10705 vss.t147 vss.n2250 3.56757
R10706 vss.n6017 vss.n6016 3.4105
R10707 vss.n6018 vss.n6017 3.4105
R10708 vss.n6014 vss.n95 3.4105
R10709 vss.n6018 vss.n95 3.4105
R10710 vss.n6016 vss.n6015 3.4105
R10711 vss.n6015 vss.n116 3.4105
R10712 vss.n6015 vss.n118 3.4105
R10713 vss.n6015 vss.n115 3.4105
R10714 vss.n6015 vss.n120 3.4105
R10715 vss.n6015 vss.n114 3.4105
R10716 vss.n6015 vss.n122 3.4105
R10717 vss.n6015 vss.n113 3.4105
R10718 vss.n6015 vss.n124 3.4105
R10719 vss.n6015 vss.n112 3.4105
R10720 vss.n6015 vss.n126 3.4105
R10721 vss.n6015 vss.n111 3.4105
R10722 vss.n6015 vss.n128 3.4105
R10723 vss.n6015 vss.n110 3.4105
R10724 vss.n6015 vss.n6014 3.4105
R10725 vss.n2211 vss.n2205 3.18343
R10726 vss.n3006 vss.n2343 3.18343
R10727 vss.n3020 vss.t283 2.78556
R10728 vss.n2542 vss.n413 2.71907
R10729 vss.n2655 vss.n2654 2.71907
R10730 vss.n2665 vss.n595 2.71907
R10731 vss.n775 vss.n774 2.71907
R10732 vss.n2309 vss.n2227 2.3877
R10733 vss.n4227 vss.n1303 2.3877
R10734 vss.n2966 vss.n1075 2.3877
R10735 vss.n2399 vss.n1051 2.3877
R10736 vss.n4352 vss.n4351 2.313
R10737 vss.n4575 vss.n4574 2.313
R10738 vss.n5802 vss.n5801 2.2516
R10739 vss.n5565 vss.n270 2.2505
R10740 vss.n5564 vss.n268 2.2505
R10741 vss.n5563 vss.n266 2.2505
R10742 vss.n5562 vss.n262 2.2505
R10743 vss.n5560 vss.n264 2.2505
R10744 vss.n5559 vss.n258 2.2505
R10745 vss.n5557 vss.n256 2.2505
R10746 vss.n5556 vss.n254 2.2505
R10747 vss.n5555 vss.n252 2.2505
R10748 vss.n5553 vss.n250 2.2505
R10749 vss.n5552 vss.n245 2.2505
R10750 vss.n5551 vss.n246 2.2505
R10751 vss.n5620 vss.n5619 2.2505
R10752 vss.n5621 vss.n228 2.2505
R10753 vss.n5622 vss.n233 2.2505
R10754 vss.n5624 vss.n236 2.2505
R10755 vss.n5902 vss.n5901 2.2505
R10756 vss.n5900 vss.n5899 2.2505
R10757 vss.n5638 vss.n5629 2.2505
R10758 vss.n5639 vss.n5634 2.2505
R10759 vss.n5891 vss.n5890 2.2505
R10760 vss.n5888 vss.n5887 2.2505
R10761 vss.n5644 vss.n5641 2.2505
R10762 vss.n5658 vss.n5651 2.2505
R10763 vss.n5660 vss.n5654 2.2505
R10764 vss.n5875 vss.n5874 2.2505
R10765 vss.n5873 vss.n5872 2.2505
R10766 vss.n5664 vss.n5661 2.2505
R10767 vss.n5675 vss.n5670 2.2505
R10768 vss.n5864 vss.n5863 2.2505
R10769 vss.n5862 vss.n5861 2.2505
R10770 vss.n5695 vss.n5680 2.2505
R10771 vss.n5696 vss.n5687 2.2505
R10772 vss.n5697 vss.n5690 2.2505
R10773 vss.n5849 vss.n5848 2.2505
R10774 vss.n5847 vss.n5846 2.2505
R10775 vss.n5702 vss.n5699 2.2505
R10776 vss.n5713 vss.n5707 2.2505
R10777 vss.n5838 vss.n5837 2.2505
R10778 vss.n5836 vss.n5835 2.2505
R10779 vss.n5734 vss.n5718 2.2505
R10780 vss.n5735 vss.n5726 2.2505
R10781 vss.n5736 vss.n5729 2.2505
R10782 vss.n5823 vss.n5822 2.2505
R10783 vss.n5821 vss.n5820 2.2505
R10784 vss.n5741 vss.n5738 2.2505
R10785 vss.n5752 vss.n5746 2.2505
R10786 vss.n5812 vss.n5811 2.2505
R10787 vss.n5810 vss.n5809 2.2505
R10788 vss.n5759 vss.n5756 2.2505
R10789 vss.n5570 vss.n273 2.2505
R10790 vss.n4353 vss.n4352 2.2505
R10791 vss.n4355 vss.n4326 2.2505
R10792 vss.n4359 vss.n4358 2.2505
R10793 vss.n4386 vss.n4385 2.2505
R10794 vss.n4389 vss.n4321 2.2505
R10795 vss.n4392 vss.n4391 2.2505
R10796 vss.n4395 vss.n4394 2.2505
R10797 vss.n4398 vss.n4397 2.2505
R10798 vss.n4401 vss.n4400 2.2505
R10799 vss.n4406 vss.n4405 2.2505
R10800 vss.n4409 vss.n4408 2.2505
R10801 vss.n4413 vss.n4412 2.2505
R10802 vss.n4415 vss.n4414 2.2505
R10803 vss.n4418 vss.n4310 2.2505
R10804 vss.n4421 vss.n4420 2.2505
R10805 vss.n4423 vss.n4422 2.2505
R10806 vss.n4426 vss.n4425 2.2505
R10807 vss.n4430 vss.n4429 2.2505
R10808 vss.n4432 vss.n4303 2.2505
R10809 vss.n4436 vss.n4435 2.2505
R10810 vss.n4440 vss.n4439 2.2505
R10811 vss.n4443 vss.n4301 2.2505
R10812 vss.n4446 vss.n4445 2.2505
R10813 vss.n4450 vss.n4449 2.2505
R10814 vss.n4452 vss.n4298 2.2505
R10815 vss.n4456 vss.n4455 2.2505
R10816 vss.n4460 vss.n4459 2.2505
R10817 vss.n4463 vss.n4296 2.2505
R10818 vss.n4466 vss.n4465 2.2505
R10819 vss.n4470 vss.n4469 2.2505
R10820 vss.n4472 vss.n4293 2.2505
R10821 vss.n4476 vss.n4475 2.2505
R10822 vss.n4480 vss.n4479 2.2505
R10823 vss.n4483 vss.n4291 2.2505
R10824 vss.n4489 vss.n4488 2.2505
R10825 vss.n4490 vss.n4290 2.2505
R10826 vss.n4494 vss.n4492 2.2505
R10827 vss.n4496 vss.n4289 2.2505
R10828 vss.n4500 vss.n4499 2.2505
R10829 vss.n4502 vss.n4501 2.2505
R10830 vss.n4505 vss.n4287 2.2505
R10831 vss.n4508 vss.n4507 2.2505
R10832 vss.n4512 vss.n4511 2.2505
R10833 vss.n4514 vss.n4283 2.2505
R10834 vss.n4518 vss.n4517 2.2505
R10835 vss.n4522 vss.n4521 2.2505
R10836 vss.n4525 vss.n4281 2.2505
R10837 vss.n4528 vss.n4527 2.2505
R10838 vss.n4532 vss.n4531 2.2505
R10839 vss.n4534 vss.n4278 2.2505
R10840 vss.n4538 vss.n4537 2.2505
R10841 vss.n4542 vss.n4541 2.2505
R10842 vss.n4545 vss.n4276 2.2505
R10843 vss.n4548 vss.n4547 2.2505
R10844 vss.n4552 vss.n4551 2.2505
R10845 vss.n4554 vss.n4273 2.2505
R10846 vss.n4558 vss.n4557 2.2505
R10847 vss.n4562 vss.n4561 2.2505
R10848 vss.n4565 vss.n4271 2.2505
R10849 vss.n4568 vss.n4567 2.2505
R10850 vss.n4570 vss.n4569 2.2505
R10851 vss.n4574 vss.n4573 2.2505
R10852 vss.n292 vss.n290 2.24726
R10853 vss.n5547 vss.n280 2.24718
R10854 vss.n291 vss.n280 2.24718
R10855 vss.n288 vss.n280 2.24718
R10856 vss.n5545 vss.n281 2.24718
R10857 vss.n5545 vss.n294 2.24718
R10858 vss.n5545 vss.n293 2.24718
R10859 vss.n5567 vss.n5566 2.24671
R10860 vss.n5567 vss.n5546 2.24671
R10861 vss.n4361 vss.n4324 2.24547
R10862 vss.n4393 vss.n4312 2.24547
R10863 vss.n4399 vss.n4312 2.24547
R10864 vss.n4407 vss.n4312 2.24547
R10865 vss.n4322 vss.n4318 2.24547
R10866 vss.n4322 vss.n4315 2.24547
R10867 vss.n4322 vss.n4313 2.24547
R10868 vss.n5149 vss.n5148 2.14772
R10869 vss.n939 vss.n938 2.14772
R10870 vss.n1258 vss.n1116 2.14772
R10871 vss.n907 vss.n906 2.14772
R10872 vss.n5144 vss.n1103 2.14772
R10873 vss.n965 vss.n964 2.14772
R10874 vss.n1285 vss.n1261 2.14772
R10875 vss.n5330 vss.n5329 2.14772
R10876 vss.n5141 vss.n5022 2.14772
R10877 vss.n995 vss.n994 2.14772
R10878 vss.n4745 vss.n4743 2.14772
R10879 vss.n4865 vss.n4864 2.14772
R10880 vss.n5019 vss.n4235 2.14772
R10881 vss.n4237 vss.n4236 2.14772
R10882 vss.n4591 vss.n4589 2.14772
R10883 vss.n4711 vss.n4710 2.14772
R10884 vss.n4331 vss.n4329 2.14772
R10885 vss.n2238 vss.n2235 2.08676
R10886 vss.n2226 vss.n2225 1.98983
R10887 vss.t41 vss.n2330 1.98983
R10888 vss.n6013 vss.n109 1.72809
R10889 vss.n106 vss.n98 1.70512
R10890 vss.n6017 vss.n105 1.69691
R10891 vss.n6017 vss.n104 1.69691
R10892 vss.n6017 vss.n103 1.69691
R10893 vss.n6017 vss.n102 1.69691
R10894 vss.n6017 vss.n101 1.69691
R10895 vss.n6017 vss.n100 1.69691
R10896 vss.n127 vss.n95 1.69691
R10897 vss.n125 vss.n95 1.69691
R10898 vss.n121 vss.n95 1.69691
R10899 vss.n119 vss.n95 1.69691
R10900 vss.n117 vss.n95 1.69691
R10901 vss.n107 vss.n95 1.69691
R10902 vss.n6015 vss.n97 1.69691
R10903 vss.n6017 vss.n99 1.6968
R10904 vss.n123 vss.n95 1.6968
R10905 vss.n2274 vss.n2273 1.59196
R10906 vss.n2234 vss.n2216 1.59196
R10907 vss.n4205 vss.n4204 1.59196
R10908 vss.n3601 vss.n3081 1.53201
R10909 vss.n6013 vss.n6012 1.5005
R10910 vss.n3603 vss.n3602 1.5005
R10911 vss.n3082 vss.n3079 1.5005
R10912 vss.n3598 vss.n3074 1.5005
R10913 vss.n3597 vss.n3071 1.5005
R10914 vss.n3596 vss.n3068 1.5005
R10915 vss.n3084 vss.n3065 1.5005
R10916 vss.n3592 vss.n3062 1.5005
R10917 vss.n3591 vss.n3059 1.5005
R10918 vss.n3590 vss.n3056 1.5005
R10919 vss.n3086 vss.n3053 1.5005
R10920 vss.n3586 vss.n3050 1.5005
R10921 vss.n3585 vss.n3047 1.5005
R10922 vss.n3584 vss.n3043 1.5005
R10923 vss.n3088 vss.n3045 1.5005
R10924 vss.n3580 vss.n2186 1.5005
R10925 vss.n3579 vss.n2182 1.5005
R10926 vss.n3578 vss.n2178 1.5005
R10927 vss.n3090 vss.n2174 1.5005
R10928 vss.n3574 vss.n2170 1.5005
R10929 vss.n3573 vss.n2166 1.5005
R10930 vss.n3572 vss.n2162 1.5005
R10931 vss.n3092 vss.n2158 1.5005
R10932 vss.n3568 vss.n2153 1.5005
R10933 vss.n3567 vss.n2155 1.5005
R10934 vss.n3566 vss.n2142 1.5005
R10935 vss.n3094 vss.n2138 1.5005
R10936 vss.n3562 vss.n2134 1.5005
R10937 vss.n3561 vss.n2130 1.5005
R10938 vss.n3560 vss.n2126 1.5005
R10939 vss.n3096 vss.n2122 1.5005
R10940 vss.n3556 vss.n2118 1.5005
R10941 vss.n3555 vss.n2114 1.5005
R10942 vss.n3554 vss.n2110 1.5005
R10943 vss.n3098 vss.n2105 1.5005
R10944 vss.n3549 vss.n2107 1.5005
R10945 vss.n3548 vss.n2084 1.5005
R10946 vss.n3547 vss.n2080 1.5005
R10947 vss.n3103 vss.n2076 1.5005
R10948 vss.n3542 vss.n2072 1.5005
R10949 vss.n3541 vss.n2068 1.5005
R10950 vss.n3540 vss.n2064 1.5005
R10951 vss.n3108 vss.n2060 1.5005
R10952 vss.n3536 vss.n2056 1.5005
R10953 vss.n3535 vss.n2051 1.5005
R10954 vss.n3534 vss.n2053 1.5005
R10955 vss.n3114 vss.n2030 1.5005
R10956 vss.n3530 vss.n2026 1.5005
R10957 vss.n3529 vss.n2022 1.5005
R10958 vss.n3528 vss.n2018 1.5005
R10959 vss.n3120 vss.n2014 1.5005
R10960 vss.n3524 vss.n2010 1.5005
R10961 vss.n3523 vss.n2006 1.5005
R10962 vss.n3129 vss.n2002 1.5005
R10963 vss.n3519 vss.n1997 1.5005
R10964 vss.n3518 vss.n1999 1.5005
R10965 vss.n3517 vss.n1975 1.5005
R10966 vss.n3131 vss.n1971 1.5005
R10967 vss.n3513 vss.n1967 1.5005
R10968 vss.n3512 vss.n1963 1.5005
R10969 vss.n3511 vss.n1959 1.5005
R10970 vss.n3137 vss.n1955 1.5005
R10971 vss.n3507 vss.n1951 1.5005
R10972 vss.n3506 vss.n1947 1.5005
R10973 vss.n3146 vss.n1943 1.5005
R10974 vss.n3502 vss.n1938 1.5005
R10975 vss.n3501 vss.n1940 1.5005
R10976 vss.n3500 vss.n1917 1.5005
R10977 vss.n3148 vss.n1913 1.5005
R10978 vss.n3496 vss.n1909 1.5005
R10979 vss.n3495 vss.n1905 1.5005
R10980 vss.n3494 vss.n1901 1.5005
R10981 vss.n3154 vss.n1897 1.5005
R10982 vss.n3490 vss.n1893 1.5005
R10983 vss.n3489 vss.n1889 1.5005
R10984 vss.n3163 vss.n1884 1.5005
R10985 vss.n3485 vss.n1886 1.5005
R10986 vss.n3484 vss.n1863 1.5005
R10987 vss.n3483 vss.n1859 1.5005
R10988 vss.n3165 vss.n1855 1.5005
R10989 vss.n3479 vss.n1851 1.5005
R10990 vss.n3478 vss.n1847 1.5005
R10991 vss.n3477 vss.n1843 1.5005
R10992 vss.n3171 vss.n1839 1.5005
R10993 vss.n3473 vss.n1835 1.5005
R10994 vss.n3472 vss.n1830 1.5005
R10995 vss.n3180 vss.n1832 1.5005
R10996 vss.n3468 vss.n1808 1.5005
R10997 vss.n3467 vss.n1804 1.5005
R10998 vss.n3466 vss.n1800 1.5005
R10999 vss.n3182 vss.n1796 1.5005
R11000 vss.n3462 vss.n1792 1.5005
R11001 vss.n3461 vss.n1788 1.5005
R11002 vss.n3460 vss.n1784 1.5005
R11003 vss.n3191 vss.n1780 1.5005
R11004 vss.n3456 vss.n1776 1.5005
R11005 vss.n3455 vss.n1771 1.5005
R11006 vss.n3196 vss.n1773 1.5005
R11007 vss.n3451 vss.n1760 1.5005
R11008 vss.n3450 vss.n1756 1.5005
R11009 vss.n3449 vss.n1752 1.5005
R11010 vss.n3198 vss.n1748 1.5005
R11011 vss.n3445 vss.n1744 1.5005
R11012 vss.n3444 vss.n1740 1.5005
R11013 vss.n3207 vss.n1736 1.5005
R11014 vss.n3440 vss.n1732 1.5005
R11015 vss.n3439 vss.n1727 1.5005
R11016 vss.n3438 vss.n1729 1.5005
R11017 vss.n3209 vss.n1705 1.5005
R11018 vss.n3434 vss.n1701 1.5005
R11019 vss.n3433 vss.n1697 1.5005
R11020 vss.n3432 vss.n1693 1.5005
R11021 vss.n3215 vss.n1689 1.5005
R11022 vss.n3428 vss.n1685 1.5005
R11023 vss.n3427 vss.n1681 1.5005
R11024 vss.n3224 vss.n1677 1.5005
R11025 vss.n3423 vss.n1673 1.5005
R11026 vss.n3422 vss.n1668 1.5005
R11027 vss.n3421 vss.n1670 1.5005
R11028 vss.n3226 vss.n1647 1.5005
R11029 vss.n3417 vss.n1643 1.5005
R11030 vss.n3416 vss.n1639 1.5005
R11031 vss.n3415 vss.n1635 1.5005
R11032 vss.n3232 vss.n1631 1.5005
R11033 vss.n3411 vss.n1627 1.5005
R11034 vss.n3410 vss.n1623 1.5005
R11035 vss.n3241 vss.n1619 1.5005
R11036 vss.n3406 vss.n1614 1.5005
R11037 vss.n3405 vss.n1616 1.5005
R11038 vss.n3404 vss.n1593 1.5005
R11039 vss.n3243 vss.n1589 1.5005
R11040 vss.n3400 vss.n1585 1.5005
R11041 vss.n3399 vss.n1581 1.5005
R11042 vss.n3398 vss.n1577 1.5005
R11043 vss.n3249 vss.n1573 1.5005
R11044 vss.n3394 vss.n1569 1.5005
R11045 vss.n3393 vss.n1565 1.5005
R11046 vss.n3258 vss.n1560 1.5005
R11047 vss.n3389 vss.n1562 1.5005
R11048 vss.n3388 vss.n1538 1.5005
R11049 vss.n3387 vss.n1534 1.5005
R11050 vss.n3260 vss.n1530 1.5005
R11051 vss.n3383 vss.n1526 1.5005
R11052 vss.n3382 vss.n1522 1.5005
R11053 vss.n3381 vss.n1518 1.5005
R11054 vss.n3266 vss.n1514 1.5005
R11055 vss.n3377 vss.n1510 1.5005
R11056 vss.n3376 vss.n1506 1.5005
R11057 vss.n3275 vss.n1501 1.5005
R11058 vss.n3372 vss.n1503 1.5005
R11059 vss.n3371 vss.n1480 1.5005
R11060 vss.n3370 vss.n1476 1.5005
R11061 vss.n3277 vss.n1472 1.5005
R11062 vss.n3366 vss.n1468 1.5005
R11063 vss.n3365 vss.n1464 1.5005
R11064 vss.n3364 vss.n1460 1.5005
R11065 vss.n3283 vss.n1456 1.5005
R11066 vss.n3360 vss.n1452 1.5005
R11067 vss.n3359 vss.n1447 1.5005
R11068 vss.n3292 vss.n1449 1.5005
R11069 vss.n3355 vss.n1426 1.5005
R11070 vss.n3354 vss.n1422 1.5005
R11071 vss.n3353 vss.n1418 1.5005
R11072 vss.n3294 vss.n1414 1.5005
R11073 vss.n3349 vss.n1410 1.5005
R11074 vss.n3348 vss.n1406 1.5005
R11075 vss.n3303 vss.n1402 1.5005
R11076 vss.n3344 vss.n1398 1.5005
R11077 vss.n3343 vss.n1393 1.5005
R11078 vss.n3342 vss.n1395 1.5005
R11079 vss.n3305 vss.n1382 1.5005
R11080 vss.n3338 vss.n1378 1.5005
R11081 vss.n3337 vss.n1374 1.5005
R11082 vss.n3336 vss.n1370 1.5005
R11083 vss.n3309 vss.n1366 1.5005
R11084 vss.n3330 vss.n1362 1.5005
R11085 vss.n3329 vss.n1358 1.5005
R11086 vss.n3328 vss.n1355 1.5005
R11087 vss.n3313 vss.n1351 1.5005
R11088 vss.n3321 vss.n1346 1.5005
R11089 vss.n3320 vss.n1348 1.5005
R11090 vss.n3317 vss.n1333 1.5005
R11091 vss.n4200 vss.n3 1.5005
R11092 vss.n6127 vss.n4 1.5005
R11093 vss.n6126 vss.n5 1.5005
R11094 vss.n6125 vss.n6 1.5005
R11095 vss.n3002 vss.n7 1.5005
R11096 vss.n6121 vss.n9 1.5005
R11097 vss.n6120 vss.n10 1.5005
R11098 vss.n6119 vss.n11 1.5005
R11099 vss.n2954 vss.n12 1.5005
R11100 vss.n6115 vss.n14 1.5005
R11101 vss.n6114 vss.n15 1.5005
R11102 vss.n6113 vss.n16 1.5005
R11103 vss.n2465 vss.n17 1.5005
R11104 vss.n6109 vss.n19 1.5005
R11105 vss.n6108 vss.n20 1.5005
R11106 vss.n6107 vss.n21 1.5005
R11107 vss.n2480 vss.n22 1.5005
R11108 vss.n6103 vss.n24 1.5005
R11109 vss.n6102 vss.n25 1.5005
R11110 vss.n6101 vss.n26 1.5005
R11111 vss.n2506 vss.n27 1.5005
R11112 vss.n6097 vss.n29 1.5005
R11113 vss.n6096 vss.n30 1.5005
R11114 vss.n6095 vss.n31 1.5005
R11115 vss.n2905 vss.n32 1.5005
R11116 vss.n6091 vss.n34 1.5005
R11117 vss.n6090 vss.n35 1.5005
R11118 vss.n6089 vss.n36 1.5005
R11119 vss.n2541 vss.n37 1.5005
R11120 vss.n6085 vss.n39 1.5005
R11121 vss.n6084 vss.n40 1.5005
R11122 vss.n6083 vss.n41 1.5005
R11123 vss.n2881 vss.n42 1.5005
R11124 vss.n6079 vss.n44 1.5005
R11125 vss.n6078 vss.n45 1.5005
R11126 vss.n6077 vss.n46 1.5005
R11127 vss.n2587 vss.n47 1.5005
R11128 vss.n6073 vss.n49 1.5005
R11129 vss.n6072 vss.n50 1.5005
R11130 vss.n6071 vss.n51 1.5005
R11131 vss.n2613 vss.n52 1.5005
R11132 vss.n6067 vss.n54 1.5005
R11133 vss.n6066 vss.n55 1.5005
R11134 vss.n6065 vss.n56 1.5005
R11135 vss.n2630 vss.n57 1.5005
R11136 vss.n6061 vss.n59 1.5005
R11137 vss.n6060 vss.n60 1.5005
R11138 vss.n6059 vss.n61 1.5005
R11139 vss.n2833 vss.n62 1.5005
R11140 vss.n6055 vss.n64 1.5005
R11141 vss.n6054 vss.n65 1.5005
R11142 vss.n6053 vss.n66 1.5005
R11143 vss.n2821 vss.n67 1.5005
R11144 vss.n6049 vss.n69 1.5005
R11145 vss.n6048 vss.n70 1.5005
R11146 vss.n6047 vss.n71 1.5005
R11147 vss.n2695 vss.n72 1.5005
R11148 vss.n6043 vss.n74 1.5005
R11149 vss.n6042 vss.n75 1.5005
R11150 vss.n6041 vss.n76 1.5005
R11151 vss.n2714 vss.n77 1.5005
R11152 vss.n6037 vss.n79 1.5005
R11153 vss.n6036 vss.n80 1.5005
R11154 vss.n6035 vss.n81 1.5005
R11155 vss.n2741 vss.n82 1.5005
R11156 vss.n6031 vss.n84 1.5005
R11157 vss.n6030 vss.n85 1.5005
R11158 vss.n6029 vss.n86 1.5005
R11159 vss.n2760 vss.n87 1.5005
R11160 vss.n6025 vss.n89 1.5005
R11161 vss.n6024 vss.n90 1.5005
R11162 vss.n6023 vss.n91 1.5005
R11163 vss.n201 vss.n92 1.5005
R11164 vss.n6019 vss.n94 1.5005
R11165 vss.n6018 vss.n96 1.5005
R11166 vss.n191 vss.n106 1.5005
R11167 vss.n6016 vss.n108 1.5005
R11168 vss.n184 vss.n116 1.5005
R11169 vss.n180 vss.n118 1.5005
R11170 vss.n176 vss.n115 1.5005
R11171 vss.n171 vss.n120 1.5005
R11172 vss.n172 vss.n114 1.5005
R11173 vss.n159 vss.n122 1.5005
R11174 vss.n154 vss.n113 1.5005
R11175 vss.n5967 vss.n124 1.5005
R11176 vss.n5999 vss.n112 1.5005
R11177 vss.n5969 vss.n126 1.5005
R11178 vss.n5974 vss.n111 1.5005
R11179 vss.n5991 vss.n128 1.5005
R11180 vss.n5980 vss.n110 1.5005
R11181 vss.n6014 vss.n129 1.5005
R11182 vss.t23 vss.n581 1.35978
R11183 vss.n2679 vss.t0 1.35978
R11184 vss.n4225 vss.n1305 1.1941
R11185 vss.n3025 vss.n1343 1.1941
R11186 vss.n2417 vss.t42 1.1941
R11187 vss.n3334 vss.n3333 1.15283
R11188 vss.n6130 vss.n6129 1.15283
R11189 vss.n6126 vss.n2 1.13717
R11190 vss.n6125 vss.n6124 1.13717
R11191 vss.n6123 vss.n7 1.13717
R11192 vss.n6122 vss.n6121 1.13717
R11193 vss.n6120 vss.n8 1.13717
R11194 vss.n6119 vss.n6118 1.13717
R11195 vss.n6117 vss.n12 1.13717
R11196 vss.n6116 vss.n6115 1.13717
R11197 vss.n6114 vss.n13 1.13717
R11198 vss.n6113 vss.n6112 1.13717
R11199 vss.n6111 vss.n17 1.13717
R11200 vss.n6110 vss.n6109 1.13717
R11201 vss.n6108 vss.n18 1.13717
R11202 vss.n6107 vss.n6106 1.13717
R11203 vss.n6105 vss.n22 1.13717
R11204 vss.n6104 vss.n6103 1.13717
R11205 vss.n6102 vss.n23 1.13717
R11206 vss.n6101 vss.n6100 1.13717
R11207 vss.n6099 vss.n27 1.13717
R11208 vss.n6098 vss.n6097 1.13717
R11209 vss.n6096 vss.n28 1.13717
R11210 vss.n6095 vss.n6094 1.13717
R11211 vss.n6093 vss.n32 1.13717
R11212 vss.n6092 vss.n6091 1.13717
R11213 vss.n6090 vss.n33 1.13717
R11214 vss.n6089 vss.n6088 1.13717
R11215 vss.n6087 vss.n37 1.13717
R11216 vss.n6086 vss.n6085 1.13717
R11217 vss.n6084 vss.n38 1.13717
R11218 vss.n6083 vss.n6082 1.13717
R11219 vss.n6081 vss.n42 1.13717
R11220 vss.n6080 vss.n6079 1.13717
R11221 vss.n6078 vss.n43 1.13717
R11222 vss.n6077 vss.n6076 1.13717
R11223 vss.n6075 vss.n47 1.13717
R11224 vss.n6074 vss.n6073 1.13717
R11225 vss.n6072 vss.n48 1.13717
R11226 vss.n6071 vss.n6070 1.13717
R11227 vss.n6069 vss.n52 1.13717
R11228 vss.n6068 vss.n6067 1.13717
R11229 vss.n6066 vss.n53 1.13717
R11230 vss.n6065 vss.n6064 1.13717
R11231 vss.n6063 vss.n57 1.13717
R11232 vss.n6062 vss.n6061 1.13717
R11233 vss.n6060 vss.n58 1.13717
R11234 vss.n6059 vss.n6058 1.13717
R11235 vss.n6057 vss.n62 1.13717
R11236 vss.n6056 vss.n6055 1.13717
R11237 vss.n6054 vss.n63 1.13717
R11238 vss.n6053 vss.n6052 1.13717
R11239 vss.n6051 vss.n67 1.13717
R11240 vss.n6050 vss.n6049 1.13717
R11241 vss.n6048 vss.n68 1.13717
R11242 vss.n6047 vss.n6046 1.13717
R11243 vss.n6045 vss.n72 1.13717
R11244 vss.n6044 vss.n6043 1.13717
R11245 vss.n6042 vss.n73 1.13717
R11246 vss.n6041 vss.n6040 1.13717
R11247 vss.n6039 vss.n77 1.13717
R11248 vss.n6038 vss.n6037 1.13717
R11249 vss.n6036 vss.n78 1.13717
R11250 vss.n6035 vss.n6034 1.13717
R11251 vss.n6033 vss.n82 1.13717
R11252 vss.n6032 vss.n6031 1.13717
R11253 vss.n6030 vss.n83 1.13717
R11254 vss.n6029 vss.n6028 1.13717
R11255 vss.n6027 vss.n87 1.13717
R11256 vss.n6026 vss.n6025 1.13717
R11257 vss.n6024 vss.n88 1.13717
R11258 vss.n6023 vss.n6022 1.13717
R11259 vss.n6021 vss.n92 1.13717
R11260 vss.n6020 vss.n6019 1.13717
R11261 vss.n3337 vss.n3308 1.13717
R11262 vss.n3600 vss.n3082 1.13717
R11263 vss.n3599 vss.n3598 1.13717
R11264 vss.n3597 vss.n3083 1.13717
R11265 vss.n3596 vss.n3595 1.13717
R11266 vss.n3594 vss.n3084 1.13717
R11267 vss.n3593 vss.n3592 1.13717
R11268 vss.n3591 vss.n3085 1.13717
R11269 vss.n3590 vss.n3589 1.13717
R11270 vss.n3588 vss.n3086 1.13717
R11271 vss.n3587 vss.n3586 1.13717
R11272 vss.n3585 vss.n3087 1.13717
R11273 vss.n3584 vss.n3583 1.13717
R11274 vss.n3582 vss.n3088 1.13717
R11275 vss.n3581 vss.n3580 1.13717
R11276 vss.n3579 vss.n3089 1.13717
R11277 vss.n3578 vss.n3577 1.13717
R11278 vss.n3576 vss.n3090 1.13717
R11279 vss.n3575 vss.n3574 1.13717
R11280 vss.n3573 vss.n3091 1.13717
R11281 vss.n3572 vss.n3571 1.13717
R11282 vss.n3570 vss.n3092 1.13717
R11283 vss.n3569 vss.n3568 1.13717
R11284 vss.n3567 vss.n3093 1.13717
R11285 vss.n3566 vss.n3565 1.13717
R11286 vss.n3564 vss.n3094 1.13717
R11287 vss.n3563 vss.n3562 1.13717
R11288 vss.n3561 vss.n3095 1.13717
R11289 vss.n3560 vss.n3559 1.13717
R11290 vss.n3558 vss.n3096 1.13717
R11291 vss.n3557 vss.n3556 1.13717
R11292 vss.n3555 vss.n3097 1.13717
R11293 vss.n3554 vss.n3553 1.13717
R11294 vss.n3551 vss.n3098 1.13717
R11295 vss.n3550 vss.n3549 1.13717
R11296 vss.n3548 vss.n3102 1.13717
R11297 vss.n3547 vss.n3546 1.13717
R11298 vss.n3544 vss.n3103 1.13717
R11299 vss.n3543 vss.n3542 1.13717
R11300 vss.n3541 vss.n3107 1.13717
R11301 vss.n3540 vss.n3539 1.13717
R11302 vss.n3538 vss.n3108 1.13717
R11303 vss.n3537 vss.n3536 1.13717
R11304 vss.n3535 vss.n3113 1.13717
R11305 vss.n3534 vss.n3533 1.13717
R11306 vss.n3532 vss.n3114 1.13717
R11307 vss.n3531 vss.n3530 1.13717
R11308 vss.n3529 vss.n3119 1.13717
R11309 vss.n3528 vss.n3527 1.13717
R11310 vss.n3526 vss.n3120 1.13717
R11311 vss.n3525 vss.n3524 1.13717
R11312 vss.n3523 vss.n3522 1.13717
R11313 vss.n3521 vss.n3129 1.13717
R11314 vss.n3520 vss.n3519 1.13717
R11315 vss.n3518 vss.n3130 1.13717
R11316 vss.n3517 vss.n3516 1.13717
R11317 vss.n3515 vss.n3131 1.13717
R11318 vss.n3514 vss.n3513 1.13717
R11319 vss.n3512 vss.n3136 1.13717
R11320 vss.n3511 vss.n3510 1.13717
R11321 vss.n3509 vss.n3137 1.13717
R11322 vss.n3508 vss.n3507 1.13717
R11323 vss.n3506 vss.n3505 1.13717
R11324 vss.n3504 vss.n3146 1.13717
R11325 vss.n3503 vss.n3502 1.13717
R11326 vss.n3501 vss.n3147 1.13717
R11327 vss.n3500 vss.n3499 1.13717
R11328 vss.n3498 vss.n3148 1.13717
R11329 vss.n3497 vss.n3496 1.13717
R11330 vss.n3495 vss.n3153 1.13717
R11331 vss.n3494 vss.n3493 1.13717
R11332 vss.n3492 vss.n3154 1.13717
R11333 vss.n3491 vss.n3490 1.13717
R11334 vss.n3489 vss.n3488 1.13717
R11335 vss.n3487 vss.n3163 1.13717
R11336 vss.n3486 vss.n3485 1.13717
R11337 vss.n3484 vss.n3164 1.13717
R11338 vss.n3483 vss.n3482 1.13717
R11339 vss.n3481 vss.n3165 1.13717
R11340 vss.n3480 vss.n3479 1.13717
R11341 vss.n3478 vss.n3170 1.13717
R11342 vss.n3477 vss.n3476 1.13717
R11343 vss.n3475 vss.n3171 1.13717
R11344 vss.n3474 vss.n3473 1.13717
R11345 vss.n3472 vss.n3471 1.13717
R11346 vss.n3470 vss.n3180 1.13717
R11347 vss.n3469 vss.n3468 1.13717
R11348 vss.n3467 vss.n3181 1.13717
R11349 vss.n3466 vss.n3465 1.13717
R11350 vss.n3464 vss.n3182 1.13717
R11351 vss.n3463 vss.n3462 1.13717
R11352 vss.n3461 vss.n3190 1.13717
R11353 vss.n3460 vss.n3459 1.13717
R11354 vss.n3458 vss.n3191 1.13717
R11355 vss.n3457 vss.n3456 1.13717
R11356 vss.n3455 vss.n3454 1.13717
R11357 vss.n3453 vss.n3196 1.13717
R11358 vss.n3452 vss.n3451 1.13717
R11359 vss.n3450 vss.n3197 1.13717
R11360 vss.n3449 vss.n3448 1.13717
R11361 vss.n3447 vss.n3198 1.13717
R11362 vss.n3446 vss.n3445 1.13717
R11363 vss.n3444 vss.n3443 1.13717
R11364 vss.n3442 vss.n3207 1.13717
R11365 vss.n3441 vss.n3440 1.13717
R11366 vss.n3439 vss.n3208 1.13717
R11367 vss.n3438 vss.n3437 1.13717
R11368 vss.n3436 vss.n3209 1.13717
R11369 vss.n3435 vss.n3434 1.13717
R11370 vss.n3433 vss.n3214 1.13717
R11371 vss.n3432 vss.n3431 1.13717
R11372 vss.n3430 vss.n3215 1.13717
R11373 vss.n3429 vss.n3428 1.13717
R11374 vss.n3427 vss.n3426 1.13717
R11375 vss.n3425 vss.n3224 1.13717
R11376 vss.n3424 vss.n3423 1.13717
R11377 vss.n3422 vss.n3225 1.13717
R11378 vss.n3421 vss.n3420 1.13717
R11379 vss.n3419 vss.n3226 1.13717
R11380 vss.n3418 vss.n3417 1.13717
R11381 vss.n3416 vss.n3231 1.13717
R11382 vss.n3415 vss.n3414 1.13717
R11383 vss.n3413 vss.n3232 1.13717
R11384 vss.n3412 vss.n3411 1.13717
R11385 vss.n3410 vss.n3409 1.13717
R11386 vss.n3408 vss.n3241 1.13717
R11387 vss.n3407 vss.n3406 1.13717
R11388 vss.n3405 vss.n3242 1.13717
R11389 vss.n3404 vss.n3403 1.13717
R11390 vss.n3402 vss.n3243 1.13717
R11391 vss.n3401 vss.n3400 1.13717
R11392 vss.n3399 vss.n3248 1.13717
R11393 vss.n3398 vss.n3397 1.13717
R11394 vss.n3396 vss.n3249 1.13717
R11395 vss.n3395 vss.n3394 1.13717
R11396 vss.n3393 vss.n3392 1.13717
R11397 vss.n3391 vss.n3258 1.13717
R11398 vss.n3390 vss.n3389 1.13717
R11399 vss.n3388 vss.n3259 1.13717
R11400 vss.n3387 vss.n3386 1.13717
R11401 vss.n3385 vss.n3260 1.13717
R11402 vss.n3384 vss.n3383 1.13717
R11403 vss.n3382 vss.n3265 1.13717
R11404 vss.n3381 vss.n3380 1.13717
R11405 vss.n3379 vss.n3266 1.13717
R11406 vss.n3378 vss.n3377 1.13717
R11407 vss.n3376 vss.n3375 1.13717
R11408 vss.n3374 vss.n3275 1.13717
R11409 vss.n3373 vss.n3372 1.13717
R11410 vss.n3371 vss.n3276 1.13717
R11411 vss.n3370 vss.n3369 1.13717
R11412 vss.n3368 vss.n3277 1.13717
R11413 vss.n3367 vss.n3366 1.13717
R11414 vss.n3365 vss.n3282 1.13717
R11415 vss.n3364 vss.n3363 1.13717
R11416 vss.n3362 vss.n3283 1.13717
R11417 vss.n3361 vss.n3360 1.13717
R11418 vss.n3359 vss.n3358 1.13717
R11419 vss.n3357 vss.n3292 1.13717
R11420 vss.n3356 vss.n3355 1.13717
R11421 vss.n3354 vss.n3293 1.13717
R11422 vss.n3353 vss.n3352 1.13717
R11423 vss.n3351 vss.n3294 1.13717
R11424 vss.n3350 vss.n3349 1.13717
R11425 vss.n3348 vss.n3347 1.13717
R11426 vss.n3346 vss.n3303 1.13717
R11427 vss.n3345 vss.n3344 1.13717
R11428 vss.n3343 vss.n3304 1.13717
R11429 vss.n3342 vss.n3341 1.13717
R11430 vss.n3340 vss.n3305 1.13717
R11431 vss.n3339 vss.n3338 1.13717
R11432 vss.n3336 vss.n3335 1.13717
R11433 vss.n3310 vss.n3309 1.13717
R11434 vss.n3331 vss.n3330 1.13717
R11435 vss.n3329 vss.n3312 1.13717
R11436 vss.n3328 vss.n3327 1.13717
R11437 vss.n3315 vss.n3313 1.13717
R11438 vss.n3322 vss.n3321 1.13717
R11439 vss.n3320 vss.n3319 1.13717
R11440 vss.n3318 vss.n3317 1.13717
R11441 vss.n3333 vss.n3332 1.13717
R11442 vss.n3314 vss.n3311 1.13717
R11443 vss.n3326 vss.n3325 1.13717
R11444 vss.n3324 vss.n3323 1.13717
R11445 vss.n3316 vss.n1 1.13717
R11446 vss.n6131 vss.n6130 1.13717
R11447 vss.n3 vss.n0 1.13717
R11448 vss.n6128 vss.n6127 1.13717
R11449 vss.n4584 vss.n4583 0.877959
R11450 vss.n2280 vss.n2249 0.796232
R11451 vss.n2217 vss.n1291 0.796232
R11452 vss.n2990 vss.n2329 0.796232
R11453 vss.n2298 vss.n2235 0.774431
R11454 vss.n5571 vss.n5570 0.620831
R11455 vss.n5541 vss.n298 0.615535
R11456 vss.n3601 vss.n3600 0.57778
R11457 vss.n3190 vss.n3189 0.549658
R11458 vss.n3552 vss.n3101 0.549658
R11459 vss.n3545 vss.n3106 0.549658
R11460 vss.n3112 vss.n3111 0.549658
R11461 vss.n3118 vss.n3117 0.549658
R11462 vss.n3124 vss.n3123 0.549658
R11463 vss.n3128 vss.n3127 0.549658
R11464 vss.n3135 vss.n3134 0.549658
R11465 vss.n3141 vss.n3140 0.549658
R11466 vss.n3145 vss.n3144 0.549658
R11467 vss.n3152 vss.n3151 0.549658
R11468 vss.n3158 vss.n3157 0.549658
R11469 vss.n3162 vss.n3161 0.549658
R11470 vss.n3169 vss.n3168 0.549658
R11471 vss.n3175 vss.n3174 0.549658
R11472 vss.n3179 vss.n3178 0.549658
R11473 vss.n3186 vss.n3185 0.549658
R11474 vss.n3195 vss.n3194 0.549658
R11475 vss.n3202 vss.n3201 0.549658
R11476 vss.n3206 vss.n3205 0.549658
R11477 vss.n3213 vss.n3212 0.549658
R11478 vss.n3219 vss.n3218 0.549658
R11479 vss.n3223 vss.n3222 0.549658
R11480 vss.n3230 vss.n3229 0.549658
R11481 vss.n3236 vss.n3235 0.549658
R11482 vss.n3240 vss.n3239 0.549658
R11483 vss.n3247 vss.n3246 0.549658
R11484 vss.n3253 vss.n3252 0.549658
R11485 vss.n3257 vss.n3256 0.549658
R11486 vss.n3264 vss.n3263 0.549658
R11487 vss.n3270 vss.n3269 0.549658
R11488 vss.n3274 vss.n3273 0.549658
R11489 vss.n3281 vss.n3280 0.549658
R11490 vss.n3287 vss.n3286 0.549658
R11491 vss.n3291 vss.n3290 0.549658
R11492 vss.n3298 vss.n3297 0.549658
R11493 vss.n3302 vss.n3301 0.549658
R11494 vss.n3307 vss.n3306 0.549658
R11495 vss.n2401 vss.n2400 0.398366
R11496 vss.n2974 vss.n1316 0.376971
R11497 vss.n2221 vss.n2218 0.347881
R11498 vss.n4221 vss.n1308 0.347881
R11499 vss.n2969 vss.n2326 0.347881
R11500 vss.n2398 vss.n2397 0.347881
R11501 vss.n2439 vss.n2382 0.347881
R11502 vss.n5532 vss.n5531 0.347881
R11503 vss.n2239 vss.n2237 0.306952
R11504 vss.n2296 vss.n2295 0.294855
R11505 vss.n2295 vss.n2237 0.294855
R11506 vss.n5795 vss.n5762 0.265206
R11507 vss.n5794 vss.n5793 0.265206
R11508 vss.n5764 vss.n5763 0.265206
R11509 vss.n5789 vss.n5767 0.265206
R11510 vss.n5788 vss.n5768 0.265206
R11511 vss.n5787 vss.n5769 0.265206
R11512 vss.n5772 vss.n5770 0.265206
R11513 vss.n5783 vss.n5773 0.265206
R11514 vss.n5782 vss.n5774 0.265206
R11515 vss.n5781 vss.n5775 0.265206
R11516 vss.n5797 vss.n5796 0.265206
R11517 vss.n5533 vss.n301 0.249932
R11518 vss.n5801 vss.n5800 0.236488
R11519 vss.n5150 vss.n1091 0.223326
R11520 vss.n5161 vss.n5160 0.223326
R11521 vss.n5162 vss.n1067 0.223326
R11522 vss.n5173 vss.n5172 0.223326
R11523 vss.n5174 vss.n1043 0.223326
R11524 vss.n5185 vss.n5184 0.223326
R11525 vss.n5186 vss.n1019 0.223326
R11526 vss.n5204 vss.n5203 0.223326
R11527 vss.n5206 vss.n5205 0.223326
R11528 vss.n320 vss.n319 0.223326
R11529 vss.n346 vss.n321 0.223326
R11530 vss.n348 vss.n347 0.223326
R11531 vss.n374 vss.n349 0.223326
R11532 vss.n376 vss.n375 0.223326
R11533 vss.n402 vss.n377 0.223326
R11534 vss.n404 vss.n403 0.223326
R11535 vss.n430 vss.n405 0.223326
R11536 vss.n432 vss.n431 0.223326
R11537 vss.n458 vss.n433 0.223326
R11538 vss.n460 vss.n459 0.223326
R11539 vss.n486 vss.n461 0.223326
R11540 vss.n488 vss.n487 0.223326
R11541 vss.n514 vss.n489 0.223326
R11542 vss.n516 vss.n515 0.223326
R11543 vss.n542 vss.n517 0.223326
R11544 vss.n544 vss.n543 0.223326
R11545 vss.n570 vss.n545 0.223326
R11546 vss.n572 vss.n571 0.223326
R11547 vss.n598 vss.n573 0.223326
R11548 vss.n600 vss.n599 0.223326
R11549 vss.n626 vss.n601 0.223326
R11550 vss.n628 vss.n627 0.223326
R11551 vss.n654 vss.n629 0.223326
R11552 vss.n656 vss.n655 0.223326
R11553 vss.n682 vss.n657 0.223326
R11554 vss.n684 vss.n683 0.223326
R11555 vss.n710 vss.n685 0.223326
R11556 vss.n712 vss.n711 0.223326
R11557 vss.n737 vss.n713 0.223326
R11558 vss.n739 vss.n738 0.223326
R11559 vss.n915 vss.n913 0.223326
R11560 vss.n918 vss.n916 0.223326
R11561 vss.n921 vss.n919 0.223326
R11562 vss.n924 vss.n922 0.223326
R11563 vss.n927 vss.n925 0.223326
R11564 vss.n930 vss.n928 0.223326
R11565 vss.n933 vss.n931 0.223326
R11566 vss.n935 vss.n934 0.223326
R11567 vss.n937 vss.n936 0.223326
R11568 vss.n1257 vss.n1256 0.223326
R11569 vss.n1254 vss.n1253 0.223326
R11570 vss.n1251 vss.n1250 0.223326
R11571 vss.n1248 vss.n1247 0.223326
R11572 vss.n1245 vss.n1244 0.223326
R11573 vss.n1242 vss.n1241 0.223326
R11574 vss.n1239 vss.n1238 0.223326
R11575 vss.n1236 vss.n1235 0.223326
R11576 vss.n1233 vss.n1232 0.223326
R11577 vss.n1230 vss.n1229 0.223326
R11578 vss.n1227 vss.n1226 0.223326
R11579 vss.n1224 vss.n1223 0.223326
R11580 vss.n1221 vss.n1220 0.223326
R11581 vss.n1218 vss.n1217 0.223326
R11582 vss.n1215 vss.n1214 0.223326
R11583 vss.n1212 vss.n1211 0.223326
R11584 vss.n1209 vss.n1208 0.223326
R11585 vss.n1206 vss.n1205 0.223326
R11586 vss.n1203 vss.n1202 0.223326
R11587 vss.n1200 vss.n1199 0.223326
R11588 vss.n1197 vss.n1196 0.223326
R11589 vss.n1194 vss.n1193 0.223326
R11590 vss.n1191 vss.n1190 0.223326
R11591 vss.n1188 vss.n1187 0.223326
R11592 vss.n1185 vss.n1184 0.223326
R11593 vss.n1182 vss.n1181 0.223326
R11594 vss.n1179 vss.n1178 0.223326
R11595 vss.n1176 vss.n1175 0.223326
R11596 vss.n1173 vss.n1172 0.223326
R11597 vss.n1170 vss.n1169 0.223326
R11598 vss.n1167 vss.n1166 0.223326
R11599 vss.n1164 vss.n1163 0.223326
R11600 vss.n1161 vss.n1160 0.223326
R11601 vss.n1158 vss.n1157 0.223326
R11602 vss.n1155 vss.n1154 0.223326
R11603 vss.n1152 vss.n1151 0.223326
R11604 vss.n1149 vss.n1148 0.223326
R11605 vss.n1146 vss.n1145 0.223326
R11606 vss.n1143 vss.n1142 0.223326
R11607 vss.n1140 vss.n1139 0.223326
R11608 vss.n1138 vss.n1137 0.223326
R11609 vss.n1135 vss.n1134 0.223326
R11610 vss.n1132 vss.n1131 0.223326
R11611 vss.n1129 vss.n1128 0.223326
R11612 vss.n1126 vss.n1125 0.223326
R11613 vss.n1123 vss.n1122 0.223326
R11614 vss.n1120 vss.n1119 0.223326
R11615 vss.n1117 vss.n903 0.223326
R11616 vss.n905 vss.n904 0.223326
R11617 vss.n5155 vss.n5154 0.223326
R11618 vss.n5156 vss.n1079 0.223326
R11619 vss.n5167 vss.n5166 0.223326
R11620 vss.n5168 vss.n1055 0.223326
R11621 vss.n5179 vss.n5178 0.223326
R11622 vss.n5180 vss.n1031 0.223326
R11623 vss.n5191 vss.n5190 0.223326
R11624 vss.n5198 vss.n5192 0.223326
R11625 vss.n5197 vss.n5196 0.223326
R11626 vss.n5194 vss.n5193 0.223326
R11627 vss.n334 vss.n333 0.223326
R11628 vss.n360 vss.n335 0.223326
R11629 vss.n362 vss.n361 0.223326
R11630 vss.n388 vss.n363 0.223326
R11631 vss.n390 vss.n389 0.223326
R11632 vss.n416 vss.n391 0.223326
R11633 vss.n418 vss.n417 0.223326
R11634 vss.n444 vss.n419 0.223326
R11635 vss.n446 vss.n445 0.223326
R11636 vss.n472 vss.n447 0.223326
R11637 vss.n474 vss.n473 0.223326
R11638 vss.n500 vss.n475 0.223326
R11639 vss.n502 vss.n501 0.223326
R11640 vss.n528 vss.n503 0.223326
R11641 vss.n530 vss.n529 0.223326
R11642 vss.n556 vss.n531 0.223326
R11643 vss.n558 vss.n557 0.223326
R11644 vss.n584 vss.n559 0.223326
R11645 vss.n586 vss.n585 0.223326
R11646 vss.n612 vss.n587 0.223326
R11647 vss.n614 vss.n613 0.223326
R11648 vss.n640 vss.n615 0.223326
R11649 vss.n642 vss.n641 0.223326
R11650 vss.n668 vss.n643 0.223326
R11651 vss.n670 vss.n669 0.223326
R11652 vss.n696 vss.n671 0.223326
R11653 vss.n698 vss.n697 0.223326
R11654 vss.n724 vss.n699 0.223326
R11655 vss.n726 vss.n725 0.223326
R11656 vss.n757 vss.n727 0.223326
R11657 vss.n759 vss.n758 0.223326
R11658 vss.n944 vss.n760 0.223326
R11659 vss.n947 vss.n945 0.223326
R11660 vss.n950 vss.n948 0.223326
R11661 vss.n953 vss.n951 0.223326
R11662 vss.n956 vss.n954 0.223326
R11663 vss.n959 vss.n957 0.223326
R11664 vss.n961 vss.n960 0.223326
R11665 vss.n963 vss.n962 0.223326
R11666 vss.n1284 vss.n1283 0.223326
R11667 vss.n1281 vss.n1280 0.223326
R11668 vss.n1278 vss.n1277 0.223326
R11669 vss.n1275 vss.n1274 0.223326
R11670 vss.n1272 vss.n1271 0.223326
R11671 vss.n1269 vss.n1268 0.223326
R11672 vss.n1266 vss.n1265 0.223326
R11673 vss.n1263 vss.n1262 0.223326
R11674 vss.n5211 vss.n1007 0.223326
R11675 vss.n5214 vss.n5212 0.223326
R11676 vss.n5217 vss.n5215 0.223326
R11677 vss.n5220 vss.n5218 0.223326
R11678 vss.n5223 vss.n5221 0.223326
R11679 vss.n5226 vss.n5224 0.223326
R11680 vss.n5229 vss.n5227 0.223326
R11681 vss.n5232 vss.n5230 0.223326
R11682 vss.n5235 vss.n5233 0.223326
R11683 vss.n5238 vss.n5236 0.223326
R11684 vss.n5241 vss.n5239 0.223326
R11685 vss.n5244 vss.n5242 0.223326
R11686 vss.n5247 vss.n5245 0.223326
R11687 vss.n5250 vss.n5248 0.223326
R11688 vss.n5253 vss.n5251 0.223326
R11689 vss.n5256 vss.n5254 0.223326
R11690 vss.n5259 vss.n5257 0.223326
R11691 vss.n5262 vss.n5260 0.223326
R11692 vss.n5265 vss.n5263 0.223326
R11693 vss.n5268 vss.n5266 0.223326
R11694 vss.n5271 vss.n5269 0.223326
R11695 vss.n5274 vss.n5272 0.223326
R11696 vss.n5277 vss.n5275 0.223326
R11697 vss.n5280 vss.n5278 0.223326
R11698 vss.n5283 vss.n5281 0.223326
R11699 vss.n5286 vss.n5284 0.223326
R11700 vss.n5289 vss.n5287 0.223326
R11701 vss.n5292 vss.n5290 0.223326
R11702 vss.n5295 vss.n5293 0.223326
R11703 vss.n5298 vss.n5296 0.223326
R11704 vss.n5301 vss.n5299 0.223326
R11705 vss.n5303 vss.n5302 0.223326
R11706 vss.n5306 vss.n5304 0.223326
R11707 vss.n5309 vss.n5307 0.223326
R11708 vss.n5312 vss.n5310 0.223326
R11709 vss.n5315 vss.n5313 0.223326
R11710 vss.n5318 vss.n5316 0.223326
R11711 vss.n5321 vss.n5319 0.223326
R11712 vss.n5324 vss.n5322 0.223326
R11713 vss.n5326 vss.n5325 0.223326
R11714 vss.n5328 vss.n5327 0.223326
R11715 vss.n5140 vss.n5139 0.223326
R11716 vss.n5137 vss.n5136 0.223326
R11717 vss.n5134 vss.n5133 0.223326
R11718 vss.n5131 vss.n5130 0.223326
R11719 vss.n5128 vss.n5127 0.223326
R11720 vss.n5125 vss.n5124 0.223326
R11721 vss.n5122 vss.n5121 0.223326
R11722 vss.n5119 vss.n5118 0.223326
R11723 vss.n5116 vss.n5115 0.223326
R11724 vss.n5113 vss.n5112 0.223326
R11725 vss.n5110 vss.n5109 0.223326
R11726 vss.n5107 vss.n5106 0.223326
R11727 vss.n5104 vss.n5103 0.223326
R11728 vss.n5101 vss.n5100 0.223326
R11729 vss.n5098 vss.n5097 0.223326
R11730 vss.n5095 vss.n5094 0.223326
R11731 vss.n5092 vss.n5091 0.223326
R11732 vss.n5089 vss.n5088 0.223326
R11733 vss.n5086 vss.n5085 0.223326
R11734 vss.n5083 vss.n5082 0.223326
R11735 vss.n5080 vss.n5079 0.223326
R11736 vss.n5077 vss.n5076 0.223326
R11737 vss.n5074 vss.n5073 0.223326
R11738 vss.n5071 vss.n5070 0.223326
R11739 vss.n5068 vss.n5067 0.223326
R11740 vss.n5065 vss.n5064 0.223326
R11741 vss.n5062 vss.n5061 0.223326
R11742 vss.n5059 vss.n5058 0.223326
R11743 vss.n5056 vss.n5055 0.223326
R11744 vss.n5053 vss.n5052 0.223326
R11745 vss.n5050 vss.n5049 0.223326
R11746 vss.n5047 vss.n5046 0.223326
R11747 vss.n5044 vss.n5043 0.223326
R11748 vss.n5041 vss.n5040 0.223326
R11749 vss.n5038 vss.n5037 0.223326
R11750 vss.n5035 vss.n5034 0.223326
R11751 vss.n5032 vss.n5031 0.223326
R11752 vss.n5029 vss.n5028 0.223326
R11753 vss.n5026 vss.n5025 0.223326
R11754 vss.n5023 vss.n743 0.223326
R11755 vss.n971 vss.n744 0.223326
R11756 vss.n974 vss.n972 0.223326
R11757 vss.n977 vss.n975 0.223326
R11758 vss.n980 vss.n978 0.223326
R11759 vss.n983 vss.n981 0.223326
R11760 vss.n986 vss.n984 0.223326
R11761 vss.n989 vss.n987 0.223326
R11762 vss.n991 vss.n990 0.223326
R11763 vss.n993 vss.n992 0.223326
R11764 vss.n4748 vss.n4746 0.223326
R11765 vss.n4751 vss.n4749 0.223326
R11766 vss.n4754 vss.n4752 0.223326
R11767 vss.n4757 vss.n4755 0.223326
R11768 vss.n4760 vss.n4758 0.223326
R11769 vss.n4763 vss.n4761 0.223326
R11770 vss.n4766 vss.n4764 0.223326
R11771 vss.n4769 vss.n4767 0.223326
R11772 vss.n4772 vss.n4770 0.223326
R11773 vss.n4775 vss.n4773 0.223326
R11774 vss.n4778 vss.n4776 0.223326
R11775 vss.n4781 vss.n4779 0.223326
R11776 vss.n4784 vss.n4782 0.223326
R11777 vss.n4787 vss.n4785 0.223326
R11778 vss.n4790 vss.n4788 0.223326
R11779 vss.n4793 vss.n4791 0.223326
R11780 vss.n4796 vss.n4794 0.223326
R11781 vss.n4799 vss.n4797 0.223326
R11782 vss.n4802 vss.n4800 0.223326
R11783 vss.n4805 vss.n4803 0.223326
R11784 vss.n4808 vss.n4806 0.223326
R11785 vss.n4811 vss.n4809 0.223326
R11786 vss.n4814 vss.n4812 0.223326
R11787 vss.n4817 vss.n4815 0.223326
R11788 vss.n4820 vss.n4818 0.223326
R11789 vss.n4823 vss.n4821 0.223326
R11790 vss.n4826 vss.n4824 0.223326
R11791 vss.n4829 vss.n4827 0.223326
R11792 vss.n4832 vss.n4830 0.223326
R11793 vss.n4835 vss.n4833 0.223326
R11794 vss.n4838 vss.n4836 0.223326
R11795 vss.n4841 vss.n4839 0.223326
R11796 vss.n4844 vss.n4842 0.223326
R11797 vss.n4847 vss.n4845 0.223326
R11798 vss.n4850 vss.n4848 0.223326
R11799 vss.n4853 vss.n4851 0.223326
R11800 vss.n4856 vss.n4854 0.223326
R11801 vss.n4859 vss.n4857 0.223326
R11802 vss.n4862 vss.n4860 0.223326
R11803 vss.n4894 vss.n4863 0.223326
R11804 vss.n4893 vss.n4892 0.223326
R11805 vss.n4890 vss.n4889 0.223326
R11806 vss.n4887 vss.n4886 0.223326
R11807 vss.n4884 vss.n4883 0.223326
R11808 vss.n4881 vss.n4880 0.223326
R11809 vss.n4878 vss.n4877 0.223326
R11810 vss.n4875 vss.n4874 0.223326
R11811 vss.n4872 vss.n4871 0.223326
R11812 vss.n4870 vss.n4869 0.223326
R11813 vss.n5018 vss.n5017 0.223326
R11814 vss.n5015 vss.n5014 0.223326
R11815 vss.n5012 vss.n5011 0.223326
R11816 vss.n5009 vss.n5008 0.223326
R11817 vss.n5006 vss.n5005 0.223326
R11818 vss.n5003 vss.n5002 0.223326
R11819 vss.n5000 vss.n4999 0.223326
R11820 vss.n4997 vss.n4996 0.223326
R11821 vss.n4994 vss.n4993 0.223326
R11822 vss.n4991 vss.n4990 0.223326
R11823 vss.n4988 vss.n4987 0.223326
R11824 vss.n4985 vss.n4984 0.223326
R11825 vss.n4982 vss.n4981 0.223326
R11826 vss.n4979 vss.n4978 0.223326
R11827 vss.n4976 vss.n4975 0.223326
R11828 vss.n4973 vss.n4972 0.223326
R11829 vss.n4970 vss.n4969 0.223326
R11830 vss.n4967 vss.n4966 0.223326
R11831 vss.n4964 vss.n4963 0.223326
R11832 vss.n4961 vss.n4960 0.223326
R11833 vss.n4958 vss.n4957 0.223326
R11834 vss.n4955 vss.n4954 0.223326
R11835 vss.n4952 vss.n4951 0.223326
R11836 vss.n4949 vss.n4948 0.223326
R11837 vss.n4946 vss.n4945 0.223326
R11838 vss.n4943 vss.n4942 0.223326
R11839 vss.n4940 vss.n4939 0.223326
R11840 vss.n4937 vss.n4936 0.223326
R11841 vss.n4934 vss.n4933 0.223326
R11842 vss.n4931 vss.n4930 0.223326
R11843 vss.n4928 vss.n4927 0.223326
R11844 vss.n4925 vss.n4924 0.223326
R11845 vss.n4922 vss.n4921 0.223326
R11846 vss.n4919 vss.n4918 0.223326
R11847 vss.n4916 vss.n4915 0.223326
R11848 vss.n4913 vss.n4912 0.223326
R11849 vss.n4910 vss.n4909 0.223326
R11850 vss.n4907 vss.n4906 0.223326
R11851 vss.n4904 vss.n4903 0.223326
R11852 vss.n4901 vss.n4900 0.223326
R11853 vss.n4265 vss.n4264 0.223326
R11854 vss.n4262 vss.n4261 0.223326
R11855 vss.n4259 vss.n4258 0.223326
R11856 vss.n4256 vss.n4255 0.223326
R11857 vss.n4253 vss.n4252 0.223326
R11858 vss.n4250 vss.n4249 0.223326
R11859 vss.n4247 vss.n4246 0.223326
R11860 vss.n4244 vss.n4243 0.223326
R11861 vss.n4242 vss.n4241 0.223326
R11862 vss.n4594 vss.n4592 0.223326
R11863 vss.n4597 vss.n4595 0.223326
R11864 vss.n4600 vss.n4598 0.223326
R11865 vss.n4603 vss.n4601 0.223326
R11866 vss.n4606 vss.n4604 0.223326
R11867 vss.n4609 vss.n4607 0.223326
R11868 vss.n4612 vss.n4610 0.223326
R11869 vss.n4615 vss.n4613 0.223326
R11870 vss.n4618 vss.n4616 0.223326
R11871 vss.n4621 vss.n4619 0.223326
R11872 vss.n4624 vss.n4622 0.223326
R11873 vss.n4627 vss.n4625 0.223326
R11874 vss.n4630 vss.n4628 0.223326
R11875 vss.n4633 vss.n4631 0.223326
R11876 vss.n4636 vss.n4634 0.223326
R11877 vss.n4639 vss.n4637 0.223326
R11878 vss.n4642 vss.n4640 0.223326
R11879 vss.n4645 vss.n4643 0.223326
R11880 vss.n4648 vss.n4646 0.223326
R11881 vss.n4651 vss.n4649 0.223326
R11882 vss.n4654 vss.n4652 0.223326
R11883 vss.n4657 vss.n4655 0.223326
R11884 vss.n4660 vss.n4658 0.223326
R11885 vss.n4663 vss.n4661 0.223326
R11886 vss.n4666 vss.n4664 0.223326
R11887 vss.n4669 vss.n4667 0.223326
R11888 vss.n4672 vss.n4670 0.223326
R11889 vss.n4675 vss.n4673 0.223326
R11890 vss.n4678 vss.n4676 0.223326
R11891 vss.n4681 vss.n4679 0.223326
R11892 vss.n4684 vss.n4682 0.223326
R11893 vss.n4687 vss.n4685 0.223326
R11894 vss.n4690 vss.n4688 0.223326
R11895 vss.n4693 vss.n4691 0.223326
R11896 vss.n4696 vss.n4694 0.223326
R11897 vss.n4699 vss.n4697 0.223326
R11898 vss.n4702 vss.n4700 0.223326
R11899 vss.n4705 vss.n4703 0.223326
R11900 vss.n4708 vss.n4706 0.223326
R11901 vss.n4740 vss.n4709 0.223326
R11902 vss.n4739 vss.n4738 0.223326
R11903 vss.n4736 vss.n4735 0.223326
R11904 vss.n4733 vss.n4732 0.223326
R11905 vss.n4730 vss.n4729 0.223326
R11906 vss.n4727 vss.n4726 0.223326
R11907 vss.n4724 vss.n4723 0.223326
R11908 vss.n4721 vss.n4720 0.223326
R11909 vss.n4718 vss.n4717 0.223326
R11910 vss.n4716 vss.n4715 0.223326
R11911 vss.n4334 vss.n4332 0.223326
R11912 vss.n4337 vss.n4335 0.223326
R11913 vss.n4340 vss.n4338 0.223326
R11914 vss.n4343 vss.n4341 0.223326
R11915 vss.n4346 vss.n4344 0.223326
R11916 vss.n4349 vss.n4347 0.223326
R11917 vss.n2220 vss.n2208 0.207022
R11918 vss.n4220 vss.n4219 0.207022
R11919 vss.n2977 vss.n2976 0.207022
R11920 vss.n2407 vss.n2406 0.207022
R11921 vss.n2441 vss.n2440 0.207022
R11922 vss.n5778 vss.n5777 0.206263
R11923 vss.n4366 vss.n4365 0.20611
R11924 vss.n5800 vss.n5799 0.20461
R11925 vss.n5799 vss.n5798 0.201088
R11926 vss.n5765 vss.n5762 0.201088
R11927 vss.n5793 vss.n5792 0.201088
R11928 vss.n5791 vss.n5764 0.201088
R11929 vss.n5790 vss.n5789 0.201088
R11930 vss.n5788 vss.n5766 0.201088
R11931 vss.n5787 vss.n5786 0.201088
R11932 vss.n5785 vss.n5770 0.201088
R11933 vss.n5784 vss.n5783 0.201088
R11934 vss.n5782 vss.n5771 0.201088
R11935 vss.n5781 vss.n5780 0.201088
R11936 vss.n5779 vss.n5776 0.201088
R11937 vss.n5797 vss.n5761 0.201088
R11938 vss.n2221 vss.n2220 0.19887
R11939 vss.n4221 vss.n4220 0.19887
R11940 vss.n2976 vss.n2969 0.19887
R11941 vss.n2406 vss.n2397 0.19887
R11942 vss.n2440 vss.n2439 0.19887
R11943 vss.n5533 vss.n5532 0.19887
R11944 vss.n301 vss.n297 0.196396
R11945 vss.n5150 vss.n5149 0.196152
R11946 vss.n5160 vss.n1091 0.196152
R11947 vss.n5162 vss.n5161 0.196152
R11948 vss.n5172 vss.n1067 0.196152
R11949 vss.n5174 vss.n5173 0.196152
R11950 vss.n5184 vss.n1043 0.196152
R11951 vss.n5186 vss.n5185 0.196152
R11952 vss.n5203 vss.n1019 0.196152
R11953 vss.n5206 vss.n5204 0.196152
R11954 vss.n5205 vss.n319 0.196152
R11955 vss.n321 vss.n320 0.196152
R11956 vss.n347 vss.n346 0.196152
R11957 vss.n349 vss.n348 0.196152
R11958 vss.n375 vss.n374 0.196152
R11959 vss.n377 vss.n376 0.196152
R11960 vss.n403 vss.n402 0.196152
R11961 vss.n405 vss.n404 0.196152
R11962 vss.n431 vss.n430 0.196152
R11963 vss.n433 vss.n432 0.196152
R11964 vss.n459 vss.n458 0.196152
R11965 vss.n461 vss.n460 0.196152
R11966 vss.n487 vss.n486 0.196152
R11967 vss.n489 vss.n488 0.196152
R11968 vss.n515 vss.n514 0.196152
R11969 vss.n517 vss.n516 0.196152
R11970 vss.n543 vss.n542 0.196152
R11971 vss.n545 vss.n544 0.196152
R11972 vss.n571 vss.n570 0.196152
R11973 vss.n573 vss.n572 0.196152
R11974 vss.n599 vss.n598 0.196152
R11975 vss.n601 vss.n600 0.196152
R11976 vss.n627 vss.n626 0.196152
R11977 vss.n629 vss.n628 0.196152
R11978 vss.n655 vss.n654 0.196152
R11979 vss.n657 vss.n656 0.196152
R11980 vss.n683 vss.n682 0.196152
R11981 vss.n685 vss.n684 0.196152
R11982 vss.n711 vss.n710 0.196152
R11983 vss.n713 vss.n712 0.196152
R11984 vss.n738 vss.n737 0.196152
R11985 vss.n913 vss.n739 0.196152
R11986 vss.n916 vss.n915 0.196152
R11987 vss.n919 vss.n918 0.196152
R11988 vss.n922 vss.n921 0.196152
R11989 vss.n925 vss.n924 0.196152
R11990 vss.n928 vss.n927 0.196152
R11991 vss.n931 vss.n930 0.196152
R11992 vss.n934 vss.n933 0.196152
R11993 vss.n936 vss.n935 0.196152
R11994 vss.n938 vss.n937 0.196152
R11995 vss.n1258 vss.n1257 0.196152
R11996 vss.n1256 vss.n1254 0.196152
R11997 vss.n1253 vss.n1251 0.196152
R11998 vss.n1250 vss.n1248 0.196152
R11999 vss.n1247 vss.n1245 0.196152
R12000 vss.n1244 vss.n1242 0.196152
R12001 vss.n1241 vss.n1239 0.196152
R12002 vss.n1238 vss.n1236 0.196152
R12003 vss.n1235 vss.n1233 0.196152
R12004 vss.n1232 vss.n1230 0.196152
R12005 vss.n1229 vss.n1227 0.196152
R12006 vss.n1226 vss.n1224 0.196152
R12007 vss.n1223 vss.n1221 0.196152
R12008 vss.n1220 vss.n1218 0.196152
R12009 vss.n1217 vss.n1215 0.196152
R12010 vss.n1214 vss.n1212 0.196152
R12011 vss.n1211 vss.n1209 0.196152
R12012 vss.n1208 vss.n1206 0.196152
R12013 vss.n1205 vss.n1203 0.196152
R12014 vss.n1202 vss.n1200 0.196152
R12015 vss.n1199 vss.n1197 0.196152
R12016 vss.n1196 vss.n1194 0.196152
R12017 vss.n1193 vss.n1191 0.196152
R12018 vss.n1190 vss.n1188 0.196152
R12019 vss.n1187 vss.n1185 0.196152
R12020 vss.n1184 vss.n1182 0.196152
R12021 vss.n1181 vss.n1179 0.196152
R12022 vss.n1178 vss.n1176 0.196152
R12023 vss.n1175 vss.n1173 0.196152
R12024 vss.n1172 vss.n1170 0.196152
R12025 vss.n1169 vss.n1167 0.196152
R12026 vss.n1166 vss.n1164 0.196152
R12027 vss.n1163 vss.n1161 0.196152
R12028 vss.n1160 vss.n1158 0.196152
R12029 vss.n1157 vss.n1155 0.196152
R12030 vss.n1154 vss.n1152 0.196152
R12031 vss.n1151 vss.n1149 0.196152
R12032 vss.n1148 vss.n1146 0.196152
R12033 vss.n1145 vss.n1143 0.196152
R12034 vss.n1142 vss.n1140 0.196152
R12035 vss.n1139 vss.n1138 0.196152
R12036 vss.n1137 vss.n1135 0.196152
R12037 vss.n1134 vss.n1132 0.196152
R12038 vss.n1131 vss.n1129 0.196152
R12039 vss.n1128 vss.n1126 0.196152
R12040 vss.n1125 vss.n1123 0.196152
R12041 vss.n1122 vss.n1120 0.196152
R12042 vss.n1119 vss.n1117 0.196152
R12043 vss.n904 vss.n903 0.196152
R12044 vss.n906 vss.n905 0.196152
R12045 vss.n5154 vss.n1103 0.196152
R12046 vss.n5156 vss.n5155 0.196152
R12047 vss.n5166 vss.n1079 0.196152
R12048 vss.n5168 vss.n5167 0.196152
R12049 vss.n5178 vss.n1055 0.196152
R12050 vss.n5180 vss.n5179 0.196152
R12051 vss.n5190 vss.n1031 0.196152
R12052 vss.n5192 vss.n5191 0.196152
R12053 vss.n5198 vss.n5197 0.196152
R12054 vss.n5196 vss.n5194 0.196152
R12055 vss.n5193 vss.n333 0.196152
R12056 vss.n335 vss.n334 0.196152
R12057 vss.n361 vss.n360 0.196152
R12058 vss.n363 vss.n362 0.196152
R12059 vss.n389 vss.n388 0.196152
R12060 vss.n391 vss.n390 0.196152
R12061 vss.n417 vss.n416 0.196152
R12062 vss.n419 vss.n418 0.196152
R12063 vss.n445 vss.n444 0.196152
R12064 vss.n447 vss.n446 0.196152
R12065 vss.n473 vss.n472 0.196152
R12066 vss.n475 vss.n474 0.196152
R12067 vss.n501 vss.n500 0.196152
R12068 vss.n503 vss.n502 0.196152
R12069 vss.n529 vss.n528 0.196152
R12070 vss.n531 vss.n530 0.196152
R12071 vss.n557 vss.n556 0.196152
R12072 vss.n559 vss.n558 0.196152
R12073 vss.n585 vss.n584 0.196152
R12074 vss.n587 vss.n586 0.196152
R12075 vss.n613 vss.n612 0.196152
R12076 vss.n615 vss.n614 0.196152
R12077 vss.n641 vss.n640 0.196152
R12078 vss.n643 vss.n642 0.196152
R12079 vss.n669 vss.n668 0.196152
R12080 vss.n671 vss.n670 0.196152
R12081 vss.n697 vss.n696 0.196152
R12082 vss.n699 vss.n698 0.196152
R12083 vss.n725 vss.n724 0.196152
R12084 vss.n727 vss.n726 0.196152
R12085 vss.n758 vss.n757 0.196152
R12086 vss.n760 vss.n759 0.196152
R12087 vss.n945 vss.n944 0.196152
R12088 vss.n948 vss.n947 0.196152
R12089 vss.n951 vss.n950 0.196152
R12090 vss.n954 vss.n953 0.196152
R12091 vss.n957 vss.n956 0.196152
R12092 vss.n960 vss.n959 0.196152
R12093 vss.n962 vss.n961 0.196152
R12094 vss.n964 vss.n963 0.196152
R12095 vss.n1285 vss.n1284 0.196152
R12096 vss.n1283 vss.n1281 0.196152
R12097 vss.n1280 vss.n1278 0.196152
R12098 vss.n1277 vss.n1275 0.196152
R12099 vss.n1274 vss.n1272 0.196152
R12100 vss.n1271 vss.n1269 0.196152
R12101 vss.n1268 vss.n1266 0.196152
R12102 vss.n1265 vss.n1263 0.196152
R12103 vss.n1262 vss.n1007 0.196152
R12104 vss.n5212 vss.n5211 0.196152
R12105 vss.n5215 vss.n5214 0.196152
R12106 vss.n5218 vss.n5217 0.196152
R12107 vss.n5221 vss.n5220 0.196152
R12108 vss.n5224 vss.n5223 0.196152
R12109 vss.n5227 vss.n5226 0.196152
R12110 vss.n5230 vss.n5229 0.196152
R12111 vss.n5233 vss.n5232 0.196152
R12112 vss.n5236 vss.n5235 0.196152
R12113 vss.n5239 vss.n5238 0.196152
R12114 vss.n5242 vss.n5241 0.196152
R12115 vss.n5245 vss.n5244 0.196152
R12116 vss.n5248 vss.n5247 0.196152
R12117 vss.n5251 vss.n5250 0.196152
R12118 vss.n5254 vss.n5253 0.196152
R12119 vss.n5257 vss.n5256 0.196152
R12120 vss.n5260 vss.n5259 0.196152
R12121 vss.n5263 vss.n5262 0.196152
R12122 vss.n5266 vss.n5265 0.196152
R12123 vss.n5269 vss.n5268 0.196152
R12124 vss.n5272 vss.n5271 0.196152
R12125 vss.n5275 vss.n5274 0.196152
R12126 vss.n5278 vss.n5277 0.196152
R12127 vss.n5281 vss.n5280 0.196152
R12128 vss.n5284 vss.n5283 0.196152
R12129 vss.n5287 vss.n5286 0.196152
R12130 vss.n5290 vss.n5289 0.196152
R12131 vss.n5293 vss.n5292 0.196152
R12132 vss.n5296 vss.n5295 0.196152
R12133 vss.n5299 vss.n5298 0.196152
R12134 vss.n5302 vss.n5301 0.196152
R12135 vss.n5304 vss.n5303 0.196152
R12136 vss.n5307 vss.n5306 0.196152
R12137 vss.n5310 vss.n5309 0.196152
R12138 vss.n5313 vss.n5312 0.196152
R12139 vss.n5316 vss.n5315 0.196152
R12140 vss.n5319 vss.n5318 0.196152
R12141 vss.n5322 vss.n5321 0.196152
R12142 vss.n5325 vss.n5324 0.196152
R12143 vss.n5327 vss.n5326 0.196152
R12144 vss.n5329 vss.n5328 0.196152
R12145 vss.n5141 vss.n5140 0.196152
R12146 vss.n5139 vss.n5137 0.196152
R12147 vss.n5136 vss.n5134 0.196152
R12148 vss.n5133 vss.n5131 0.196152
R12149 vss.n5130 vss.n5128 0.196152
R12150 vss.n5127 vss.n5125 0.196152
R12151 vss.n5124 vss.n5122 0.196152
R12152 vss.n5121 vss.n5119 0.196152
R12153 vss.n5118 vss.n5116 0.196152
R12154 vss.n5115 vss.n5113 0.196152
R12155 vss.n5112 vss.n5110 0.196152
R12156 vss.n5109 vss.n5107 0.196152
R12157 vss.n5106 vss.n5104 0.196152
R12158 vss.n5103 vss.n5101 0.196152
R12159 vss.n5100 vss.n5098 0.196152
R12160 vss.n5097 vss.n5095 0.196152
R12161 vss.n5094 vss.n5092 0.196152
R12162 vss.n5091 vss.n5089 0.196152
R12163 vss.n5088 vss.n5086 0.196152
R12164 vss.n5085 vss.n5083 0.196152
R12165 vss.n5082 vss.n5080 0.196152
R12166 vss.n5079 vss.n5077 0.196152
R12167 vss.n5076 vss.n5074 0.196152
R12168 vss.n5073 vss.n5071 0.196152
R12169 vss.n5070 vss.n5068 0.196152
R12170 vss.n5067 vss.n5065 0.196152
R12171 vss.n5064 vss.n5062 0.196152
R12172 vss.n5061 vss.n5059 0.196152
R12173 vss.n5058 vss.n5056 0.196152
R12174 vss.n5055 vss.n5053 0.196152
R12175 vss.n5052 vss.n5050 0.196152
R12176 vss.n5049 vss.n5047 0.196152
R12177 vss.n5046 vss.n5044 0.196152
R12178 vss.n5043 vss.n5041 0.196152
R12179 vss.n5040 vss.n5038 0.196152
R12180 vss.n5037 vss.n5035 0.196152
R12181 vss.n5034 vss.n5032 0.196152
R12182 vss.n5031 vss.n5029 0.196152
R12183 vss.n5028 vss.n5026 0.196152
R12184 vss.n5025 vss.n5023 0.196152
R12185 vss.n744 vss.n743 0.196152
R12186 vss.n972 vss.n971 0.196152
R12187 vss.n975 vss.n974 0.196152
R12188 vss.n978 vss.n977 0.196152
R12189 vss.n981 vss.n980 0.196152
R12190 vss.n984 vss.n983 0.196152
R12191 vss.n987 vss.n986 0.196152
R12192 vss.n990 vss.n989 0.196152
R12193 vss.n992 vss.n991 0.196152
R12194 vss.n994 vss.n993 0.196152
R12195 vss.n4746 vss.n4745 0.196152
R12196 vss.n4749 vss.n4748 0.196152
R12197 vss.n4752 vss.n4751 0.196152
R12198 vss.n4755 vss.n4754 0.196152
R12199 vss.n4758 vss.n4757 0.196152
R12200 vss.n4761 vss.n4760 0.196152
R12201 vss.n4764 vss.n4763 0.196152
R12202 vss.n4767 vss.n4766 0.196152
R12203 vss.n4770 vss.n4769 0.196152
R12204 vss.n4773 vss.n4772 0.196152
R12205 vss.n4776 vss.n4775 0.196152
R12206 vss.n4779 vss.n4778 0.196152
R12207 vss.n4782 vss.n4781 0.196152
R12208 vss.n4785 vss.n4784 0.196152
R12209 vss.n4788 vss.n4787 0.196152
R12210 vss.n4791 vss.n4790 0.196152
R12211 vss.n4794 vss.n4793 0.196152
R12212 vss.n4797 vss.n4796 0.196152
R12213 vss.n4800 vss.n4799 0.196152
R12214 vss.n4803 vss.n4802 0.196152
R12215 vss.n4806 vss.n4805 0.196152
R12216 vss.n4809 vss.n4808 0.196152
R12217 vss.n4812 vss.n4811 0.196152
R12218 vss.n4815 vss.n4814 0.196152
R12219 vss.n4818 vss.n4817 0.196152
R12220 vss.n4821 vss.n4820 0.196152
R12221 vss.n4824 vss.n4823 0.196152
R12222 vss.n4827 vss.n4826 0.196152
R12223 vss.n4830 vss.n4829 0.196152
R12224 vss.n4833 vss.n4832 0.196152
R12225 vss.n4836 vss.n4835 0.196152
R12226 vss.n4839 vss.n4838 0.196152
R12227 vss.n4842 vss.n4841 0.196152
R12228 vss.n4845 vss.n4844 0.196152
R12229 vss.n4848 vss.n4847 0.196152
R12230 vss.n4851 vss.n4850 0.196152
R12231 vss.n4854 vss.n4853 0.196152
R12232 vss.n4857 vss.n4856 0.196152
R12233 vss.n4860 vss.n4859 0.196152
R12234 vss.n4863 vss.n4862 0.196152
R12235 vss.n4894 vss.n4893 0.196152
R12236 vss.n4892 vss.n4890 0.196152
R12237 vss.n4889 vss.n4887 0.196152
R12238 vss.n4886 vss.n4884 0.196152
R12239 vss.n4883 vss.n4881 0.196152
R12240 vss.n4880 vss.n4878 0.196152
R12241 vss.n4877 vss.n4875 0.196152
R12242 vss.n4874 vss.n4872 0.196152
R12243 vss.n4871 vss.n4870 0.196152
R12244 vss.n4869 vss.n4864 0.196152
R12245 vss.n5019 vss.n5018 0.196152
R12246 vss.n5017 vss.n5015 0.196152
R12247 vss.n5014 vss.n5012 0.196152
R12248 vss.n5011 vss.n5009 0.196152
R12249 vss.n5008 vss.n5006 0.196152
R12250 vss.n5005 vss.n5003 0.196152
R12251 vss.n5002 vss.n5000 0.196152
R12252 vss.n4999 vss.n4997 0.196152
R12253 vss.n4996 vss.n4994 0.196152
R12254 vss.n4993 vss.n4991 0.196152
R12255 vss.n4990 vss.n4988 0.196152
R12256 vss.n4987 vss.n4985 0.196152
R12257 vss.n4984 vss.n4982 0.196152
R12258 vss.n4981 vss.n4979 0.196152
R12259 vss.n4978 vss.n4976 0.196152
R12260 vss.n4975 vss.n4973 0.196152
R12261 vss.n4972 vss.n4970 0.196152
R12262 vss.n4969 vss.n4967 0.196152
R12263 vss.n4966 vss.n4964 0.196152
R12264 vss.n4963 vss.n4961 0.196152
R12265 vss.n4960 vss.n4958 0.196152
R12266 vss.n4957 vss.n4955 0.196152
R12267 vss.n4954 vss.n4952 0.196152
R12268 vss.n4951 vss.n4949 0.196152
R12269 vss.n4948 vss.n4946 0.196152
R12270 vss.n4945 vss.n4943 0.196152
R12271 vss.n4942 vss.n4940 0.196152
R12272 vss.n4939 vss.n4937 0.196152
R12273 vss.n4936 vss.n4934 0.196152
R12274 vss.n4933 vss.n4931 0.196152
R12275 vss.n4930 vss.n4928 0.196152
R12276 vss.n4927 vss.n4925 0.196152
R12277 vss.n4924 vss.n4922 0.196152
R12278 vss.n4921 vss.n4919 0.196152
R12279 vss.n4918 vss.n4916 0.196152
R12280 vss.n4915 vss.n4913 0.196152
R12281 vss.n4912 vss.n4910 0.196152
R12282 vss.n4909 vss.n4907 0.196152
R12283 vss.n4906 vss.n4904 0.196152
R12284 vss.n4903 vss.n4901 0.196152
R12285 vss.n4900 vss.n4265 0.196152
R12286 vss.n4264 vss.n4262 0.196152
R12287 vss.n4261 vss.n4259 0.196152
R12288 vss.n4258 vss.n4256 0.196152
R12289 vss.n4255 vss.n4253 0.196152
R12290 vss.n4252 vss.n4250 0.196152
R12291 vss.n4249 vss.n4247 0.196152
R12292 vss.n4246 vss.n4244 0.196152
R12293 vss.n4243 vss.n4242 0.196152
R12294 vss.n4241 vss.n4236 0.196152
R12295 vss.n4592 vss.n4591 0.196152
R12296 vss.n4595 vss.n4594 0.196152
R12297 vss.n4598 vss.n4597 0.196152
R12298 vss.n4601 vss.n4600 0.196152
R12299 vss.n4604 vss.n4603 0.196152
R12300 vss.n4607 vss.n4606 0.196152
R12301 vss.n4610 vss.n4609 0.196152
R12302 vss.n4613 vss.n4612 0.196152
R12303 vss.n4616 vss.n4615 0.196152
R12304 vss.n4619 vss.n4618 0.196152
R12305 vss.n4622 vss.n4621 0.196152
R12306 vss.n4625 vss.n4624 0.196152
R12307 vss.n4628 vss.n4627 0.196152
R12308 vss.n4631 vss.n4630 0.196152
R12309 vss.n4634 vss.n4633 0.196152
R12310 vss.n4637 vss.n4636 0.196152
R12311 vss.n4640 vss.n4639 0.196152
R12312 vss.n4643 vss.n4642 0.196152
R12313 vss.n4646 vss.n4645 0.196152
R12314 vss.n4649 vss.n4648 0.196152
R12315 vss.n4652 vss.n4651 0.196152
R12316 vss.n4655 vss.n4654 0.196152
R12317 vss.n4658 vss.n4657 0.196152
R12318 vss.n4661 vss.n4660 0.196152
R12319 vss.n4664 vss.n4663 0.196152
R12320 vss.n4667 vss.n4666 0.196152
R12321 vss.n4670 vss.n4669 0.196152
R12322 vss.n4673 vss.n4672 0.196152
R12323 vss.n4676 vss.n4675 0.196152
R12324 vss.n4679 vss.n4678 0.196152
R12325 vss.n4682 vss.n4681 0.196152
R12326 vss.n4685 vss.n4684 0.196152
R12327 vss.n4688 vss.n4687 0.196152
R12328 vss.n4691 vss.n4690 0.196152
R12329 vss.n4694 vss.n4693 0.196152
R12330 vss.n4697 vss.n4696 0.196152
R12331 vss.n4700 vss.n4699 0.196152
R12332 vss.n4703 vss.n4702 0.196152
R12333 vss.n4706 vss.n4705 0.196152
R12334 vss.n4709 vss.n4708 0.196152
R12335 vss.n4740 vss.n4739 0.196152
R12336 vss.n4738 vss.n4736 0.196152
R12337 vss.n4735 vss.n4733 0.196152
R12338 vss.n4732 vss.n4730 0.196152
R12339 vss.n4729 vss.n4727 0.196152
R12340 vss.n4726 vss.n4724 0.196152
R12341 vss.n4723 vss.n4721 0.196152
R12342 vss.n4720 vss.n4718 0.196152
R12343 vss.n4717 vss.n4716 0.196152
R12344 vss.n4715 vss.n4710 0.196152
R12345 vss.n4332 vss.n4331 0.196152
R12346 vss.n4335 vss.n4334 0.196152
R12347 vss.n4338 vss.n4337 0.196152
R12348 vss.n4341 vss.n4340 0.196152
R12349 vss.n4344 vss.n4343 0.196152
R12350 vss.n4347 vss.n4346 0.196152
R12351 vss.n4350 vss.n4349 0.192188
R12352 vss.n5796 vss.n5760 0.141503
R12353 vss.n5777 vss.n5775 0.141503
R12354 vss.n5542 vss.n5541 0.13856
R12355 vss.n4371 vss.n4365 0.13856
R12356 vss.n4372 vss.n4371 0.13856
R12357 vss.n4381 vss.n4378 0.0900522
R12358 vss.n4377 vss.n4360 0.0881866
R12359 vss.n4585 vss.n4584 0.0755
R12360 vss.n298 vss.n295 0.0688282
R12361 vss.n4585 vss.n4575 0.0674118
R12362 vss.n4369 vss.n4364 0.0647361
R12363 vss.n5565 vss.n5564 0.063
R12364 vss.n5564 vss.n5563 0.063
R12365 vss.n5563 vss.n5562 0.063
R12366 vss.n5560 vss.n5559 0.063
R12367 vss.n5557 vss.n5556 0.063
R12368 vss.n5556 vss.n5555 0.063
R12369 vss.n5553 vss.n5552 0.063
R12370 vss.n5552 vss.n5551 0.063
R12371 vss.n5621 vss.n5620 0.063
R12372 vss.n5622 vss.n5621 0.063
R12373 vss.n5901 vss.n5624 0.063
R12374 vss.n5901 vss.n5900 0.063
R12375 vss.n5639 vss.n5638 0.063
R12376 vss.n5890 vss.n5639 0.063
R12377 vss.n5888 vss.n5641 0.063
R12378 vss.n5658 vss.n5641 0.063
R12379 vss.n5874 vss.n5660 0.063
R12380 vss.n5874 vss.n5873 0.063
R12381 vss.n5873 vss.n5661 0.063
R12382 vss.n5675 vss.n5661 0.063
R12383 vss.n5863 vss.n5675 0.063
R12384 vss.n5863 vss.n5862 0.063
R12385 vss.n5696 vss.n5695 0.063
R12386 vss.n5697 vss.n5696 0.063
R12387 vss.n5848 vss.n5847 0.063
R12388 vss.n5847 vss.n5699 0.063
R12389 vss.n5837 vss.n5713 0.063
R12390 vss.n5837 vss.n5836 0.063
R12391 vss.n5735 vss.n5734 0.063
R12392 vss.n5736 vss.n5735 0.063
R12393 vss.n5822 vss.n5821 0.063
R12394 vss.n5821 vss.n5738 0.063
R12395 vss.n5811 vss.n5752 0.063
R12396 vss.n5811 vss.n5810 0.063
R12397 vss.n5801 vss.n5759 0.063
R12398 vss.n4352 vss.n4326 0.063
R12399 vss.n4414 vss.n4310 0.063
R12400 vss.n4421 vss.n4310 0.063
R12401 vss.n4422 vss.n4421 0.063
R12402 vss.n4429 vss.n4426 0.063
R12403 vss.n4436 vss.n4303 0.063
R12404 vss.n4439 vss.n4436 0.063
R12405 vss.n4446 vss.n4301 0.063
R12406 vss.n4449 vss.n4446 0.063
R12407 vss.n4456 vss.n4298 0.063
R12408 vss.n4459 vss.n4456 0.063
R12409 vss.n4466 vss.n4296 0.063
R12410 vss.n4469 vss.n4466 0.063
R12411 vss.n4476 vss.n4293 0.063
R12412 vss.n4479 vss.n4476 0.063
R12413 vss.n4489 vss.n4291 0.063
R12414 vss.n4490 vss.n4489 0.063
R12415 vss.n4492 vss.n4289 0.063
R12416 vss.n4500 vss.n4289 0.063
R12417 vss.n4501 vss.n4500 0.063
R12418 vss.n4501 vss.n4287 0.063
R12419 vss.n4508 vss.n4287 0.063
R12420 vss.n4511 vss.n4508 0.063
R12421 vss.n4518 vss.n4283 0.063
R12422 vss.n4521 vss.n4518 0.063
R12423 vss.n4528 vss.n4281 0.063
R12424 vss.n4531 vss.n4528 0.063
R12425 vss.n4538 vss.n4278 0.063
R12426 vss.n4541 vss.n4538 0.063
R12427 vss.n4548 vss.n4276 0.063
R12428 vss.n4551 vss.n4548 0.063
R12429 vss.n4558 vss.n4273 0.063
R12430 vss.n4561 vss.n4558 0.063
R12431 vss.n4568 vss.n4271 0.063
R12432 vss.n4569 vss.n4568 0.063
R12433 vss.n5561 vss.n5560 0.0614375
R12434 vss.n5559 vss.n5558 0.0614375
R12435 vss.n4426 vss.n4307 0.0614375
R12436 vss.n4429 vss.n4428 0.0614375
R12437 vss.n5862 vss.n5677 0.059875
R12438 vss.n4511 vss.n4510 0.059875
R12439 vss.n4494 vss.n4290 0.0593235
R12440 vss.n4573 vss.n4570 0.0593235
R12441 vss.n4382 vss.n4381 0.0583358
R12442 vss.n5555 vss.n5554 0.0583125
R12443 vss.n4439 vss.n4438 0.0583125
R12444 vss.n4405 vss.n4402 0.0578529
R12445 vss.n4411 vss.n4409 0.0578529
R12446 vss.n5698 vss.n5697 0.05675
R12447 vss.n4521 vss.n4520 0.05675
R12448 vss.n4488 vss.n4484 0.0563824
R12449 vss.n5551 vss.n242 0.0551875
R12450 vss.n4449 vss.n4448 0.0551875
R12451 vss.n4498 vss.n4496 0.0549118
R12452 vss.n4567 vss.n4566 0.0549118
R12453 vss.n5712 vss.n5699 0.053625
R12454 vss.n4531 vss.n4530 0.053625
R12455 vss.n4397 vss.n4396 0.0534412
R12456 vss.n4404 vss.n4314 0.0534412
R12457 vss.n4417 vss.n4415 0.0534412
R12458 vss.n4487 vss.n4485 0.0534412
R12459 vss.n4495 vss.n4494 0.0534412
R12460 vss.n4570 vss.n4270 0.0534412
R12461 vss.n4572 vss.n4267 0.0534412
R12462 vss.n4580 vss.n4579 0.0533351
R12463 vss.n790 vss.n789 0.0533351
R12464 vss.n823 vss.n791 0.0533351
R12465 vss.n825 vss.n824 0.0533351
R12466 vss.n855 vss.n826 0.0533351
R12467 vss.n857 vss.n856 0.0533351
R12468 vss.n5335 vss.n858 0.0533351
R12469 vss.n5337 vss.n5336 0.0533351
R12470 vss.n5339 vss.n5338 0.0533351
R12471 vss.n2296 vss.n2235 0.0529194
R12472 vss.n5623 vss.n5622 0.0520625
R12473 vss.n4459 vss.n4458 0.0520625
R12474 vss.n4401 vss.n4317 0.0519706
R12475 vss.n4412 vss.n4311 0.0519706
R12476 vss.n4480 vss.n4292 0.0519706
R12477 vss.n4372 vss.n4360 0.0508731
R12478 vss.n5836 vss.n5715 0.0505
R12479 vss.n4541 vss.n4540 0.0505
R12480 vss.n4483 vss.n4482 0.0505
R12481 vss.n4504 vss.n4502 0.0505
R12482 vss.n4562 vss.n4272 0.0505
R12483 vss.n5545 vss.n5544 0.0492504
R12484 vss.n4391 vss.n4390 0.0490294
R12485 vss.n4420 vss.n4309 0.0490294
R12486 vss.n4499 vss.n4288 0.0490294
R12487 vss.n4565 vss.n4564 0.0490294
R12488 vss.n4378 vss.n4377 0.0490075
R12489 vss.n5900 vss.n5626 0.0489375
R12490 vss.n4469 vss.n4468 0.0489375
R12491 vss.n4395 vss.n4320 0.0475588
R12492 vss.n4419 vss.n4418 0.0475588
R12493 vss.n4472 vss.n4471 0.0475588
R12494 vss.n5737 vss.n5736 0.047375
R12495 vss.n4551 vss.n4550 0.047375
R12496 vss.n4583 vss.n4580 0.0468918
R12497 vss.n4579 vss.n789 0.0468918
R12498 vss.n791 vss.n790 0.0468918
R12499 vss.n824 vss.n823 0.0468918
R12500 vss.n826 vss.n825 0.0468918
R12501 vss.n856 vss.n855 0.0468918
R12502 vss.n858 vss.n857 0.0468918
R12503 vss.n5336 vss.n5335 0.0468918
R12504 vss.n5338 vss.n5337 0.0468918
R12505 vss.n5348 vss.n5339 0.0468918
R12506 vss.n4475 vss.n4474 0.0460882
R12507 vss.n4507 vss.n4285 0.0460882
R12508 vss.n4554 vss.n4553 0.0460882
R12509 vss.n5890 vss.n5889 0.0458125
R12510 vss.n4479 vss.n4478 0.0458125
R12511 vss.n4359 vss.n4326 0.0453569
R12512 vss.n4386 vss.n4323 0.0446176
R12513 vss.n4425 vss.n4305 0.0446176
R12514 vss.n4506 vss.n4505 0.0446176
R12515 vss.n4557 vss.n4556 0.0446176
R12516 vss.n4414 vss.n4413 0.0443487
R12517 vss.n5751 vss.n5738 0.04425
R12518 vss.n4561 vss.n4560 0.04425
R12519 vss.n4389 vss.n4388 0.0431471
R12520 vss.n4424 vss.n4423 0.0431471
R12521 vss.n4465 vss.n4464 0.0431471
R12522 vss.n5659 vss.n5658 0.0426875
R12523 vss.n4491 vss.n4490 0.0426875
R12524 vss.n4361 vss.n4325 0.0421667
R12525 vss.n4470 vss.n4295 0.0416765
R12526 vss.n4516 vss.n4514 0.0416765
R12527 vss.n4547 vss.n4546 0.0416765
R12528 vss.n4362 vss.n4360 0.0412986
R12529 vss.n5567 vss.n5565 0.0411764
R12530 vss.n5810 vss.n5753 0.041125
R12531 vss.n4569 vss.n4268 0.041125
R12532 vss.n4355 vss.n4354 0.0402059
R12533 vss.n4434 vss.n4432 0.0402059
R12534 vss.n4513 vss.n4512 0.0402059
R12535 vss.n4552 vss.n4275 0.0402059
R12536 vss.n5595 vss.n260 0.0399737
R12537 vss.n5910 vss.n230 0.0399737
R12538 vss.n5883 vss.n5649 0.0399737
R12539 vss.n5857 vss.n5685 0.0399737
R12540 vss.n5831 vss.n5724 0.0399737
R12541 vss.n5542 vss.n297 0.0396791
R12542 vss.n279 vss.n277 0.039413
R12543 vss.n5598 vss.n258 0.0388772
R12544 vss.n5906 vss.n233 0.0388772
R12545 vss.n5879 vss.n5651 0.0388772
R12546 vss.n5853 vss.n5687 0.0388772
R12547 vss.n5827 vss.n5726 0.0388772
R12548 vss.n4358 vss.n4357 0.0387353
R12549 vss.n4431 vss.n4430 0.0387353
R12550 vss.n4460 vss.n4297 0.0387353
R12551 vss.n3602 vss.n3082 0.0375036
R12552 vss.n3591 vss.n3590 0.0375036
R12553 vss.n3580 vss.n3579 0.0375036
R12554 vss.n3568 vss.n3092 0.0375036
R12555 vss.n3560 vss.n3096 0.0375036
R12556 vss.n3548 vss.n3547 0.0375036
R12557 vss.n3536 vss.n3535 0.0375036
R12558 vss.n3524 vss.n3120 0.0375036
R12559 vss.n3513 vss.n3131 0.0375036
R12560 vss.n3502 vss.n3146 0.0375036
R12561 vss.n3494 vss.n3154 0.0375036
R12562 vss.n3483 vss.n3165 0.0375036
R12563 vss.n3472 vss.n3180 0.0375036
R12564 vss.n3461 vss.n3460 0.0375036
R12565 vss.n3450 vss.n3449 0.0375036
R12566 vss.n3428 vss.n3215 0.0375036
R12567 vss.n3417 vss.n3226 0.0375036
R12568 vss.n3406 vss.n3241 0.0375036
R12569 vss.n3398 vss.n3249 0.0375036
R12570 vss.n3387 vss.n3260 0.0375036
R12571 vss.n3376 vss.n3275 0.0375036
R12572 vss.n3365 vss.n3364 0.0375036
R12573 vss.n3354 vss.n3353 0.0375036
R12574 vss.n3343 vss.n3342 0.0375036
R12575 vss.n3330 vss.n3329 0.0375036
R12576 vss.n6127 vss.n3 0.0375036
R12577 vss.n6119 vss.n12 0.0375036
R12578 vss.n6108 vss.n6107 0.0375036
R12579 vss.n6097 vss.n6096 0.0375036
R12580 vss.n6085 vss.n37 0.0375036
R12581 vss.n6077 vss.n47 0.0375036
R12582 vss.n6066 vss.n6065 0.0375036
R12583 vss.n6055 vss.n6054 0.0375036
R12584 vss.n6043 vss.n72 0.0375036
R12585 vss.n6035 vss.n82 0.0375036
R12586 vss.n6024 vss.n6023 0.0375036
R12587 vss.n4463 vss.n4462 0.0372647
R12588 vss.n4524 vss.n4522 0.0372647
R12589 vss.n4542 vss.n4277 0.0372647
R12590 vss.n3598 vss.n3082 0.0370523
R12591 vss.n3598 vss.n3597 0.0370523
R12592 vss.n3597 vss.n3596 0.0370523
R12593 vss.n3596 vss.n3084 0.0370523
R12594 vss.n3592 vss.n3084 0.0370523
R12595 vss.n3592 vss.n3591 0.0370523
R12596 vss.n3590 vss.n3086 0.0370523
R12597 vss.n3586 vss.n3086 0.0370523
R12598 vss.n3586 vss.n3585 0.0370523
R12599 vss.n3585 vss.n3584 0.0370523
R12600 vss.n3584 vss.n3088 0.0370523
R12601 vss.n3580 vss.n3088 0.0370523
R12602 vss.n3579 vss.n3578 0.0370523
R12603 vss.n3578 vss.n3090 0.0370523
R12604 vss.n3574 vss.n3090 0.0370523
R12605 vss.n3574 vss.n3573 0.0370523
R12606 vss.n3573 vss.n3572 0.0370523
R12607 vss.n3572 vss.n3092 0.0370523
R12608 vss.n3568 vss.n3567 0.0370523
R12609 vss.n3567 vss.n3566 0.0370523
R12610 vss.n3566 vss.n3094 0.0370523
R12611 vss.n3562 vss.n3094 0.0370523
R12612 vss.n3562 vss.n3561 0.0370523
R12613 vss.n3561 vss.n3560 0.0370523
R12614 vss.n3556 vss.n3096 0.0370523
R12615 vss.n3556 vss.n3555 0.0370523
R12616 vss.n3555 vss.n3554 0.0370523
R12617 vss.n3554 vss.n3098 0.0370523
R12618 vss.n3549 vss.n3098 0.0370523
R12619 vss.n3549 vss.n3548 0.0370523
R12620 vss.n3547 vss.n3103 0.0370523
R12621 vss.n3542 vss.n3103 0.0370523
R12622 vss.n3542 vss.n3541 0.0370523
R12623 vss.n3541 vss.n3540 0.0370523
R12624 vss.n3540 vss.n3108 0.0370523
R12625 vss.n3536 vss.n3108 0.0370523
R12626 vss.n3535 vss.n3534 0.0370523
R12627 vss.n3534 vss.n3114 0.0370523
R12628 vss.n3530 vss.n3114 0.0370523
R12629 vss.n3530 vss.n3529 0.0370523
R12630 vss.n3529 vss.n3528 0.0370523
R12631 vss.n3528 vss.n3120 0.0370523
R12632 vss.n3524 vss.n3523 0.0370523
R12633 vss.n3523 vss.n3129 0.0370523
R12634 vss.n3519 vss.n3129 0.0370523
R12635 vss.n3519 vss.n3518 0.0370523
R12636 vss.n3518 vss.n3517 0.0370523
R12637 vss.n3517 vss.n3131 0.0370523
R12638 vss.n3513 vss.n3512 0.0370523
R12639 vss.n3512 vss.n3511 0.0370523
R12640 vss.n3511 vss.n3137 0.0370523
R12641 vss.n3507 vss.n3137 0.0370523
R12642 vss.n3507 vss.n3506 0.0370523
R12643 vss.n3506 vss.n3146 0.0370523
R12644 vss.n3502 vss.n3501 0.0370523
R12645 vss.n3501 vss.n3500 0.0370523
R12646 vss.n3500 vss.n3148 0.0370523
R12647 vss.n3496 vss.n3148 0.0370523
R12648 vss.n3496 vss.n3495 0.0370523
R12649 vss.n3495 vss.n3494 0.0370523
R12650 vss.n3490 vss.n3154 0.0370523
R12651 vss.n3490 vss.n3489 0.0370523
R12652 vss.n3489 vss.n3163 0.0370523
R12653 vss.n3485 vss.n3163 0.0370523
R12654 vss.n3485 vss.n3484 0.0370523
R12655 vss.n3484 vss.n3483 0.0370523
R12656 vss.n3479 vss.n3165 0.0370523
R12657 vss.n3479 vss.n3478 0.0370523
R12658 vss.n3478 vss.n3477 0.0370523
R12659 vss.n3477 vss.n3171 0.0370523
R12660 vss.n3473 vss.n3171 0.0370523
R12661 vss.n3473 vss.n3472 0.0370523
R12662 vss.n3468 vss.n3180 0.0370523
R12663 vss.n3468 vss.n3467 0.0370523
R12664 vss.n3467 vss.n3466 0.0370523
R12665 vss.n3466 vss.n3182 0.0370523
R12666 vss.n3462 vss.n3182 0.0370523
R12667 vss.n3462 vss.n3461 0.0370523
R12668 vss.n3460 vss.n3191 0.0370523
R12669 vss.n3456 vss.n3191 0.0370523
R12670 vss.n3456 vss.n3455 0.0370523
R12671 vss.n3455 vss.n3196 0.0370523
R12672 vss.n3451 vss.n3196 0.0370523
R12673 vss.n3451 vss.n3450 0.0370523
R12674 vss.n3449 vss.n3198 0.0370523
R12675 vss.n3445 vss.n3198 0.0370523
R12676 vss.n3445 vss.n3444 0.0370523
R12677 vss.n3444 vss.n3207 0.0370523
R12678 vss.n3440 vss.n3207 0.0370523
R12679 vss.n3440 vss.n3439 0.0370523
R12680 vss.n3439 vss.n3438 0.0370523
R12681 vss.n3438 vss.n3209 0.0370523
R12682 vss.n3434 vss.n3209 0.0370523
R12683 vss.n3434 vss.n3433 0.0370523
R12684 vss.n3433 vss.n3432 0.0370523
R12685 vss.n3432 vss.n3215 0.0370523
R12686 vss.n3428 vss.n3427 0.0370523
R12687 vss.n3427 vss.n3224 0.0370523
R12688 vss.n3423 vss.n3224 0.0370523
R12689 vss.n3423 vss.n3422 0.0370523
R12690 vss.n3422 vss.n3421 0.0370523
R12691 vss.n3421 vss.n3226 0.0370523
R12692 vss.n3417 vss.n3416 0.0370523
R12693 vss.n3416 vss.n3415 0.0370523
R12694 vss.n3415 vss.n3232 0.0370523
R12695 vss.n3411 vss.n3232 0.0370523
R12696 vss.n3411 vss.n3410 0.0370523
R12697 vss.n3410 vss.n3241 0.0370523
R12698 vss.n3406 vss.n3405 0.0370523
R12699 vss.n3405 vss.n3404 0.0370523
R12700 vss.n3404 vss.n3243 0.0370523
R12701 vss.n3400 vss.n3243 0.0370523
R12702 vss.n3400 vss.n3399 0.0370523
R12703 vss.n3399 vss.n3398 0.0370523
R12704 vss.n3394 vss.n3249 0.0370523
R12705 vss.n3394 vss.n3393 0.0370523
R12706 vss.n3393 vss.n3258 0.0370523
R12707 vss.n3389 vss.n3258 0.0370523
R12708 vss.n3389 vss.n3388 0.0370523
R12709 vss.n3388 vss.n3387 0.0370523
R12710 vss.n3383 vss.n3260 0.0370523
R12711 vss.n3383 vss.n3382 0.0370523
R12712 vss.n3382 vss.n3381 0.0370523
R12713 vss.n3381 vss.n3266 0.0370523
R12714 vss.n3377 vss.n3266 0.0370523
R12715 vss.n3377 vss.n3376 0.0370523
R12716 vss.n3372 vss.n3275 0.0370523
R12717 vss.n3372 vss.n3371 0.0370523
R12718 vss.n3371 vss.n3370 0.0370523
R12719 vss.n3370 vss.n3277 0.0370523
R12720 vss.n3366 vss.n3277 0.0370523
R12721 vss.n3366 vss.n3365 0.0370523
R12722 vss.n3364 vss.n3283 0.0370523
R12723 vss.n3360 vss.n3283 0.0370523
R12724 vss.n3360 vss.n3359 0.0370523
R12725 vss.n3359 vss.n3292 0.0370523
R12726 vss.n3355 vss.n3292 0.0370523
R12727 vss.n3355 vss.n3354 0.0370523
R12728 vss.n3353 vss.n3294 0.0370523
R12729 vss.n3349 vss.n3294 0.0370523
R12730 vss.n3349 vss.n3348 0.0370523
R12731 vss.n3348 vss.n3303 0.0370523
R12732 vss.n3344 vss.n3303 0.0370523
R12733 vss.n3344 vss.n3343 0.0370523
R12734 vss.n3342 vss.n3305 0.0370523
R12735 vss.n3338 vss.n3305 0.0370523
R12736 vss.n3338 vss.n3337 0.0370523
R12737 vss.n3337 vss.n3336 0.0370523
R12738 vss.n3336 vss.n3309 0.0370523
R12739 vss.n3330 vss.n3309 0.0370523
R12740 vss.n3329 vss.n3328 0.0370523
R12741 vss.n3328 vss.n3313 0.0370523
R12742 vss.n3321 vss.n3313 0.0370523
R12743 vss.n3321 vss.n3320 0.0370523
R12744 vss.n3320 vss.n3317 0.0370523
R12745 vss.n3317 vss.n3 0.0370523
R12746 vss.n6127 vss.n6126 0.0370523
R12747 vss.n6126 vss.n6125 0.0370523
R12748 vss.n6125 vss.n7 0.0370523
R12749 vss.n6121 vss.n7 0.0370523
R12750 vss.n6121 vss.n6120 0.0370523
R12751 vss.n6120 vss.n6119 0.0370523
R12752 vss.n6115 vss.n12 0.0370523
R12753 vss.n6115 vss.n6114 0.0370523
R12754 vss.n6114 vss.n6113 0.0370523
R12755 vss.n6113 vss.n17 0.0370523
R12756 vss.n6109 vss.n17 0.0370523
R12757 vss.n6109 vss.n6108 0.0370523
R12758 vss.n6107 vss.n22 0.0370523
R12759 vss.n6103 vss.n22 0.0370523
R12760 vss.n6103 vss.n6102 0.0370523
R12761 vss.n6102 vss.n6101 0.0370523
R12762 vss.n6101 vss.n27 0.0370523
R12763 vss.n6097 vss.n27 0.0370523
R12764 vss.n6096 vss.n6095 0.0370523
R12765 vss.n6095 vss.n32 0.0370523
R12766 vss.n6091 vss.n32 0.0370523
R12767 vss.n6091 vss.n6090 0.0370523
R12768 vss.n6090 vss.n6089 0.0370523
R12769 vss.n6089 vss.n37 0.0370523
R12770 vss.n6085 vss.n6084 0.0370523
R12771 vss.n6084 vss.n6083 0.0370523
R12772 vss.n6083 vss.n42 0.0370523
R12773 vss.n6079 vss.n42 0.0370523
R12774 vss.n6079 vss.n6078 0.0370523
R12775 vss.n6078 vss.n6077 0.0370523
R12776 vss.n6073 vss.n47 0.0370523
R12777 vss.n6073 vss.n6072 0.0370523
R12778 vss.n6072 vss.n6071 0.0370523
R12779 vss.n6071 vss.n52 0.0370523
R12780 vss.n6067 vss.n52 0.0370523
R12781 vss.n6067 vss.n6066 0.0370523
R12782 vss.n6065 vss.n57 0.0370523
R12783 vss.n6061 vss.n57 0.0370523
R12784 vss.n6061 vss.n6060 0.0370523
R12785 vss.n6060 vss.n6059 0.0370523
R12786 vss.n6059 vss.n62 0.0370523
R12787 vss.n6055 vss.n62 0.0370523
R12788 vss.n6054 vss.n6053 0.0370523
R12789 vss.n6053 vss.n67 0.0370523
R12790 vss.n6049 vss.n67 0.0370523
R12791 vss.n6049 vss.n6048 0.0370523
R12792 vss.n6048 vss.n6047 0.0370523
R12793 vss.n6047 vss.n72 0.0370523
R12794 vss.n6043 vss.n6042 0.0370523
R12795 vss.n6042 vss.n6041 0.0370523
R12796 vss.n6041 vss.n77 0.0370523
R12797 vss.n6037 vss.n77 0.0370523
R12798 vss.n6037 vss.n6036 0.0370523
R12799 vss.n6036 vss.n6035 0.0370523
R12800 vss.n6031 vss.n82 0.0370523
R12801 vss.n6031 vss.n6030 0.0370523
R12802 vss.n6030 vss.n6029 0.0370523
R12803 vss.n6029 vss.n87 0.0370523
R12804 vss.n6025 vss.n87 0.0370523
R12805 vss.n6025 vss.n6024 0.0370523
R12806 vss.n6023 vss.n92 0.0370523
R12807 vss.n6019 vss.n92 0.0370523
R12808 vss.n6019 vss.n6018 0.0370523
R12809 vss.n6016 vss.n106 0.0370523
R12810 vss.n6014 vss.n6013 0.0370523
R12811 vss.n5591 vss.n264 0.0366842
R12812 vss.n5618 vss.n228 0.0366842
R12813 vss.n5886 vss.n5644 0.0366842
R12814 vss.n5860 vss.n5680 0.0366842
R12815 vss.n5834 vss.n5718 0.0366842
R12816 vss.n5808 vss.n5756 0.0366842
R12817 vss.n4214 vss.n4213 0.0361445
R12818 vss.n2449 vss.n2377 0.0361445
R12819 vss.n4351 vss.n4350 0.0357941
R12820 vss.n4442 vss.n4440 0.0357941
R12821 vss.n4517 vss.n4282 0.0357941
R12822 vss.n4545 vss.n4544 0.0357941
R12823 vss.n5573 vss.n5571 0.0357412
R12824 vss.n4209 vss.n1318 0.0356562
R12825 vss.n4210 vss.n1315 0.035168
R12826 vss.n5601 vss.n256 0.0344912
R12827 vss.n5903 vss.n236 0.0344912
R12828 vss.n5876 vss.n5654 0.0344912
R12829 vss.n5850 vss.n5690 0.0344912
R12830 vss.n5824 vss.n5729 0.0344912
R12831 vss.n4353 vss.n4328 0.0343235
R12832 vss.n4435 vss.n4302 0.0343235
R12833 vss.n4452 vss.n4451 0.0343235
R12834 vss.n4455 vss.n4454 0.0328529
R12835 vss.n4527 vss.n4280 0.0328529
R12836 vss.n4534 vss.n4533 0.0328529
R12837 vss.n4217 vss.n1312 0.0327266
R12838 vss.n5803 vss.n5802 0.0324147
R12839 vss.n5587 vss.n262 0.0322982
R12840 vss.n5619 vss.n243 0.0322982
R12841 vss.n5887 vss.n5637 0.0322982
R12842 vss.n5861 vss.n5673 0.0322982
R12843 vss.n5835 vss.n5710 0.0322982
R12844 vss.n5809 vss.n5749 0.0322982
R12845 vss.n2986 vss.n2985 0.03175
R12846 vss.n3613 vss.n3071 0.03175
R12847 vss.n3617 vss.n3071 0.03175
R12848 vss.n3650 vss.n2190 0.03175
R12849 vss.n3683 vss.n2146 0.03175
R12850 vss.n3719 vss.n2088 0.03175
R12851 vss.n3752 vss.n2034 0.03175
R12852 vss.n3785 vss.n1979 0.03175
R12853 vss.n3821 vss.n1921 0.03175
R12854 vss.n3854 vss.n1867 0.03175
R12855 vss.n3887 vss.n1812 0.03175
R12856 vss.n3923 vss.n1764 0.03175
R12857 vss.n3956 vss.n1709 0.03175
R12858 vss.n3992 vss.n1651 0.03175
R12859 vss.n4025 vss.n1597 0.03175
R12860 vss.n4058 vss.n1542 0.03175
R12861 vss.n4094 vss.n1484 0.03175
R12862 vss.n4127 vss.n1430 0.03175
R12863 vss.n4160 vss.n1386 0.03175
R12864 vss.n4196 vss.n1338 0.03175
R12865 vss.n2953 vss.n2362 0.03175
R12866 vss.n2922 vss.n26 0.03175
R12867 vss.n2918 vss.n26 0.03175
R12868 vss.n2889 vss.n2888 0.03175
R12869 vss.n2859 vss.n2606 0.03175
R12870 vss.n2829 vss.n65 0.03175
R12871 vss.n2825 vss.n65 0.03175
R12872 vss.n2796 vss.n2795 0.03175
R12873 vss.n5924 vss.n208 0.03175
R12874 vss.n5960 vss.n164 0.03175
R12875 vss.n4445 vss.n4300 0.0313824
R12876 vss.n4526 vss.n4525 0.0313824
R12877 vss.n4537 vss.n4536 0.0313824
R12878 vss.n3713 vss.n2107 0.0313277
R12879 vss.n3788 vss.n1975 0.0313277
R12880 vss.n3815 vss.n1940 0.0313277
R12881 vss.n3890 vss.n1808 0.0313277
R12882 vss.n3986 vss.n1670 0.0313277
R12883 vss.n4061 vss.n1538 0.0313277
R12884 vss.n4088 vss.n1503 0.0313277
R12885 vss.n4163 vss.n1382 0.0313277
R12886 vss.n5954 vss.n172 0.0313277
R12887 vss.n2978 vss.n2968 0.0312617
R12888 vss.n3686 vss.n2142 0.0309054
R12889 vss.n3917 vss.n1773 0.0309054
R12890 vss.n3959 vss.n1705 0.0309054
R12891 vss.n4190 vss.n1348 0.0309054
R12892 vss.n2892 vss.n39 0.0309054
R12893 vss.n2855 vss.n2613 0.0309054
R12894 vss.n5927 vss.n91 0.0309054
R12895 vss.n3644 vss.n3045 0.0304831
R12896 vss.n3746 vss.n2053 0.0304831
R12897 vss.n3857 vss.n1863 0.0304831
R12898 vss.n4019 vss.n1616 0.0304831
R12899 vss.n4130 vss.n1426 0.0304831
R12900 vss.n2949 vss.n14 0.0304831
R12901 vss.n2799 vss.n2714 0.0304831
R12902 vss.n5604 vss.n254 0.0301053
R12903 vss.n5902 vss.n239 0.0301053
R12904 vss.n5875 vss.n5657 0.0301053
R12905 vss.n5849 vss.n5693 0.0301053
R12906 vss.n5823 vss.n5732 0.0301053
R12907 vss.n3653 vss.n2186 0.0300608
R12908 vss.n3755 vss.n2030 0.0300608
R12909 vss.n3848 vss.n1886 0.0300608
R12910 vss.n4028 vss.n1593 0.0300608
R12911 vss.n4121 vss.n1449 0.0300608
R12912 vss.n2955 vss.n2954 0.0300608
R12913 vss.n2792 vss.n79 0.0300608
R12914 vss.n6012 vss.n130 0.0300608
R12915 vss.n5570 vss.n5569 0.0299698
R12916 vss.n4444 vss.n4443 0.0299118
R12917 vss.n4445 vss.n4444 0.0299118
R12918 vss.n5537 vss.n299 0.0297969
R12919 vss.n3677 vss.n2155 0.0296385
R12920 vss.n3926 vss.n1760 0.0296385
R12921 vss.n3950 vss.n1729 0.0296385
R12922 vss.n4199 vss.n1333 0.0296385
R12923 vss.n2885 vss.n40 0.0296385
R12924 vss.n2862 vss.n51 0.0296385
R12925 vss.n2316 vss.n1299 0.0293086
R12926 vss.n3722 vss.n2084 0.0292162
R12927 vss.n3779 vss.n1999 0.0292162
R12928 vss.n3824 vss.n1917 0.0292162
R12929 vss.n3881 vss.n1832 0.0292162
R12930 vss.n3995 vss.n1647 0.0292162
R12931 vss.n4052 vss.n1562 0.0292162
R12932 vss.n4097 vss.n1480 0.0292162
R12933 vss.n4154 vss.n1395 0.0292162
R12934 vss.n2768 vss.n90 0.0292162
R12935 vss.n5963 vss.n159 0.0292162
R12936 vss.n2319 vss.n1300 0.0288203
R12937 vss.n3609 vss.n3074 0.0287939
R12938 vss.n3620 vss.n3068 0.0287939
R12939 vss.n2925 vss.n25 0.0287939
R12940 vss.n2915 vss.n2506 0.0287939
R12941 vss.n2822 vss.n66 0.0287939
R12942 vss.n4450 vss.n4300 0.0284412
R12943 vss.n4527 vss.n4526 0.0284412
R12944 vss.n4536 vss.n4534 0.0284412
R12945 vss.n3710 vss.n2105 0.0283716
R12946 vss.n3791 vss.n1971 0.0283716
R12947 vss.n3812 vss.n1938 0.0283716
R12948 vss.n3893 vss.n1804 0.0283716
R12949 vss.n3983 vss.n1668 0.0283716
R12950 vss.n4064 vss.n1534 0.0283716
R12951 vss.n4085 vss.n1501 0.0283716
R12952 vss.n4166 vss.n1378 0.0283716
R12953 vss.n2832 vss.n64 0.0283716
R12954 vss.n5951 vss.n171 0.0283716
R12955 vss.n3689 vss.n2138 0.0279493
R12956 vss.n3914 vss.n1771 0.0279493
R12957 vss.n3962 vss.n1701 0.0279493
R12958 vss.n4187 vss.n1346 0.0279493
R12959 vss.n2852 vss.n54 0.0279493
R12960 vss.n5930 vss.n201 0.0279493
R12961 vss.n5584 vss.n266 0.0279123
R12962 vss.n5614 vss.n246 0.0279123
R12963 vss.n5892 vss.n5891 0.0279123
R12964 vss.n5865 vss.n5864 0.0279123
R12965 vss.n5839 vss.n5838 0.0279123
R12966 vss.n5813 vss.n5812 0.0279123
R12967 vss.n3010 vss.n2337 0.0278438
R12968 vss.n3641 vss.n3043 0.027527
R12969 vss.n3743 vss.n2051 0.027527
R12970 vss.n3860 vss.n1859 0.027527
R12971 vss.n4016 vss.n1614 0.027527
R12972 vss.n4133 vss.n1422 0.027527
R12973 vss.n2946 vss.n15 0.027527
R12974 vss.n2895 vss.n2541 0.027527
R12975 vss.n2802 vss.n76 0.027527
R12976 vss.n4384 vss.n4325 0.0274097
R12977 vss.n3011 vss.n2335 0.0273555
R12978 vss.n3758 vss.n2026 0.0271047
R12979 vss.n3845 vss.n1884 0.0271047
R12980 vss.n4031 vss.n1589 0.0271047
R12981 vss.n4118 vss.n1447 0.0271047
R12982 vss.n2789 vss.n80 0.0271047
R12983 vss.n5987 vss.n129 0.0271047
R12984 vss.n4454 vss.n4452 0.0269706
R12985 vss.n4532 vss.n4280 0.0269706
R12986 vss.n4533 vss.n4532 0.0269706
R12987 vss.n3656 vss.n2182 0.0266824
R12988 vss.n3674 vss.n2153 0.0266824
R12989 vss.n3929 vss.n1756 0.0266824
R12990 vss.n3947 vss.n1727 0.0266824
R12991 vss.n4201 vss.n4200 0.0266824
R12992 vss.n2958 vss.n11 0.0266824
R12993 vss.n2882 vss.n41 0.0266824
R12994 vss.n2865 vss.n50 0.0266824
R12995 vss.n3776 vss.n1997 0.0262601
R12996 vss.n3827 vss.n1913 0.0262601
R12997 vss.n4049 vss.n1560 0.0262601
R12998 vss.n4100 vss.n1476 0.0262601
R12999 vss.n2771 vss.n89 0.0262601
R13000 vss.n5966 vss.n154 0.0262601
R13001 vss.n3606 vss.n3079 0.0258378
R13002 vss.n3623 vss.n3065 0.0258378
R13003 vss.n3725 vss.n2080 0.0258378
R13004 vss.n3878 vss.n1830 0.0258378
R13005 vss.n3998 vss.n1643 0.0258378
R13006 vss.n4151 vss.n1393 0.0258378
R13007 vss.n2928 vss.n24 0.0258378
R13008 vss.n2912 vss.n29 0.0258378
R13009 vss.n2821 vss.n2820 0.0258378
R13010 vss.n5607 vss.n252 0.0257193
R13011 vss.n5899 vss.n5898 0.0257193
R13012 vss.n5872 vss.n5871 0.0257193
R13013 vss.n5846 vss.n5845 0.0257193
R13014 vss.n5820 vss.n5819 0.0257193
R13015 vss.n4351 vss.n4328 0.0255
R13016 vss.n4440 vss.n4302 0.0255
R13017 vss.n4451 vss.n4450 0.0255
R13018 vss.n3707 vss.n2110 0.0254155
R13019 vss.n3896 vss.n1800 0.0254155
R13020 vss.n3980 vss.n1673 0.0254155
R13021 vss.n4169 vss.n1374 0.0254155
R13022 vss.n2834 vss.n2833 0.0254155
R13023 vss.n5948 vss.n176 0.0254155
R13024 vss.n5778 vss.n109 0.0252351
R13025 vss.n3692 vss.n2134 0.0249932
R13026 vss.n3794 vss.n1967 0.0249932
R13027 vss.n3809 vss.n1943 0.0249932
R13028 vss.n3911 vss.n1776 0.0249932
R13029 vss.n3965 vss.n1697 0.0249932
R13030 vss.n4067 vss.n1530 0.0249932
R13031 vss.n4082 vss.n1506 0.0249932
R13032 vss.n4184 vss.n1351 0.0249932
R13033 vss.n2849 vss.n55 0.0249932
R13034 vss.n5933 vss.n94 0.0249932
R13035 vss.n2314 vss.n1298 0.0249141
R13036 vss.n4219 vss.n1310 0.0249141
R13037 vss.n3638 vss.n3047 0.0245709
R13038 vss.n2943 vss.n16 0.0245709
R13039 vss.n2898 vss.n36 0.0245709
R13040 vss.n2805 vss.n75 0.0245709
R13041 vss.n3740 vss.n2056 0.0241486
R13042 vss.n3761 vss.n2022 0.0241486
R13043 vss.n3842 vss.n1889 0.0241486
R13044 vss.n3863 vss.n1855 0.0241486
R13045 vss.n4013 vss.n1619 0.0241486
R13046 vss.n4034 vss.n1585 0.0241486
R13047 vss.n4115 vss.n1452 0.0241486
R13048 vss.n4136 vss.n1418 0.0241486
R13049 vss.n2786 vss.n81 0.0241486
R13050 vss.n5990 vss.n5980 0.0241486
R13051 vss.n4443 vss.n4442 0.0240294
R13052 vss.n4522 vss.n4282 0.0240294
R13053 vss.n4544 vss.n4542 0.0240294
R13054 vss.n2393 vss.n2391 0.0239375
R13055 vss.n4364 vss.n4360 0.0239375
R13056 vss.n3659 vss.n2178 0.0237264
R13057 vss.n3944 vss.n1732 0.0237264
R13058 vss.n2961 vss.n10 0.0237264
R13059 vss.n2881 vss.n2880 0.0237264
R13060 vss.n2868 vss.n49 0.0237264
R13061 vss.n5581 vss.n268 0.0235263
R13062 vss.n5610 vss.n245 0.0235263
R13063 vss.n5895 vss.n5634 0.0235263
R13064 vss.n5868 vss.n5670 0.0235263
R13065 vss.n5842 vss.n5707 0.0235263
R13066 vss.n5816 vss.n5746 0.0235263
R13067 vss.n5573 vss.n273 0.0235263
R13068 vss.n2409 vss.n2408 0.0234492
R13069 vss.n3671 vss.n2158 0.0233041
R13070 vss.n3773 vss.n2002 0.0233041
R13071 vss.n3830 vss.n1909 0.0233041
R13072 vss.n3932 vss.n1752 0.0233041
R13073 vss.n4046 vss.n1565 0.0233041
R13074 vss.n4103 vss.n1472 0.0233041
R13075 vss.n2995 vss.n4 0.0233041
R13076 vss.n2774 vss.n2760 0.0233041
R13077 vss.n6000 vss.n5967 0.0233041
R13078 vss.n4367 vss.n4366 0.0232009
R13079 vss.n4362 vss.n4361 0.0230694
R13080 vss.n3626 vss.n3062 0.0228818
R13081 vss.n3728 vss.n2076 0.0228818
R13082 vss.n3875 vss.n1835 0.0228818
R13083 vss.n4001 vss.n1639 0.0228818
R13084 vss.n4148 vss.n1398 0.0228818
R13085 vss.n2931 vss.n2480 0.0228818
R13086 vss.n2817 vss.n69 0.0228818
R13087 vss.n4385 vss.n4321 0.0226729
R13088 vss.n4392 vss.n4321 0.0226729
R13089 vss.n4462 vss.n4460 0.0225588
R13090 vss.n4525 vss.n4524 0.0225588
R13091 vss.n4537 vss.n4277 0.0225588
R13092 vss.n3603 vss.n3081 0.0224595
R13093 vss.n3704 vss.n2114 0.0224595
R13094 vss.n3899 vss.n1796 0.0224595
R13095 vss.n3977 vss.n1677 0.0224595
R13096 vss.n4172 vss.n1370 0.0224595
R13097 vss.n2909 vss.n30 0.0224595
R13098 vss.n2837 vss.n61 0.0224595
R13099 vss.n5945 vss.n180 0.0224595
R13100 vss.n5759 vss.n5753 0.022375
R13101 vss.n4574 vss.n4268 0.022375
R13102 vss.n3695 vss.n2130 0.0220372
R13103 vss.n3797 vss.n1963 0.0220372
R13104 vss.n3806 vss.n1947 0.0220372
R13105 vss.n3908 vss.n1780 0.0220372
R13106 vss.n3968 vss.n1693 0.0220372
R13107 vss.n4070 vss.n1526 0.0220372
R13108 vss.n4079 vss.n1510 0.0220372
R13109 vss.n4181 vss.n1355 0.0220372
R13110 vss.n5936 vss.n96 0.0220372
R13111 vss.n3635 vss.n3050 0.0216149
R13112 vss.n2940 vss.n2465 0.0216149
R13113 vss.n2901 vss.n35 0.0216149
R13114 vss.n2846 vss.n56 0.0216149
R13115 vss.n2808 vss.n74 0.0216149
R13116 vss.n2244 vss.n2243 0.0214961
R13117 vss.n5581 vss.n270 0.0213333
R13118 vss.n5610 vss.n250 0.0213333
R13119 vss.n5895 vss.n5629 0.0213333
R13120 vss.n5868 vss.n5664 0.0213333
R13121 vss.n5842 vss.n5702 0.0213333
R13122 vss.n5816 vss.n5741 0.0213333
R13123 vss.n3737 vss.n2060 0.0211926
R13124 vss.n3764 vss.n2018 0.0211926
R13125 vss.n3839 vss.n1893 0.0211926
R13126 vss.n3866 vss.n1851 0.0211926
R13127 vss.n4010 vss.n1623 0.0211926
R13128 vss.n4037 vss.n1581 0.0211926
R13129 vss.n4112 vss.n1456 0.0211926
R13130 vss.n4139 vss.n1414 0.0211926
R13131 vss.n5992 vss.n5991 0.0211926
R13132 vss.n4357 vss.n4355 0.0210882
R13133 vss.n4432 vss.n4431 0.0210882
R13134 vss.n4455 vss.n4297 0.0210882
R13135 vss.n2306 vss.n2230 0.0210078
R13136 vss.n2443 vss.n2442 0.0210078
R13137 vss.n5660 vss.n5659 0.0208125
R13138 vss.n4492 vss.n4491 0.0208125
R13139 vss.n3662 vss.n2174 0.0207703
R13140 vss.n3941 vss.n1736 0.0207703
R13141 vss.n3003 vss.n9 0.0207703
R13142 vss.n2877 vss.n44 0.0207703
R13143 vss.n2871 vss.n2587 0.0207703
R13144 vss.n2783 vss.n2741 0.0207703
R13145 vss.n2450 vss.n2375 0.0205195
R13146 vss.n3668 vss.n2162 0.020348
R13147 vss.n3770 vss.n2006 0.020348
R13148 vss.n3833 vss.n1905 0.020348
R13149 vss.n3935 vss.n1748 0.020348
R13150 vss.n4043 vss.n1569 0.020348
R13151 vss.n4106 vss.n1468 0.020348
R13152 vss.n2998 vss.n5 0.020348
R13153 vss.n2777 vss.n86 0.020348
R13154 vss.n2443 vss.n2380 0.0200312
R13155 vss.n3629 vss.n3059 0.0199257
R13156 vss.n3731 vss.n2072 0.0199257
R13157 vss.n3872 vss.n1839 0.0199257
R13158 vss.n4004 vss.n1635 0.0199257
R13159 vss.n4145 vss.n1402 0.0199257
R13160 vss.n2934 vss.n21 0.0199257
R13161 vss.n2814 vss.n70 0.0199257
R13162 vss.n5999 vss.n5998 0.0199257
R13163 vss.n4354 vss.n4353 0.0196176
R13164 vss.n4435 vss.n4434 0.0196176
R13165 vss.n4514 vss.n4513 0.0196176
R13166 vss.n4547 vss.n4275 0.0196176
R13167 vss.n2289 vss.n2244 0.019543
R13168 vss.n2426 vss.n2425 0.019543
R13169 vss.n3701 vss.n2118 0.0195034
R13170 vss.n3902 vss.n1792 0.0195034
R13171 vss.n3974 vss.n1681 0.0195034
R13172 vss.n4175 vss.n1366 0.0195034
R13173 vss.n2906 vss.n31 0.0195034
R13174 vss.n2840 vss.n60 0.0195034
R13175 vss.n116 vss.n99 0.019402
R13176 vss.n123 vss.n112 0.019402
R13177 vss.n118 vss.n99 0.019402
R13178 vss.n124 vss.n123 0.019402
R13179 vss.n5752 vss.n5751 0.01925
R13180 vss.n4560 vss.n4271 0.01925
R13181 vss.n3602 vss.n3601 0.0192033
R13182 vss.n6018 vss.n97 0.0191787
R13183 vss.n116 vss.n107 0.0191787
R13184 vss.n117 vss.n115 0.0191787
R13185 vss.n115 vss.n100 0.0191787
R13186 vss.n119 vss.n114 0.0191787
R13187 vss.n114 vss.n101 0.0191787
R13188 vss.n121 vss.n113 0.0191787
R13189 vss.n113 vss.n102 0.0191787
R13190 vss.n112 vss.n103 0.0191787
R13191 vss.n125 vss.n111 0.0191787
R13192 vss.n111 vss.n104 0.0191787
R13193 vss.n127 vss.n110 0.0191787
R13194 vss.n110 vss.n105 0.0191787
R13195 vss.n6014 vss.n105 0.0191787
R13196 vss.n128 vss.n104 0.0191787
R13197 vss.n126 vss.n103 0.0191787
R13198 vss.n124 vss.n102 0.0191787
R13199 vss.n122 vss.n101 0.0191787
R13200 vss.n120 vss.n100 0.0191787
R13201 vss.n128 vss.n127 0.0191787
R13202 vss.n126 vss.n125 0.0191787
R13203 vss.n122 vss.n121 0.0191787
R13204 vss.n120 vss.n119 0.0191787
R13205 vss.n118 vss.n117 0.0191787
R13206 vss.n6016 vss.n107 0.0191787
R13207 vss.n106 vss.n97 0.0191787
R13208 vss.n5607 vss.n250 0.0191404
R13209 vss.n5898 vss.n5629 0.0191404
R13210 vss.n5871 vss.n5664 0.0191404
R13211 vss.n5845 vss.n5702 0.0191404
R13212 vss.n5819 vss.n5741 0.0191404
R13213 vss.n3698 vss.n2126 0.0190811
R13214 vss.n3800 vss.n1959 0.0190811
R13215 vss.n3803 vss.n1951 0.0190811
R13216 vss.n3905 vss.n1784 0.0190811
R13217 vss.n3971 vss.n1689 0.0190811
R13218 vss.n4073 vss.n1522 0.0190811
R13219 vss.n4076 vss.n1514 0.0190811
R13220 vss.n4178 vss.n1358 0.0190811
R13221 vss.n5939 vss.n191 0.0190811
R13222 vss.n5942 vss.n184 0.0190811
R13223 vss.n2290 vss.n2240 0.0190547
R13224 vss.n3632 vss.n3053 0.0186588
R13225 vss.n2937 vss.n19 0.0186588
R13226 vss.n2904 vss.n34 0.0186588
R13227 vss.n2843 vss.n2630 0.0186588
R13228 vss.n3734 vss.n2064 0.0182365
R13229 vss.n3767 vss.n2014 0.0182365
R13230 vss.n3836 vss.n1897 0.0182365
R13231 vss.n3869 vss.n1847 0.0182365
R13232 vss.n4007 vss.n1627 0.0182365
R13233 vss.n4040 vss.n1577 0.0182365
R13234 vss.n4109 vss.n1460 0.0182365
R13235 vss.n4142 vss.n1410 0.0182365
R13236 vss.n2811 vss.n2695 0.0182365
R13237 vss.n5995 vss.n5974 0.0182365
R13238 vss.n4465 vss.n4295 0.0181471
R13239 vss.n4517 vss.n4516 0.0181471
R13240 vss.n4546 vss.n4545 0.0181471
R13241 vss.n3665 vss.n2170 0.0178142
R13242 vss.n3938 vss.n1740 0.0178142
R13243 vss.n3002 vss.n3001 0.0178142
R13244 vss.n2874 vss.n45 0.0178142
R13245 vss.n2780 vss.n84 0.0178142
R13246 vss.n5889 vss.n5888 0.0176875
R13247 vss.n4478 vss.n4291 0.0176875
R13248 vss.n3665 vss.n2166 0.0173919
R13249 vss.n3767 vss.n2010 0.0173919
R13250 vss.n3836 vss.n1901 0.0173919
R13251 vss.n3938 vss.n1744 0.0173919
R13252 vss.n4040 vss.n1573 0.0173919
R13253 vss.n4109 vss.n1464 0.0173919
R13254 vss.n3001 vss.n6 0.0173919
R13255 vss.n2874 vss.n46 0.0173919
R13256 vss.n2780 vss.n85 0.0173919
R13257 vss.n2290 vss.n2289 0.0171016
R13258 vss.n2426 vss.n2391 0.0171016
R13259 vss.n3734 vss.n2068 0.0169696
R13260 vss.n3869 vss.n1843 0.0169696
R13261 vss.n4007 vss.n1631 0.0169696
R13262 vss.n4142 vss.n1406 0.0169696
R13263 vss.n2811 vss.n71 0.0169696
R13264 vss.n5995 vss.n5969 0.0169696
R13265 vss.n5584 vss.n268 0.0169474
R13266 vss.n5614 vss.n245 0.0169474
R13267 vss.n5892 vss.n5634 0.0169474
R13268 vss.n5865 vss.n5670 0.0169474
R13269 vss.n5839 vss.n5707 0.0169474
R13270 vss.n5813 vss.n5746 0.0169474
R13271 vss.n5576 vss.n273 0.0169474
R13272 vss.n5568 vss.n269 0.0167446
R13273 vss.n4388 vss.n4386 0.0166765
R13274 vss.n4425 vss.n4424 0.0166765
R13275 vss.n4464 vss.n4463 0.0166765
R13276 vss.n2425 vss.n2380 0.0166133
R13277 vss.n3632 vss.n3056 0.0165473
R13278 vss.n3698 vss.n2122 0.0165473
R13279 vss.n3905 vss.n1788 0.0165473
R13280 vss.n3971 vss.n1685 0.0165473
R13281 vss.n4178 vss.n1362 0.0165473
R13282 vss.n2937 vss.n20 0.0165473
R13283 vss.n2905 vss.n2904 0.0165473
R13284 vss.n2843 vss.n59 0.0165473
R13285 vss.n3333 vss.n3311 0.0161667
R13286 vss.n3325 vss.n3311 0.0161667
R13287 vss.n3325 vss.n3324 0.0161667
R13288 vss.n3324 vss.n1 0.0161667
R13289 vss.n6130 vss.n1 0.0161667
R13290 vss.n5822 vss.n5737 0.016125
R13291 vss.n2450 vss.n2449 0.016125
R13292 vss.n4550 vss.n4273 0.016125
R13293 vss.n3800 vss.n1955 0.016125
R13294 vss.n3803 vss.n1955 0.016125
R13295 vss.n4073 vss.n1518 0.016125
R13296 vss.n4076 vss.n1518 0.016125
R13297 vss.n5939 vss.n108 0.016125
R13298 vss.n5942 vss.n108 0.016125
R13299 vss.n275 vss.n271 0.0159348
R13300 vss.n3629 vss.n3056 0.0157027
R13301 vss.n3701 vss.n2122 0.0157027
R13302 vss.n3902 vss.n1788 0.0157027
R13303 vss.n3974 vss.n1685 0.0157027
R13304 vss.n4175 vss.n1362 0.0157027
R13305 vss.n2934 vss.n20 0.0157027
R13306 vss.n2906 vss.n2905 0.0157027
R13307 vss.n2840 vss.n59 0.0157027
R13308 vss.n2306 vss.n2305 0.0156367
R13309 vss.n5544 vss.n295 0.0154435
R13310 vss.n4367 vss.n4363 0.0154435
R13311 vss.n4374 vss.n4363 0.0154435
R13312 vss.n4375 vss.n4374 0.0154435
R13313 vss.n3731 vss.n2068 0.0152804
R13314 vss.n3872 vss.n1843 0.0152804
R13315 vss.n4004 vss.n1631 0.0152804
R13316 vss.n4145 vss.n1406 0.0152804
R13317 vss.n2814 vss.n71 0.0152804
R13318 vss.n5998 vss.n5969 0.0152804
R13319 vss.n4358 vss.n4323 0.0152059
R13320 vss.n4430 vss.n4305 0.0152059
R13321 vss.n4507 vss.n4506 0.0152059
R13322 vss.n4556 vss.n4554 0.0152059
R13323 vss.n6015 vss.n109 0.0151515
R13324 vss.n2243 vss.n2230 0.0151484
R13325 vss.n3668 vss.n2166 0.0148581
R13326 vss.n3770 vss.n2010 0.0148581
R13327 vss.n3833 vss.n1901 0.0148581
R13328 vss.n3935 vss.n1744 0.0148581
R13329 vss.n4043 vss.n1573 0.0148581
R13330 vss.n4106 vss.n1464 0.0148581
R13331 vss.n2998 vss.n6 0.0148581
R13332 vss.n2871 vss.n46 0.0148581
R13333 vss.n2777 vss.n85 0.0148581
R13334 vss.n5604 vss.n252 0.0147544
R13335 vss.n5899 vss.n239 0.0147544
R13336 vss.n5872 vss.n5657 0.0147544
R13337 vss.n5846 vss.n5693 0.0147544
R13338 vss.n5820 vss.n5732 0.0147544
R13339 vss.n5638 vss.n5626 0.0145625
R13340 vss.n4468 vss.n4293 0.0145625
R13341 vss.n3662 vss.n2170 0.0144358
R13342 vss.n3941 vss.n1740 0.0144358
R13343 vss.n3003 vss.n3002 0.0144358
R13344 vss.n2877 vss.n45 0.0144358
R13345 vss.n2783 vss.n84 0.0144358
R13346 vss.n6118 vss.n6117 0.0144134
R13347 vss.n6106 vss.n18 0.0144134
R13348 vss.n6098 vss.n28 0.0144134
R13349 vss.n6087 vss.n6086 0.0144134
R13350 vss.n6076 vss.n6075 0.0144134
R13351 vss.n6064 vss.n53 0.0144134
R13352 vss.n6056 vss.n63 0.0144134
R13353 vss.n6045 vss.n6044 0.0144134
R13354 vss.n6034 vss.n6033 0.0144134
R13355 vss.n6022 vss.n88 0.0144134
R13356 vss.n3589 vss.n3085 0.0144134
R13357 vss.n3581 vss.n3089 0.0144134
R13358 vss.n3570 vss.n3569 0.0144134
R13359 vss.n3559 vss.n3558 0.0144134
R13360 vss.n3546 vss.n3102 0.0144134
R13361 vss.n3537 vss.n3113 0.0144134
R13362 vss.n3526 vss.n3525 0.0144134
R13363 vss.n3515 vss.n3514 0.0144134
R13364 vss.n3504 vss.n3503 0.0144134
R13365 vss.n3493 vss.n3492 0.0144134
R13366 vss.n3482 vss.n3481 0.0144134
R13367 vss.n3471 vss.n3470 0.0144134
R13368 vss.n3459 vss.n3190 0.0144134
R13369 vss.n3430 vss.n3429 0.0144134
R13370 vss.n3419 vss.n3418 0.0144134
R13371 vss.n3408 vss.n3407 0.0144134
R13372 vss.n3397 vss.n3396 0.0144134
R13373 vss.n3386 vss.n3385 0.0144134
R13374 vss.n3375 vss.n3374 0.0144134
R13375 vss.n6124 vss.n2 0.0142437
R13376 vss.n6124 vss.n6123 0.0142437
R13377 vss.n6123 vss.n6122 0.0142437
R13378 vss.n6122 vss.n8 0.0142437
R13379 vss.n6118 vss.n8 0.0142437
R13380 vss.n6117 vss.n6116 0.0142437
R13381 vss.n6116 vss.n13 0.0142437
R13382 vss.n6112 vss.n13 0.0142437
R13383 vss.n6112 vss.n6111 0.0142437
R13384 vss.n6111 vss.n6110 0.0142437
R13385 vss.n6110 vss.n18 0.0142437
R13386 vss.n6106 vss.n6105 0.0142437
R13387 vss.n6105 vss.n6104 0.0142437
R13388 vss.n6104 vss.n23 0.0142437
R13389 vss.n6100 vss.n23 0.0142437
R13390 vss.n6100 vss.n6099 0.0142437
R13391 vss.n6099 vss.n6098 0.0142437
R13392 vss.n6094 vss.n28 0.0142437
R13393 vss.n6094 vss.n6093 0.0142437
R13394 vss.n6093 vss.n6092 0.0142437
R13395 vss.n6092 vss.n33 0.0142437
R13396 vss.n6088 vss.n33 0.0142437
R13397 vss.n6088 vss.n6087 0.0142437
R13398 vss.n6086 vss.n38 0.0142437
R13399 vss.n6082 vss.n38 0.0142437
R13400 vss.n6082 vss.n6081 0.0142437
R13401 vss.n6081 vss.n6080 0.0142437
R13402 vss.n6080 vss.n43 0.0142437
R13403 vss.n6076 vss.n43 0.0142437
R13404 vss.n6075 vss.n6074 0.0142437
R13405 vss.n6074 vss.n48 0.0142437
R13406 vss.n6070 vss.n48 0.0142437
R13407 vss.n6070 vss.n6069 0.0142437
R13408 vss.n6069 vss.n6068 0.0142437
R13409 vss.n6068 vss.n53 0.0142437
R13410 vss.n6064 vss.n6063 0.0142437
R13411 vss.n6063 vss.n6062 0.0142437
R13412 vss.n6062 vss.n58 0.0142437
R13413 vss.n6058 vss.n58 0.0142437
R13414 vss.n6058 vss.n6057 0.0142437
R13415 vss.n6057 vss.n6056 0.0142437
R13416 vss.n6052 vss.n63 0.0142437
R13417 vss.n6052 vss.n6051 0.0142437
R13418 vss.n6051 vss.n6050 0.0142437
R13419 vss.n6050 vss.n68 0.0142437
R13420 vss.n6046 vss.n68 0.0142437
R13421 vss.n6046 vss.n6045 0.0142437
R13422 vss.n6044 vss.n73 0.0142437
R13423 vss.n6040 vss.n73 0.0142437
R13424 vss.n6040 vss.n6039 0.0142437
R13425 vss.n6039 vss.n6038 0.0142437
R13426 vss.n6038 vss.n78 0.0142437
R13427 vss.n6034 vss.n78 0.0142437
R13428 vss.n6033 vss.n6032 0.0142437
R13429 vss.n6032 vss.n83 0.0142437
R13430 vss.n6028 vss.n83 0.0142437
R13431 vss.n6028 vss.n6027 0.0142437
R13432 vss.n6027 vss.n6026 0.0142437
R13433 vss.n6026 vss.n88 0.0142437
R13434 vss.n6022 vss.n6021 0.0142437
R13435 vss.n6021 vss.n6020 0.0142437
R13436 vss.n3600 vss.n3599 0.0142437
R13437 vss.n3599 vss.n3083 0.0142437
R13438 vss.n3595 vss.n3083 0.0142437
R13439 vss.n3595 vss.n3594 0.0142437
R13440 vss.n3594 vss.n3593 0.0142437
R13441 vss.n3593 vss.n3085 0.0142437
R13442 vss.n3589 vss.n3588 0.0142437
R13443 vss.n3588 vss.n3587 0.0142437
R13444 vss.n3587 vss.n3087 0.0142437
R13445 vss.n3583 vss.n3087 0.0142437
R13446 vss.n3583 vss.n3582 0.0142437
R13447 vss.n3582 vss.n3581 0.0142437
R13448 vss.n3577 vss.n3089 0.0142437
R13449 vss.n3577 vss.n3576 0.0142437
R13450 vss.n3576 vss.n3575 0.0142437
R13451 vss.n3575 vss.n3091 0.0142437
R13452 vss.n3571 vss.n3091 0.0142437
R13453 vss.n3571 vss.n3570 0.0142437
R13454 vss.n3569 vss.n3093 0.0142437
R13455 vss.n3565 vss.n3093 0.0142437
R13456 vss.n3565 vss.n3564 0.0142437
R13457 vss.n3564 vss.n3563 0.0142437
R13458 vss.n3563 vss.n3095 0.0142437
R13459 vss.n3559 vss.n3095 0.0142437
R13460 vss.n3558 vss.n3557 0.0142437
R13461 vss.n3557 vss.n3097 0.0142437
R13462 vss.n3553 vss.n3097 0.0142437
R13463 vss.n3551 vss.n3550 0.0142437
R13464 vss.n3550 vss.n3102 0.0142437
R13465 vss.n3544 vss.n3543 0.0142437
R13466 vss.n3543 vss.n3107 0.0142437
R13467 vss.n3539 vss.n3538 0.0142437
R13468 vss.n3538 vss.n3537 0.0142437
R13469 vss.n3533 vss.n3532 0.0142437
R13470 vss.n3532 vss.n3531 0.0142437
R13471 vss.n3531 vss.n3119 0.0142437
R13472 vss.n3527 vss.n3526 0.0142437
R13473 vss.n3522 vss.n3521 0.0142437
R13474 vss.n3521 vss.n3520 0.0142437
R13475 vss.n3520 vss.n3130 0.0142437
R13476 vss.n3516 vss.n3515 0.0142437
R13477 vss.n3514 vss.n3136 0.0142437
R13478 vss.n3510 vss.n3509 0.0142437
R13479 vss.n3509 vss.n3508 0.0142437
R13480 vss.n3505 vss.n3504 0.0142437
R13481 vss.n3503 vss.n3147 0.0142437
R13482 vss.n3499 vss.n3498 0.0142437
R13483 vss.n3498 vss.n3497 0.0142437
R13484 vss.n3497 vss.n3153 0.0142437
R13485 vss.n3492 vss.n3491 0.0142437
R13486 vss.n3488 vss.n3487 0.0142437
R13487 vss.n3487 vss.n3486 0.0142437
R13488 vss.n3486 vss.n3164 0.0142437
R13489 vss.n3481 vss.n3480 0.0142437
R13490 vss.n3480 vss.n3170 0.0142437
R13491 vss.n3476 vss.n3475 0.0142437
R13492 vss.n3475 vss.n3474 0.0142437
R13493 vss.n3470 vss.n3469 0.0142437
R13494 vss.n3469 vss.n3181 0.0142437
R13495 vss.n3465 vss.n3464 0.0142437
R13496 vss.n3464 vss.n3463 0.0142437
R13497 vss.n3463 vss.n3190 0.0142437
R13498 vss.n3459 vss.n3458 0.0142437
R13499 vss.n3458 vss.n3457 0.0142437
R13500 vss.n3454 vss.n3453 0.0142437
R13501 vss.n3453 vss.n3452 0.0142437
R13502 vss.n3452 vss.n3197 0.0142437
R13503 vss.n3448 vss.n3447 0.0142437
R13504 vss.n3447 vss.n3446 0.0142437
R13505 vss.n3443 vss.n3442 0.0142437
R13506 vss.n3442 vss.n3441 0.0142437
R13507 vss.n3441 vss.n3208 0.0142437
R13508 vss.n3437 vss.n3436 0.0142437
R13509 vss.n3436 vss.n3435 0.0142437
R13510 vss.n3435 vss.n3214 0.0142437
R13511 vss.n3431 vss.n3430 0.0142437
R13512 vss.n3426 vss.n3425 0.0142437
R13513 vss.n3425 vss.n3424 0.0142437
R13514 vss.n3424 vss.n3225 0.0142437
R13515 vss.n3420 vss.n3419 0.0142437
R13516 vss.n3418 vss.n3231 0.0142437
R13517 vss.n3414 vss.n3413 0.0142437
R13518 vss.n3413 vss.n3412 0.0142437
R13519 vss.n3409 vss.n3408 0.0142437
R13520 vss.n3407 vss.n3242 0.0142437
R13521 vss.n3403 vss.n3402 0.0142437
R13522 vss.n3402 vss.n3401 0.0142437
R13523 vss.n3401 vss.n3248 0.0142437
R13524 vss.n3396 vss.n3395 0.0142437
R13525 vss.n3392 vss.n3391 0.0142437
R13526 vss.n3391 vss.n3390 0.0142437
R13527 vss.n3390 vss.n3259 0.0142437
R13528 vss.n3385 vss.n3384 0.0142437
R13529 vss.n3384 vss.n3265 0.0142437
R13530 vss.n3380 vss.n3379 0.0142437
R13531 vss.n3379 vss.n3378 0.0142437
R13532 vss.n3374 vss.n3373 0.0142437
R13533 vss.n3373 vss.n3276 0.0142437
R13534 vss.n3369 vss.n3368 0.0142437
R13535 vss.n3368 vss.n3367 0.0142437
R13536 vss.n3367 vss.n3282 0.0142437
R13537 vss.n3363 vss.n3362 0.0142437
R13538 vss.n3362 vss.n3361 0.0142437
R13539 vss.n3358 vss.n3357 0.0142437
R13540 vss.n3357 vss.n3356 0.0142437
R13541 vss.n3356 vss.n3293 0.0142437
R13542 vss.n3352 vss.n3351 0.0142437
R13543 vss.n3351 vss.n3350 0.0142437
R13544 vss.n3347 vss.n3346 0.0142437
R13545 vss.n3346 vss.n3345 0.0142437
R13546 vss.n3345 vss.n3304 0.0142437
R13547 vss.n3341 vss.n3340 0.0142437
R13548 vss.n3340 vss.n3339 0.0142437
R13549 vss.n3339 vss.n3308 0.0142437
R13550 vss.n3363 vss.n3287 0.014074
R13551 vss.n6128 vss.n2 0.0140468
R13552 vss.n3737 vss.n2064 0.0140135
R13553 vss.n3764 vss.n2014 0.0140135
R13554 vss.n3839 vss.n1897 0.0140135
R13555 vss.n3866 vss.n1847 0.0140135
R13556 vss.n4010 vss.n1627 0.0140135
R13557 vss.n4037 vss.n1577 0.0140135
R13558 vss.n4112 vss.n1460 0.0140135
R13559 vss.n4139 vss.n1410 0.0140135
R13560 vss.n2808 vss.n2695 0.0140135
R13561 vss.n5992 vss.n5974 0.0140135
R13562 vss.n3335 vss.n3308 0.0139483
R13563 vss.n4474 vss.n4472 0.0137353
R13564 vss.n4512 vss.n4285 0.0137353
R13565 vss.n4553 vss.n4552 0.0137353
R13566 vss.n3350 vss.n3302 0.0137347
R13567 vss.n5576 vss.n275 0.0136579
R13568 vss.n3635 vss.n3053 0.0135912
R13569 vss.n2940 vss.n19 0.0135912
R13570 vss.n2901 vss.n34 0.0135912
R13571 vss.n2846 vss.n2630 0.0135912
R13572 vss.n3476 vss.n3175 0.013565
R13573 vss.n3446 vss.n3206 0.0133953
R13574 vss.n3112 vss.n3107 0.0132256
R13575 vss.n3380 vss.n3270 0.0132256
R13576 vss.n2305 vss.n2208 0.0131953
R13577 vss.n3695 vss.n2126 0.0131689
R13578 vss.n3797 vss.n1959 0.0131689
R13579 vss.n3806 vss.n1951 0.0131689
R13580 vss.n3908 vss.n1784 0.0131689
R13581 vss.n3968 vss.n1689 0.0131689
R13582 vss.n4070 vss.n1522 0.0131689
R13583 vss.n4079 vss.n1514 0.0131689
R13584 vss.n4181 vss.n1358 0.0131689
R13585 vss.n5936 vss.n191 0.0131689
R13586 vss.n5945 vss.n184 0.0131689
R13587 vss.n5734 vss.n5715 0.013
R13588 vss.n4540 vss.n4276 0.013
R13589 vss.n3704 vss.n2118 0.0127466
R13590 vss.n3899 vss.n1792 0.0127466
R13591 vss.n3977 vss.n1681 0.0127466
R13592 vss.n4172 vss.n1366 0.0127466
R13593 vss.n2909 vss.n31 0.0127466
R13594 vss.n2837 vss.n60 0.0127466
R13595 vss.n3493 vss.n3158 0.0127166
R13596 vss.n3429 vss.n3223 0.0127166
R13597 vss.n2240 vss.n2239 0.012707
R13598 vss.n2313 vss.n2208 0.012707
R13599 vss.n2407 vss.n2337 0.012707
R13600 vss.n2409 vss.n2393 0.012707
R13601 vss.n5587 vss.n266 0.0125614
R13602 vss.n246 vss.n243 0.0125614
R13603 vss.n5891 vss.n5637 0.0125614
R13604 vss.n5864 vss.n5673 0.0125614
R13605 vss.n5838 vss.n5710 0.0125614
R13606 vss.n5812 vss.n5749 0.0125614
R13607 vss.n3331 vss.n3312 0.0123951
R13608 vss.n3525 vss.n3128 0.0123773
R13609 vss.n3397 vss.n3253 0.0123773
R13610 vss.n3626 vss.n3059 0.0123243
R13611 vss.n3728 vss.n2072 0.0123243
R13612 vss.n3875 vss.n1839 0.0123243
R13613 vss.n4001 vss.n1635 0.0123243
R13614 vss.n4148 vss.n1402 0.0123243
R13615 vss.n2931 vss.n21 0.0123243
R13616 vss.n2817 vss.n70 0.0123243
R13617 vss.n6000 vss.n5999 0.0123243
R13618 vss.n4391 vss.n4320 0.0122647
R13619 vss.n4420 vss.n4419 0.0122647
R13620 vss.n4471 vss.n4470 0.0122647
R13621 vss.n3319 vss.n3318 0.01225
R13622 vss.n2441 vss.n2375 0.0122188
R13623 vss.n6020 vss.n93 0.0122076
R13624 vss.n4385 vss.n4324 0.0120592
R13625 vss.n4394 vss.n4393 0.0120592
R13626 vss.n4394 vss.n4318 0.0120592
R13627 vss.n4400 vss.n4399 0.0120592
R13628 vss.n4400 vss.n4315 0.0120592
R13629 vss.n4408 vss.n4407 0.0120592
R13630 vss.n4408 vss.n4313 0.0120592
R13631 vss.n4359 vss.n4324 0.0120592
R13632 vss.n4393 vss.n4392 0.0120592
R13633 vss.n4399 vss.n4398 0.0120592
R13634 vss.n4407 vss.n4406 0.0120592
R13635 vss.n4398 vss.n4318 0.0120592
R13636 vss.n4406 vss.n4315 0.0120592
R13637 vss.n4413 vss.n4313 0.0120592
R13638 vss.n3510 vss.n3141 0.0120379
R13639 vss.n3412 vss.n3240 0.0120379
R13640 vss.n3671 vss.n2162 0.011902
R13641 vss.n3773 vss.n2006 0.011902
R13642 vss.n3830 vss.n1905 0.011902
R13643 vss.n3932 vss.n1748 0.011902
R13644 vss.n4046 vss.n1569 0.011902
R13645 vss.n4103 vss.n1468 0.011902
R13646 vss.n2995 vss.n5 0.011902
R13647 vss.n2774 vss.n86 0.011902
R13648 vss.n2316 vss.n1298 0.0117305
R13649 vss.n3508 vss.n3145 0.0116986
R13650 vss.n3414 vss.n3236 0.0116986
R13651 vss.n3327 vss.n3314 0.0116698
R13652 vss.n3659 vss.n2174 0.0114797
R13653 vss.n3944 vss.n1736 0.0114797
R13654 vss.n2961 vss.n9 0.0114797
R13655 vss.n2880 vss.n44 0.0114797
R13656 vss.n2868 vss.n2587 0.0114797
R13657 vss.n2786 vss.n2741 0.0114797
R13658 vss.n5624 vss.n5623 0.0114375
R13659 vss.n4458 vss.n4296 0.0114375
R13660 vss.n2314 vss.n2313 0.0112422
R13661 vss.n3527 vss.n3124 0.0111895
R13662 vss.n3395 vss.n3257 0.0111895
R13663 vss.n3322 vss.n3316 0.0110895
R13664 vss.n3740 vss.n2060 0.0110574
R13665 vss.n3761 vss.n2018 0.0110574
R13666 vss.n3842 vss.n1893 0.0110574
R13667 vss.n3863 vss.n1851 0.0110574
R13668 vss.n4013 vss.n1623 0.0110574
R13669 vss.n4034 vss.n1581 0.0110574
R13670 vss.n4115 vss.n1456 0.0110574
R13671 vss.n4136 vss.n1414 0.0110574
R13672 vss.n5991 vss.n5990 0.0110574
R13673 vss.n3491 vss.n3162 0.0108502
R13674 vss.n3431 vss.n3219 0.0108502
R13675 vss.n4390 vss.n4389 0.0107941
R13676 vss.n4423 vss.n4309 0.0107941
R13677 vss.n4502 vss.n4288 0.0107941
R13678 vss.n4564 vss.n4562 0.0107941
R13679 vss.n3638 vss.n3050 0.0106351
R13680 vss.n2943 vss.n2465 0.0106351
R13681 vss.n2898 vss.n35 0.0106351
R13682 vss.n2849 vss.n56 0.0106351
R13683 vss.n2805 vss.n74 0.0106351
R13684 vss.n3545 vss.n3544 0.0105108
R13685 vss.n3378 vss.n3274 0.0105108
R13686 vss.n5601 vss.n254 0.0103684
R13687 vss.n5903 vss.n5902 0.0103684
R13688 vss.n5876 vss.n5875 0.0103684
R13689 vss.n5850 vss.n5849 0.0103684
R13690 vss.n5824 vss.n5823 0.0103684
R13691 vss.n3448 vss.n3202 0.0103412
R13692 vss.n3692 vss.n2130 0.0102128
R13693 vss.n3794 vss.n1963 0.0102128
R13694 vss.n3809 vss.n1947 0.0102128
R13695 vss.n3911 vss.n1780 0.0102128
R13696 vss.n3965 vss.n1693 0.0102128
R13697 vss.n4067 vss.n1526 0.0102128
R13698 vss.n4082 vss.n1510 0.0102128
R13699 vss.n4184 vss.n1355 0.0102128
R13700 vss.n5933 vss.n96 0.0102128
R13701 vss.n4379 vss.n4312 0.0101931
R13702 vss.n3474 vss.n3179 0.0101715
R13703 vss.n6131 vss.n0 0.0100741
R13704 vss.n3352 vss.n3298 0.0100018
R13705 vss.n5713 vss.n5712 0.009875
R13706 vss.n4530 vss.n4278 0.009875
R13707 vss.n5798 vss.n5797 0.00986599
R13708 vss.n5797 vss.n5762 0.00986599
R13709 vss.n5793 vss.n5762 0.00986599
R13710 vss.n5793 vss.n5764 0.00986599
R13711 vss.n5789 vss.n5764 0.00986599
R13712 vss.n5789 vss.n5788 0.00986599
R13713 vss.n5788 vss.n5787 0.00986599
R13714 vss.n5787 vss.n5770 0.00986599
R13715 vss.n5783 vss.n5770 0.00986599
R13716 vss.n5783 vss.n5782 0.00986599
R13717 vss.n5782 vss.n5781 0.00986599
R13718 vss.n5781 vss.n5776 0.00986599
R13719 vss.n3606 vss.n3603 0.00979054
R13720 vss.n3707 vss.n2114 0.00979054
R13721 vss.n3896 vss.n1796 0.00979054
R13722 vss.n3980 vss.n1677 0.00979054
R13723 vss.n4169 vss.n1370 0.00979054
R13724 vss.n2912 vss.n30 0.00979054
R13725 vss.n2834 vss.n61 0.00979054
R13726 vss.n5948 vss.n180 0.00979054
R13727 vss.n3361 vss.n3291 0.00966245
R13728 vss.n3332 vss.n3310 0.00963889
R13729 vss.n5566 vss.n282 0.0095706
R13730 vss.n5546 vss.n5545 0.0095706
R13731 vss.n5566 vss.n277 0.0095706
R13732 vss.n5546 vss.n278 0.0095706
R13733 vss.n3465 vss.n3186 0.00949278
R13734 vss.n3623 vss.n3062 0.00936824
R13735 vss.n3725 vss.n2076 0.00936824
R13736 vss.n3878 vss.n1835 0.00936824
R13737 vss.n3998 vss.n1639 0.00936824
R13738 vss.n4151 vss.n1398 0.00936824
R13739 vss.n2928 vss.n2480 0.00936824
R13740 vss.n2820 vss.n69 0.00936824
R13741 vss.n4482 vss.n4480 0.00932353
R13742 vss.n4505 vss.n4504 0.00932353
R13743 vss.n4557 vss.n4272 0.00932353
R13744 vss.n3457 vss.n3195 0.00932311
R13745 vss.n2985 vss.n2335 0.00928906
R13746 vss.n3553 vss.n3552 0.00915343
R13747 vss.n3369 vss.n3281 0.00915343
R13748 vss.n5805 vss.n5803 0.00902497
R13749 vss.n3307 vss.n3304 0.00898375
R13750 vss.n3674 vss.n2158 0.00894595
R13751 vss.n3776 vss.n2002 0.00894595
R13752 vss.n3827 vss.n1909 0.00894595
R13753 vss.n3929 vss.n1752 0.00894595
R13754 vss.n4049 vss.n1565 0.00894595
R13755 vss.n4100 vss.n1472 0.00894595
R13756 vss.n4201 vss.n4 0.00894595
R13757 vss.n2771 vss.n2760 0.00894595
R13758 vss.n5967 vss.n5966 0.00894595
R13759 vss.n5794 vss.n5763 0.0088871
R13760 vss.n5796 vss.n5795 0.0088871
R13761 vss.n5795 vss.n5794 0.0088871
R13762 vss.n5767 vss.n5763 0.0088871
R13763 vss.n5768 vss.n5767 0.0088871
R13764 vss.n5769 vss.n5768 0.0088871
R13765 vss.n5772 vss.n5769 0.0088871
R13766 vss.n5773 vss.n5772 0.0088871
R13767 vss.n5774 vss.n5773 0.0088871
R13768 vss.n5775 vss.n5774 0.0088871
R13769 vss.n4219 vss.n4218 0.00880078
R13770 vss.n3011 vss.n3010 0.00880078
R13771 vss.n5538 vss.n297 0.00880078
R13772 vss.n3482 vss.n3169 0.0086444
R13773 vss.n3213 vss.n3208 0.0086444
R13774 vss.n285 vss.n281 0.00864396
R13775 vss.n288 vss.n285 0.00864396
R13776 vss.n294 vss.n289 0.00864396
R13777 vss.n291 vss.n284 0.00864396
R13778 vss.n293 vss.n292 0.00864396
R13779 vss.n5547 vss.n283 0.00864396
R13780 vss.n5567 vss.n5547 0.00864396
R13781 vss.n292 vss.n291 0.00864396
R13782 vss.n289 vss.n288 0.00864396
R13783 vss.n294 vss.n284 0.00864396
R13784 vss.n293 vss.n283 0.00864396
R13785 vss.n5569 vss.n281 0.00864396
R13786 vss.n3656 vss.n2178 0.00852365
R13787 vss.n3947 vss.n1732 0.00852365
R13788 vss.n2958 vss.n10 0.00852365
R13789 vss.n2882 vss.n2881 0.00852365
R13790 vss.n2865 vss.n49 0.00852365
R13791 vss.n290 vss.n278 0.00848752
R13792 vss.n290 vss.n282 0.00848752
R13793 vss.n3326 vss.n3315 0.00833333
R13794 vss.n5620 vss.n242 0.0083125
R13795 vss.n4448 vss.n4298 0.0083125
R13796 vss.n3118 vss.n3113 0.00830505
R13797 vss.n3386 vss.n3264 0.00830505
R13798 vss.n5591 vss.n262 0.00817544
R13799 vss.n5619 vss.n5618 0.00817544
R13800 vss.n5887 vss.n5886 0.00817544
R13801 vss.n5861 vss.n5860 0.00817544
R13802 vss.n5835 vss.n5834 0.00817544
R13803 vss.n5809 vss.n5808 0.00817544
R13804 vss.n3743 vss.n2056 0.00810135
R13805 vss.n3758 vss.n2022 0.00810135
R13806 vss.n3845 vss.n1889 0.00810135
R13807 vss.n3860 vss.n1855 0.00810135
R13808 vss.n4016 vss.n1619 0.00810135
R13809 vss.n4031 vss.n1585 0.00810135
R13810 vss.n4118 vss.n1452 0.00810135
R13811 vss.n4133 vss.n1418 0.00810135
R13812 vss.n2789 vss.n81 0.00810135
R13813 vss.n5987 vss.n5980 0.00810135
R13814 vss.n3499 vss.n3152 0.0079657
R13815 vss.n3230 vss.n3225 0.0079657
R13816 vss.n4397 vss.n4317 0.00785294
R13817 vss.n4415 vss.n4311 0.00785294
R13818 vss.n4475 vss.n4292 0.00785294
R13819 vss.n1310 vss.n1300 0.00782422
R13820 vss.n3323 vss.n3315 0.00775309
R13821 vss.n3641 vss.n3047 0.00767905
R13822 vss.n2946 vss.n16 0.00767905
R13823 vss.n2895 vss.n36 0.00767905
R13824 vss.n2802 vss.n75 0.00767905
R13825 vss.n3135 vss.n3130 0.00762635
R13826 vss.n3403 vss.n3247 0.00762635
R13827 vss.n2319 vss.n1299 0.00733594
R13828 vss.n3689 vss.n2134 0.00725676
R13829 vss.n3791 vss.n1967 0.00725676
R13830 vss.n3812 vss.n1943 0.00725676
R13831 vss.n3914 vss.n1776 0.00725676
R13832 vss.n3962 vss.n1697 0.00725676
R13833 vss.n4064 vss.n1530 0.00725676
R13834 vss.n4085 vss.n1506 0.00725676
R13835 vss.n4187 vss.n1351 0.00725676
R13836 vss.n2852 vss.n55 0.00725676
R13837 vss.n5930 vss.n94 0.00725676
R13838 vss.n3516 vss.n3135 0.00711733
R13839 vss.n3247 vss.n3242 0.00711733
R13840 vss.n6129 vss.n6128 0.00688272
R13841 vss.n2377 vss.n299 0.00684766
R13842 vss.n3710 vss.n2110 0.00683446
R13843 vss.n3893 vss.n1800 0.00683446
R13844 vss.n3983 vss.n1673 0.00683446
R13845 vss.n4166 vss.n1374 0.00683446
R13846 vss.n2833 vss.n2832 0.00683446
R13847 vss.n5951 vss.n176 0.00683446
R13848 vss.n3152 vss.n3147 0.00677798
R13849 vss.n3420 vss.n3230 0.00677798
R13850 vss.n4379 vss.n4322 0.0067601
R13851 vss.n5848 vss.n5698 0.00675
R13852 vss.n4520 vss.n4281 0.00675
R13853 vss.n3334 vss.n3310 0.00644753
R13854 vss.n3533 vss.n3118 0.00643863
R13855 vss.n3264 vss.n3259 0.00643863
R13856 vss.n3609 vss.n3079 0.00641216
R13857 vss.n3620 vss.n3065 0.00641216
R13858 vss.n3722 vss.n2080 0.00641216
R13859 vss.n3881 vss.n1830 0.00641216
R13860 vss.n3995 vss.n1643 0.00641216
R13861 vss.n4154 vss.n1393 0.00641216
R13862 vss.n2925 vss.n24 0.00641216
R13863 vss.n2915 vss.n29 0.00641216
R13864 vss.n2822 vss.n2821 0.00641216
R13865 vss.n4396 vss.n4395 0.00638235
R13866 vss.n4418 vss.n4417 0.00638235
R13867 vss.n4496 vss.n4495 0.00638235
R13868 vss.n4567 vss.n4270 0.00638235
R13869 vss.n5538 vss.n5537 0.00635938
R13870 vss.n3335 vss.n3334 0.00630247
R13871 vss.n3169 vss.n3164 0.00609928
R13872 vss.n3437 vss.n3213 0.00609928
R13873 vss.n6129 vss.n0 0.00601235
R13874 vss.n3779 vss.n1997 0.00598986
R13875 vss.n3824 vss.n1913 0.00598986
R13876 vss.n4052 vss.n1560 0.00598986
R13877 vss.n4097 vss.n1476 0.00598986
R13878 vss.n2768 vss.n89 0.00598986
R13879 vss.n5963 vss.n154 0.00598986
R13880 vss.n5598 vss.n256 0.00598246
R13881 vss.n5906 vss.n236 0.00598246
R13882 vss.n5879 vss.n5654 0.00598246
R13883 vss.n5853 vss.n5690 0.00598246
R13884 vss.n5827 vss.n5729 0.00598246
R13885 vss.n3341 vss.n3307 0.0059296
R13886 vss.n4375 vss.n4312 0.0057504
R13887 vss.n5800 vss.n5760 0.00567462
R13888 vss.n5571 vss.n276 0.00561727
R13889 vss.n3552 vss.n3551 0.00559025
R13890 vss.n3281 vss.n3276 0.00559025
R13891 vss.n3653 vss.n2182 0.00556757
R13892 vss.n3677 vss.n2153 0.00556757
R13893 vss.n3926 vss.n1756 0.00556757
R13894 vss.n3950 vss.n1727 0.00556757
R13895 vss.n4200 vss.n4199 0.00556757
R13896 vss.n2955 vss.n11 0.00556757
R13897 vss.n2885 vss.n41 0.00556757
R13898 vss.n2862 vss.n50 0.00556757
R13899 vss.n5798 vss.n5760 0.00553105
R13900 vss.n5777 vss.n5776 0.00553105
R13901 vss.n3454 vss.n3195 0.00542058
R13902 vss.n2239 vss.n2238 0.00538281
R13903 vss.n3186 vss.n3181 0.0052509
R13904 vss.n5554 vss.n5553 0.0051875
R13905 vss.n4438 vss.n4301 0.0051875
R13906 vss.n3755 vss.n2026 0.00514527
R13907 vss.n3848 vss.n1884 0.00514527
R13908 vss.n4028 vss.n1589 0.00514527
R13909 vss.n4121 vss.n1447 0.00514527
R13910 vss.n2792 vss.n80 0.00514527
R13911 vss.n130 vss.n129 0.00514527
R13912 vss.n3358 vss.n3291 0.00508123
R13913 vss.n3323 vss.n3322 0.00499691
R13914 vss.n4488 vss.n4487 0.00491176
R13915 vss.n4499 vss.n4498 0.00491176
R13916 vss.n4566 vss.n4565 0.00491176
R13917 vss.n4575 vss.n4267 0.00491176
R13918 vss.n3298 vss.n3293 0.00491155
R13919 vss.n2978 vss.n2977 0.00489453
R13920 vss.n2986 vss.n2968 0.00489453
R13921 vss.n3644 vss.n3043 0.00472297
R13922 vss.n3746 vss.n2051 0.00472297
R13923 vss.n3857 vss.n1859 0.00472297
R13924 vss.n4019 vss.n1614 0.00472297
R13925 vss.n4130 vss.n1422 0.00472297
R13926 vss.n2949 vss.n15 0.00472297
R13927 vss.n2892 vss.n2541 0.00472297
R13928 vss.n2799 vss.n76 0.00472297
R13929 vss.n3471 vss.n3179 0.0045722
R13930 vss.n3202 vss.n3197 0.0045722
R13931 vss.n3327 vss.n3326 0.00441667
R13932 vss.n3686 vss.n2138 0.00430068
R13933 vss.n3917 vss.n1771 0.00430068
R13934 vss.n3959 vss.n1701 0.00430068
R13935 vss.n4190 vss.n1346 0.00430068
R13936 vss.n2855 vss.n54 0.00430068
R13937 vss.n5927 vss.n201 0.00430068
R13938 vss.n3546 vss.n3545 0.00423285
R13939 vss.n3375 vss.n3274 0.00423285
R13940 vss.n5799 vss.n5761 0.00402161
R13941 vss.n5765 vss.n5761 0.00402161
R13942 vss.n5792 vss.n5765 0.00402161
R13943 vss.n5792 vss.n5791 0.00402161
R13944 vss.n5791 vss.n5790 0.00402161
R13945 vss.n5790 vss.n5766 0.00402161
R13946 vss.n5786 vss.n5766 0.00402161
R13947 vss.n5786 vss.n5785 0.00402161
R13948 vss.n5785 vss.n5784 0.00402161
R13949 vss.n5784 vss.n5771 0.00402161
R13950 vss.n5780 vss.n5771 0.00402161
R13951 vss.n5780 vss.n5779 0.00402103
R13952 vss.n5779 vss.n5778 0.00401908
R13953 vss.n4366 vss.n298 0.00401879
R13954 vss.n6015 vss.n93 0.00398524
R13955 vss.n4214 vss.n1312 0.00391797
R13956 vss.n2442 vss.n2441 0.00391797
R13957 vss.n3488 vss.n3162 0.0038935
R13958 vss.n3219 vss.n3214 0.0038935
R13959 vss.n3713 vss.n2105 0.00387838
R13960 vss.n3788 vss.n1971 0.00387838
R13961 vss.n3815 vss.n1938 0.00387838
R13962 vss.n3890 vss.n1804 0.00387838
R13963 vss.n3986 vss.n1668 0.00387838
R13964 vss.n4061 vss.n1534 0.00387838
R13965 vss.n4088 vss.n1501 0.00387838
R13966 vss.n4163 vss.n1378 0.00387838
R13967 vss.n2829 vss.n64 0.00387838
R13968 vss.n5954 vss.n171 0.00387838
R13969 vss.n264 vss.n260 0.00378947
R13970 vss.n5910 vss.n228 0.00378947
R13971 vss.n5883 vss.n5644 0.00378947
R13972 vss.n5857 vss.n5680 0.00378947
R13973 vss.n5831 vss.n5718 0.00378947
R13974 vss.n5805 vss.n5756 0.00378947
R13975 vss.n5695 vss.n5677 0.003625
R13976 vss.n4510 vss.n4283 0.003625
R13977 vss.n3124 vss.n3119 0.00355415
R13978 vss.n3392 vss.n3257 0.00355415
R13979 vss.n3613 vss.n3074 0.00345608
R13980 vss.n3617 vss.n3068 0.00345608
R13981 vss.n2922 vss.n25 0.00345608
R13982 vss.n2918 vss.n2506 0.00345608
R13983 vss.n2825 vss.n66 0.00345608
R13984 vss.n4405 vss.n4404 0.00344118
R13985 vss.n4409 vss.n4314 0.00344118
R13986 vss.n4484 vss.n4483 0.00344118
R13987 vss.n4218 vss.n4217 0.00342969
R13988 vss.n3332 vss.n3331 0.00311111
R13989 vss.n3505 vss.n3145 0.00304513
R13990 vss.n3236 vss.n3231 0.00304513
R13991 vss.n3719 vss.n2084 0.00303378
R13992 vss.n1999 vss.n1979 0.00303378
R13993 vss.n3821 vss.n1917 0.00303378
R13994 vss.n1832 vss.n1812 0.00303378
R13995 vss.n3992 vss.n1647 0.00303378
R13996 vss.n1562 vss.n1542 0.00303378
R13997 vss.n4094 vss.n1480 0.00303378
R13998 vss.n1395 vss.n1386 0.00303378
R13999 vss.n208 vss.n90 0.00303378
R14000 vss.n5960 vss.n159 0.00303378
R14001 vss.n98 vss.n95 0.00275863
R14002 vss.n6017 vss.n98 0.00275863
R14003 vss.n3141 vss.n3136 0.00270578
R14004 vss.n3409 vss.n3240 0.00270578
R14005 vss.n2155 vss.n2146 0.00261149
R14006 vss.n3923 vss.n1760 0.00261149
R14007 vss.n1729 vss.n1709 0.00261149
R14008 vss.n4196 vss.n1333 0.00261149
R14009 vss.n2888 vss.n40 0.00261149
R14010 vss.n2859 vss.n51 0.00261149
R14011 vss.n3522 vss.n3128 0.00236643
R14012 vss.n3253 vss.n3248 0.00236643
R14013 vss.n3650 vss.n2186 0.00218919
R14014 vss.n3752 vss.n2030 0.00218919
R14015 vss.n1886 vss.n1867 0.00218919
R14016 vss.n4025 vss.n1593 0.00218919
R14017 vss.n1449 vss.n1430 0.00218919
R14018 vss.n2954 vss.n2953 0.00218919
R14019 vss.n2795 vss.n79 0.00218919
R14020 vss.n6012 vss.n6011 0.00218919
R14021 vss.n3318 vss 0.00209568
R14022 vss.n5562 vss.n5561 0.0020625
R14023 vss.n5558 vss.n5557 0.0020625
R14024 vss.n4422 vss.n4307 0.0020625
R14025 vss.n4428 vss.n4303 0.0020625
R14026 vss.n3158 vss.n3153 0.00202708
R14027 vss.n3426 vss.n3223 0.00202708
R14028 vss.n4402 vss.n4401 0.00197059
R14029 vss.n4412 vss.n4411 0.00197059
R14030 vss.n4485 vss.n4290 0.00197059
R14031 vss.n4573 vss.n4572 0.00197059
R14032 vss.n3045 vss.n2190 0.00176689
R14033 vss.n2053 vss.n2034 0.00176689
R14034 vss.n3854 vss.n1863 0.00176689
R14035 vss.n1616 vss.n1597 0.00176689
R14036 vss.n4127 vss.n1426 0.00176689
R14037 vss.n2362 vss.n14 0.00176689
R14038 vss.n2796 vss.n2714 0.00176689
R14039 vss.n3319 vss.n3316 0.00166049
R14040 vss.n5595 vss.n258 0.00159649
R14041 vss.n233 vss.n230 0.00159649
R14042 vss.n5651 vss.n5649 0.00159649
R14043 vss.n5687 vss.n5685 0.00159649
R14044 vss.n5726 vss.n5724 0.00159649
R14045 vss.n280 vss.n279 0.00158696
R14046 vss.n3539 vss.n3112 0.00151805
R14047 vss.n3270 vss.n3265 0.00151805
R14048 vss.n4213 vss.n1315 0.00147656
R14049 vss.n3443 vss.n3206 0.00134837
R14050 vss.n3683 vss.n2142 0.00134459
R14051 vss.n1773 vss.n1764 0.00134459
R14052 vss.n3956 vss.n1705 0.00134459
R14053 vss.n1348 vss.n1338 0.00134459
R14054 vss.n2889 vss.n39 0.00134459
R14055 vss.n2613 vss.n2606 0.00134459
R14056 vss.n5924 vss.n91 0.00134459
R14057 vss.n5578 vss.n271 0.00130979
R14058 vss.n287 vss.n286 0.00130979
R14059 vss.n3175 vss.n3170 0.0011787
R14060 vss.n5568 vss.n287 0.00115217
R14061 vss.n287 vss.n275 0.00115217
R14062 vss.n280 vss.n271 0.00115217
R14063 vss.n3314 vss.n3312 0.00108025
R14064 vss.n6131 vss 0.00108025
R14065 vss.n3347 vss.n3302 0.00100902
R14066 vss.n4210 vss.n4209 0.000988281
R14067 vss.n2977 vss.n1318 0.000988281
R14068 vss.n2408 vss.n2407 0.000988281
R14069 vss.n2107 vss.n2088 0.000922297
R14070 vss.n3785 vss.n1975 0.000922297
R14071 vss.n1940 vss.n1921 0.000922297
R14072 vss.n3887 vss.n1808 0.000922297
R14073 vss.n1670 vss.n1651 0.000922297
R14074 vss.n4058 vss.n1538 0.000922297
R14075 vss.n1503 vss.n1484 0.000922297
R14076 vss.n4160 vss.n1382 0.000922297
R14077 vss.n172 vss.n164 0.000922297
R14078 vss.n3287 vss.n3282 0.00083935
R14079 vss.n6017 vss.n93 0.000533837
R14080 vin_n.n196 vin_n.t133 321.697
R14081 vin_n.n196 vin_n.t130 321.697
R14082 vin_n.n194 vin_n.t136 321.697
R14083 vin_n.n194 vin_n.t135 321.697
R14084 vin_n.n192 vin_n.t119 321.697
R14085 vin_n.n192 vin_n.t117 321.697
R14086 vin_n.n190 vin_n.t191 321.697
R14087 vin_n.n190 vin_n.t189 321.697
R14088 vin_n.n188 vin_n.t45 321.697
R14089 vin_n.n188 vin_n.t44 321.697
R14090 vin_n.n186 vin_n.t51 321.697
R14091 vin_n.n186 vin_n.t49 321.697
R14092 vin_n.n184 vin_n.t55 321.697
R14093 vin_n.n184 vin_n.t53 321.697
R14094 vin_n.n182 vin_n.t61 321.697
R14095 vin_n.n182 vin_n.t59 321.697
R14096 vin_n.n180 vin_n.t128 321.697
R14097 vin_n.n180 vin_n.t127 321.697
R14098 vin_n.n178 vin_n.t186 321.697
R14099 vin_n.n178 vin_n.t185 321.697
R14100 vin_n.n176 vin_n.t173 321.697
R14101 vin_n.n176 vin_n.t170 321.697
R14102 vin_n.n174 vin_n.t177 321.697
R14103 vin_n.n174 vin_n.t176 321.697
R14104 vin_n.n172 vin_n.t180 321.697
R14105 vin_n.n172 vin_n.t179 321.697
R14106 vin_n.n170 vin_n.t182 321.697
R14107 vin_n.n170 vin_n.t181 321.697
R14108 vin_n.n168 vin_n.t99 321.697
R14109 vin_n.n168 vin_n.t98 321.697
R14110 vin_n.n166 vin_n.t103 321.697
R14111 vin_n.n166 vin_n.t102 321.697
R14112 vin_n.n164 vin_n.t108 321.697
R14113 vin_n.n164 vin_n.t106 321.697
R14114 vin_n.n162 vin_n.t112 321.697
R14115 vin_n.n162 vin_n.t110 321.697
R14116 vin_n.n160 vin_n.t120 321.697
R14117 vin_n.n160 vin_n.t118 321.697
R14118 vin_n.n158 vin_n.t157 321.697
R14119 vin_n.n158 vin_n.t155 321.697
R14120 vin_n.n156 vin_n.t19 321.697
R14121 vin_n.n156 vin_n.t17 321.697
R14122 vin_n.n154 vin_n.t27 321.697
R14123 vin_n.n154 vin_n.t26 321.697
R14124 vin_n.n152 vin_n.t32 321.697
R14125 vin_n.n152 vin_n.t31 321.697
R14126 vin_n.n150 vin_n.t40 321.697
R14127 vin_n.n150 vin_n.t38 321.697
R14128 vin_n.n148 vin_n.t87 321.697
R14129 vin_n.n148 vin_n.t86 321.697
R14130 vin_n.n146 vin_n.t169 321.697
R14131 vin_n.n146 vin_n.t167 321.697
R14132 vin_n.n144 vin_n.t174 321.697
R14133 vin_n.n144 vin_n.t171 321.697
R14134 vin_n.n142 vin_n.t151 321.697
R14135 vin_n.n142 vin_n.t148 321.697
R14136 vin_n.n140 vin_n.t160 321.697
R14137 vin_n.n140 vin_n.t159 321.697
R14138 vin_n.n138 vin_n.t3 321.697
R14139 vin_n.n138 vin_n.t1 321.697
R14140 vin_n.n136 vin_n.t7 321.697
R14141 vin_n.n136 vin_n.t6 321.697
R14142 vin_n.n134 vin_n.t81 321.697
R14143 vin_n.n134 vin_n.t79 321.697
R14144 vin_n.n132 vin_n.t84 321.697
R14145 vin_n.n132 vin_n.t82 321.697
R14146 vin_n.n130 vin_n.t91 321.697
R14147 vin_n.n130 vin_n.t89 321.697
R14148 vin_n.n128 vin_n.t145 321.697
R14149 vin_n.n128 vin_n.t144 321.697
R14150 vin_n.n126 vin_n.t158 321.697
R14151 vin_n.n126 vin_n.t156 321.697
R14152 vin_n.n124 vin_n.t197 321.697
R14153 vin_n.n124 vin_n.t196 321.697
R14154 vin_n.n122 vin_n.t199 321.697
R14155 vin_n.n122 vin_n.t198 321.697
R14156 vin_n.n120 vin_n.t5 321.697
R14157 vin_n.n120 vin_n.t4 321.697
R14158 vin_n.n118 vin_n.t65 321.697
R14159 vin_n.n118 vin_n.t64 321.697
R14160 vin_n.n116 vin_n.t69 321.697
R14161 vin_n.n116 vin_n.t68 321.697
R14162 vin_n.n114 vin_n.t71 321.697
R14163 vin_n.n114 vin_n.t70 321.697
R14164 vin_n.n112 vin_n.t143 321.697
R14165 vin_n.n112 vin_n.t141 321.697
R14166 vin_n.n110 vin_n.t153 321.697
R14167 vin_n.n110 vin_n.t149 321.697
R14168 vin_n.n108 vin_n.t15 321.697
R14169 vin_n.n108 vin_n.t13 321.697
R14170 vin_n.n106 vin_n.t23 321.697
R14171 vin_n.n106 vin_n.t20 321.697
R14172 vin_n.n104 vin_n.t29 321.697
R14173 vin_n.n104 vin_n.t28 321.697
R14174 vin_n.n102 vin_n.t96 321.697
R14175 vin_n.n102 vin_n.t95 321.697
R14176 vin_n.n100 vin_n.t101 321.697
R14177 vin_n.n100 vin_n.t100 321.697
R14178 vin_n.n99 vin_n.t166 321.697
R14179 vin_n.n99 vin_n.t165 321.697
R14180 vin_n.n97 vin_n.t42 321.697
R14181 vin_n.n97 vin_n.t147 321.697
R14182 vin_n.n95 vin_n.t0 321.697
R14183 vin_n.n95 vin_n.t77 321.697
R14184 vin_n.n93 vin_n.t121 321.697
R14185 vin_n.n93 vin_n.t80 321.697
R14186 vin_n.n91 vin_n.t139 321.697
R14187 vin_n.n91 vin_n.t175 321.697
R14188 vin_n.n89 vin_n.t113 321.697
R14189 vin_n.n89 vin_n.t50 321.697
R14190 vin_n.n87 vin_n.t76 321.697
R14191 vin_n.n87 vin_n.t184 321.697
R14192 vin_n.n85 vin_n.t47 321.697
R14193 vin_n.n85 vin_n.t116 321.697
R14194 vin_n.n83 vin_n.t8 321.697
R14195 vin_n.n83 vin_n.t52 321.697
R14196 vin_n.n81 vin_n.t35 321.697
R14197 vin_n.n81 vin_n.t134 321.697
R14198 vin_n.n79 vin_n.t2 321.697
R14199 vin_n.n79 vin_n.t12 321.697
R14200 vin_n.n77 vin_n.t123 321.697
R14201 vin_n.n77 vin_n.t14 321.697
R14202 vin_n.n75 vin_n.t85 321.697
R14203 vin_n.n75 vin_n.t161 321.697
R14204 vin_n.n73 vin_n.t56 321.697
R14205 vin_n.n73 vin_n.t83 321.697
R14206 vin_n.n71 vin_n.t18 321.697
R14207 vin_n.n71 vin_n.t16 321.697
R14208 vin_n.n69 vin_n.t48 321.697
R14209 vin_n.n69 vin_n.t54 321.697
R14210 vin_n.n67 vin_n.t10 321.697
R14211 vin_n.n67 vin_n.t187 321.697
R14212 vin_n.n65 vin_n.t183 321.697
R14213 vin_n.n65 vin_n.t122 321.697
R14214 vin_n.n63 vin_n.t150 321.697
R14215 vin_n.n63 vin_n.t57 321.697
R14216 vin_n.n61 vin_n.t111 321.697
R14217 vin_n.n61 vin_n.t188 321.697
R14218 vin_n.n59 vin_n.t41 321.697
R14219 vin_n.n59 vin_n.t138 321.697
R14220 vin_n.n57 vin_n.t58 321.697
R14221 vin_n.n57 vin_n.t22 321.697
R14222 vin_n.n55 vin_n.t21 321.697
R14223 vin_n.n55 vin_n.t164 321.697
R14224 vin_n.n53 vin_n.t190 321.697
R14225 vin_n.n53 vin_n.t90 321.697
R14226 vin_n.n51 vin_n.t162 321.697
R14227 vin_n.n51 vin_n.t25 321.697
R14228 vin_n.n49 vin_n.t129 321.697
R14229 vin_n.n49 vin_n.t105 321.697
R14230 vin_n.n47 vin_n.t154 321.697
R14231 vin_n.n47 vin_n.t192 321.697
R14232 vin_n.n45 vin_n.t115 321.697
R14233 vin_n.n45 vin_n.t125 321.697
R14234 vin_n.n43 vin_n.t34 321.697
R14235 vin_n.n43 vin_n.t126 321.697
R14236 vin_n.n41 vin_n.t194 321.697
R14237 vin_n.n41 vin_n.t63 321.697
R14238 vin_n.n39 vin_n.t178 321.697
R14239 vin_n.n39 vin_n.t142 321.697
R14240 vin_n.n37 vin_n.t137 321.697
R14241 vin_n.n37 vin_n.t74 321.697
R14242 vin_n.n35 vin_n.t163 321.697
R14243 vin_n.n35 vin_n.t168 321.697
R14244 vin_n.n33 vin_n.t124 321.697
R14245 vin_n.n33 vin_n.t93 321.697
R14246 vin_n.n31 vin_n.t88 321.697
R14247 vin_n.n31 vin_n.t30 321.697
R14248 vin_n.n29 vin_n.t66 321.697
R14249 vin_n.n29 vin_n.t109 321.697
R14250 vin_n.n27 vin_n.t33 321.697
R14251 vin_n.n27 vin_n.t46 321.697
R14252 vin_n.n25 vin_n.t195 321.697
R14253 vin_n.n25 vin_n.t193 321.697
R14254 vin_n.n23 vin_n.t172 321.697
R14255 vin_n.n23 vin_n.t132 321.697
R14256 vin_n.n21 vin_n.t131 321.697
R14257 vin_n.n21 vin_n.t67 321.697
R14258 vin_n.n19 vin_n.t104 321.697
R14259 vin_n.n19 vin_n.t152 321.697
R14260 vin_n.n17 vin_n.t72 321.697
R14261 vin_n.n17 vin_n.t78 321.697
R14262 vin_n.n15 vin_n.t43 321.697
R14263 vin_n.n15 vin_n.t11 321.697
R14264 vin_n.n13 vin_n.t60 321.697
R14265 vin_n.n13 vin_n.t97 321.697
R14266 vin_n.n11 vin_n.t24 321.697
R14267 vin_n.n11 vin_n.t37 321.697
R14268 vin_n.n9 vin_n.t140 321.697
R14269 vin_n.n9 vin_n.t146 321.697
R14270 vin_n.n7 vin_n.t107 321.697
R14271 vin_n.n7 vin_n.t75 321.697
R14272 vin_n.n5 vin_n.t73 321.697
R14273 vin_n.n5 vin_n.t9 321.697
R14274 vin_n.n3 vin_n.t92 321.697
R14275 vin_n.n3 vin_n.t94 321.697
R14276 vin_n.n1 vin_n.t62 321.697
R14277 vin_n.n1 vin_n.t36 321.697
R14278 vin_n.n0 vin_n.t39 321.697
R14279 vin_n.n0 vin_n.t114 321.697
R14280 vin_n.n101 vin_n.n99 67.1865
R14281 vin_n.n2 vin_n.n0 67.1865
R14282 vin_n.n197 vin_n.n196 67.0982
R14283 vin_n.n195 vin_n.n194 67.0982
R14284 vin_n.n193 vin_n.n192 67.0982
R14285 vin_n.n191 vin_n.n190 67.0982
R14286 vin_n.n189 vin_n.n188 67.0982
R14287 vin_n.n187 vin_n.n186 67.0982
R14288 vin_n.n185 vin_n.n184 67.0982
R14289 vin_n.n183 vin_n.n182 67.0982
R14290 vin_n.n181 vin_n.n180 67.0982
R14291 vin_n.n179 vin_n.n178 67.0982
R14292 vin_n.n177 vin_n.n176 67.0982
R14293 vin_n.n175 vin_n.n174 67.0982
R14294 vin_n.n173 vin_n.n172 67.0982
R14295 vin_n.n171 vin_n.n170 67.0982
R14296 vin_n.n169 vin_n.n168 67.0982
R14297 vin_n.n167 vin_n.n166 67.0982
R14298 vin_n.n165 vin_n.n164 67.0982
R14299 vin_n.n163 vin_n.n162 67.0982
R14300 vin_n.n161 vin_n.n160 67.0982
R14301 vin_n.n159 vin_n.n158 67.0982
R14302 vin_n.n157 vin_n.n156 67.0982
R14303 vin_n.n155 vin_n.n154 67.0982
R14304 vin_n.n153 vin_n.n152 67.0982
R14305 vin_n.n151 vin_n.n150 67.0982
R14306 vin_n.n149 vin_n.n148 67.0982
R14307 vin_n.n147 vin_n.n146 67.0982
R14308 vin_n.n145 vin_n.n144 67.0982
R14309 vin_n.n143 vin_n.n142 67.0982
R14310 vin_n.n141 vin_n.n140 67.0982
R14311 vin_n.n139 vin_n.n138 67.0982
R14312 vin_n.n137 vin_n.n136 67.0982
R14313 vin_n.n135 vin_n.n134 67.0982
R14314 vin_n.n133 vin_n.n132 67.0982
R14315 vin_n.n131 vin_n.n130 67.0982
R14316 vin_n.n129 vin_n.n128 67.0982
R14317 vin_n.n127 vin_n.n126 67.0982
R14318 vin_n.n125 vin_n.n124 67.0982
R14319 vin_n.n123 vin_n.n122 67.0982
R14320 vin_n.n121 vin_n.n120 67.0982
R14321 vin_n.n119 vin_n.n118 67.0982
R14322 vin_n.n117 vin_n.n116 67.0982
R14323 vin_n.n115 vin_n.n114 67.0982
R14324 vin_n.n113 vin_n.n112 67.0982
R14325 vin_n.n111 vin_n.n110 67.0982
R14326 vin_n.n109 vin_n.n108 67.0982
R14327 vin_n.n107 vin_n.n106 67.0982
R14328 vin_n.n105 vin_n.n104 67.0982
R14329 vin_n.n103 vin_n.n102 67.0982
R14330 vin_n.n101 vin_n.n100 67.0982
R14331 vin_n.n98 vin_n.n97 67.0982
R14332 vin_n.n96 vin_n.n95 67.0982
R14333 vin_n.n94 vin_n.n93 67.0982
R14334 vin_n.n92 vin_n.n91 67.0982
R14335 vin_n.n90 vin_n.n89 67.0982
R14336 vin_n.n88 vin_n.n87 67.0982
R14337 vin_n.n86 vin_n.n85 67.0982
R14338 vin_n.n84 vin_n.n83 67.0982
R14339 vin_n.n82 vin_n.n81 67.0982
R14340 vin_n.n80 vin_n.n79 67.0982
R14341 vin_n.n78 vin_n.n77 67.0982
R14342 vin_n.n76 vin_n.n75 67.0982
R14343 vin_n.n74 vin_n.n73 67.0982
R14344 vin_n.n72 vin_n.n71 67.0982
R14345 vin_n.n70 vin_n.n69 67.0982
R14346 vin_n.n68 vin_n.n67 67.0982
R14347 vin_n.n66 vin_n.n65 67.0982
R14348 vin_n.n64 vin_n.n63 67.0982
R14349 vin_n.n62 vin_n.n61 67.0982
R14350 vin_n.n60 vin_n.n59 67.0982
R14351 vin_n.n58 vin_n.n57 67.0982
R14352 vin_n.n56 vin_n.n55 67.0982
R14353 vin_n.n54 vin_n.n53 67.0982
R14354 vin_n.n52 vin_n.n51 67.0982
R14355 vin_n.n50 vin_n.n49 67.0982
R14356 vin_n.n48 vin_n.n47 67.0982
R14357 vin_n.n46 vin_n.n45 67.0982
R14358 vin_n.n44 vin_n.n43 67.0982
R14359 vin_n.n42 vin_n.n41 67.0982
R14360 vin_n.n40 vin_n.n39 67.0982
R14361 vin_n.n38 vin_n.n37 67.0982
R14362 vin_n.n36 vin_n.n35 67.0982
R14363 vin_n.n34 vin_n.n33 67.0982
R14364 vin_n.n32 vin_n.n31 67.0982
R14365 vin_n.n30 vin_n.n29 67.0982
R14366 vin_n.n28 vin_n.n27 67.0982
R14367 vin_n.n26 vin_n.n25 67.0982
R14368 vin_n.n24 vin_n.n23 67.0982
R14369 vin_n.n22 vin_n.n21 67.0982
R14370 vin_n.n20 vin_n.n19 67.0982
R14371 vin_n.n18 vin_n.n17 67.0982
R14372 vin_n.n16 vin_n.n15 67.0982
R14373 vin_n.n14 vin_n.n13 67.0982
R14374 vin_n.n12 vin_n.n11 67.0982
R14375 vin_n.n10 vin_n.n9 67.0982
R14376 vin_n.n8 vin_n.n7 67.0982
R14377 vin_n.n6 vin_n.n5 67.0982
R14378 vin_n.n4 vin_n.n3 67.0982
R14379 vin_n.n2 vin_n.n1 67.0982
R14380 vin_n.n198 vin_n.n98 1.1048
R14381 vin_n.n198 vin_n.n197 1.10331
R14382 vin_n vin_n.n198 0.59929
R14383 vin_n.n103 vin_n.n101 0.0888234
R14384 vin_n.n105 vin_n.n103 0.0888234
R14385 vin_n.n107 vin_n.n105 0.0888234
R14386 vin_n.n109 vin_n.n107 0.0888234
R14387 vin_n.n111 vin_n.n109 0.0888234
R14388 vin_n.n113 vin_n.n111 0.0888234
R14389 vin_n.n115 vin_n.n113 0.0888234
R14390 vin_n.n117 vin_n.n115 0.0888234
R14391 vin_n.n119 vin_n.n117 0.0888234
R14392 vin_n.n121 vin_n.n119 0.0888234
R14393 vin_n.n123 vin_n.n121 0.0888234
R14394 vin_n.n125 vin_n.n123 0.0888234
R14395 vin_n.n127 vin_n.n125 0.0888234
R14396 vin_n.n129 vin_n.n127 0.0888234
R14397 vin_n.n131 vin_n.n129 0.0888234
R14398 vin_n.n133 vin_n.n131 0.0888234
R14399 vin_n.n135 vin_n.n133 0.0888234
R14400 vin_n.n137 vin_n.n135 0.0888234
R14401 vin_n.n139 vin_n.n137 0.0888234
R14402 vin_n.n141 vin_n.n139 0.0888234
R14403 vin_n.n143 vin_n.n141 0.0888234
R14404 vin_n.n145 vin_n.n143 0.0888234
R14405 vin_n.n147 vin_n.n145 0.0888234
R14406 vin_n.n149 vin_n.n147 0.0888234
R14407 vin_n.n151 vin_n.n149 0.0888234
R14408 vin_n.n153 vin_n.n151 0.0888234
R14409 vin_n.n155 vin_n.n153 0.0888234
R14410 vin_n.n157 vin_n.n155 0.0888234
R14411 vin_n.n159 vin_n.n157 0.0888234
R14412 vin_n.n161 vin_n.n159 0.0888234
R14413 vin_n.n163 vin_n.n161 0.0888234
R14414 vin_n.n165 vin_n.n163 0.0888234
R14415 vin_n.n167 vin_n.n165 0.0888234
R14416 vin_n.n169 vin_n.n167 0.0888234
R14417 vin_n.n171 vin_n.n169 0.0888234
R14418 vin_n.n173 vin_n.n171 0.0888234
R14419 vin_n.n175 vin_n.n173 0.0888234
R14420 vin_n.n177 vin_n.n175 0.0888234
R14421 vin_n.n179 vin_n.n177 0.0888234
R14422 vin_n.n181 vin_n.n179 0.0888234
R14423 vin_n.n183 vin_n.n181 0.0888234
R14424 vin_n.n185 vin_n.n183 0.0888234
R14425 vin_n.n187 vin_n.n185 0.0888234
R14426 vin_n.n189 vin_n.n187 0.0888234
R14427 vin_n.n191 vin_n.n189 0.0888234
R14428 vin_n.n193 vin_n.n191 0.0888234
R14429 vin_n.n195 vin_n.n193 0.0888234
R14430 vin_n.n197 vin_n.n195 0.0888234
R14431 vin_n.n4 vin_n.n2 0.0888234
R14432 vin_n.n6 vin_n.n4 0.0888234
R14433 vin_n.n8 vin_n.n6 0.0888234
R14434 vin_n.n10 vin_n.n8 0.0888234
R14435 vin_n.n12 vin_n.n10 0.0888234
R14436 vin_n.n14 vin_n.n12 0.0888234
R14437 vin_n.n16 vin_n.n14 0.0888234
R14438 vin_n.n18 vin_n.n16 0.0888234
R14439 vin_n.n20 vin_n.n18 0.0888234
R14440 vin_n.n22 vin_n.n20 0.0888234
R14441 vin_n.n24 vin_n.n22 0.0888234
R14442 vin_n.n26 vin_n.n24 0.0888234
R14443 vin_n.n28 vin_n.n26 0.0888234
R14444 vin_n.n30 vin_n.n28 0.0888234
R14445 vin_n.n32 vin_n.n30 0.0888234
R14446 vin_n.n34 vin_n.n32 0.0888234
R14447 vin_n.n36 vin_n.n34 0.0888234
R14448 vin_n.n38 vin_n.n36 0.0888234
R14449 vin_n.n40 vin_n.n38 0.0888234
R14450 vin_n.n42 vin_n.n40 0.0888234
R14451 vin_n.n44 vin_n.n42 0.0888234
R14452 vin_n.n46 vin_n.n44 0.0888234
R14453 vin_n.n48 vin_n.n46 0.0888234
R14454 vin_n.n50 vin_n.n48 0.0888234
R14455 vin_n.n52 vin_n.n50 0.0888234
R14456 vin_n.n54 vin_n.n52 0.0888234
R14457 vin_n.n56 vin_n.n54 0.0888234
R14458 vin_n.n58 vin_n.n56 0.0888234
R14459 vin_n.n60 vin_n.n58 0.0888234
R14460 vin_n.n62 vin_n.n60 0.0888234
R14461 vin_n.n64 vin_n.n62 0.0888234
R14462 vin_n.n66 vin_n.n64 0.0888234
R14463 vin_n.n68 vin_n.n66 0.0888234
R14464 vin_n.n70 vin_n.n68 0.0888234
R14465 vin_n.n72 vin_n.n70 0.0888234
R14466 vin_n.n74 vin_n.n72 0.0888234
R14467 vin_n.n76 vin_n.n74 0.0888234
R14468 vin_n.n78 vin_n.n76 0.0888234
R14469 vin_n.n80 vin_n.n78 0.0888234
R14470 vin_n.n82 vin_n.n80 0.0888234
R14471 vin_n.n84 vin_n.n82 0.0888234
R14472 vin_n.n86 vin_n.n84 0.0888234
R14473 vin_n.n88 vin_n.n86 0.0888234
R14474 vin_n.n90 vin_n.n88 0.0888234
R14475 vin_n.n92 vin_n.n90 0.0888234
R14476 vin_n.n94 vin_n.n92 0.0888234
R14477 vin_n.n96 vin_n.n94 0.0888234
R14478 vin_n.n98 vin_n.n96 0.0888234
R14479 vbn.n228 vbn.t40 314.466
R14480 vbn.n228 vbn.t20 314.466
R14481 vbn.n230 vbn.t44 314.466
R14482 vbn.n230 vbn.t28 314.466
R14483 vbn.n232 vbn.t34 314.466
R14484 vbn.n232 vbn.t14 314.466
R14485 vbn.n235 vbn.t26 314.466
R14486 vbn.n235 vbn.t8 314.466
R14487 vbn.n237 vbn.t22 314.466
R14488 vbn.n237 vbn.t4 314.466
R14489 vbn.n240 vbn.t2 314.466
R14490 vbn.n240 vbn.t52 314.466
R14491 vbn.n242 vbn.t0 314.466
R14492 vbn.n242 vbn.t48 314.466
R14493 vbn.n245 vbn.t50 314.466
R14494 vbn.n245 vbn.t38 314.466
R14495 vbn.n247 vbn.t46 314.466
R14496 vbn.n247 vbn.t32 314.466
R14497 vbn.n114 vbn.t42 314.466
R14498 vbn.n114 vbn.t24 314.466
R14499 vbn.n222 vbn.t36 314.466
R14500 vbn.n222 vbn.t18 314.466
R14501 vbn.n220 vbn.t30 314.466
R14502 vbn.n220 vbn.t12 314.466
R14503 vbn.n99 vbn.t16 314.466
R14504 vbn.n99 vbn.t58 314.466
R14505 vbn.n255 vbn.t10 314.466
R14506 vbn.n255 vbn.t56 314.466
R14507 vbn.n257 vbn.t6 314.466
R14508 vbn.n257 vbn.t54 314.466
R14509 vbn.n95 vbn.t289 314.466
R14510 vbn.n95 vbn.t269 314.466
R14511 vbn.n93 vbn.t261 314.466
R14512 vbn.n93 vbn.t271 314.466
R14513 vbn.n91 vbn.t264 314.466
R14514 vbn.n91 vbn.t274 314.466
R14515 vbn.n89 vbn.t266 314.466
R14516 vbn.n89 vbn.t276 314.466
R14517 vbn.n87 vbn.t268 314.466
R14518 vbn.n87 vbn.t278 314.466
R14519 vbn.n85 vbn.t279 314.466
R14520 vbn.n85 vbn.t285 314.466
R14521 vbn.n83 vbn.t284 314.466
R14522 vbn.n83 vbn.t260 314.466
R14523 vbn.n81 vbn.t286 314.466
R14524 vbn.n81 vbn.t262 314.466
R14525 vbn.n79 vbn.t287 314.466
R14526 vbn.n79 vbn.t265 314.466
R14527 vbn.n77 vbn.t288 314.466
R14528 vbn.n77 vbn.t267 314.466
R14529 vbn.n75 vbn.t263 314.466
R14530 vbn.n75 vbn.t272 314.466
R14531 vbn.n73 vbn.t270 314.466
R14532 vbn.n73 vbn.t280 314.466
R14533 vbn.n71 vbn.t273 314.466
R14534 vbn.n71 vbn.t281 314.466
R14535 vbn.n69 vbn.t275 314.466
R14536 vbn.n69 vbn.t282 314.466
R14537 vbn.n68 vbn.t277 314.466
R14538 vbn.n68 vbn.t283 314.466
R14539 vbn.n14 vbn.n130 75.3571
R14540 vbn.n26 vbn.n155 75.3571
R14541 vbn.n38 vbn.n180 75.3571
R14542 vbn.n50 vbn.n205 75.3571
R14543 vbn.n64 vbn.n119 75.3477
R14544 vbn.n65 vbn.n144 75.3477
R14545 vbn.n66 vbn.n169 75.3477
R14546 vbn.n67 vbn.n194 75.3477
R14547 vbn.n64 vbn.n121 75.3376
R14548 vbn.n7 vbn.n120 75.3376
R14549 vbn.n7 vbn.n123 75.3376
R14550 vbn.n7 vbn.n122 75.3376
R14551 vbn.n23 vbn.n125 75.3376
R14552 vbn.n23 vbn.n124 75.3376
R14553 vbn.n24 vbn.n127 75.3376
R14554 vbn.n24 vbn.n126 75.3376
R14555 vbn.n22 vbn.n129 75.3376
R14556 vbn.n22 vbn.n128 75.3376
R14557 vbn.n20 vbn.n143 75.3376
R14558 vbn.n20 vbn.n142 75.3376
R14559 vbn.n19 vbn.n141 75.3376
R14560 vbn.n19 vbn.n140 75.3376
R14561 vbn.n18 vbn.n139 75.3376
R14562 vbn.n18 vbn.n138 75.3376
R14563 vbn.n17 vbn.n137 75.3376
R14564 vbn.n17 vbn.n136 75.3376
R14565 vbn.n16 vbn.n135 75.3376
R14566 vbn.n16 vbn.n134 75.3376
R14567 vbn.n15 vbn.n133 75.3376
R14568 vbn.n15 vbn.n132 75.3376
R14569 vbn.n14 vbn.n131 75.3376
R14570 vbn.n65 vbn.n146 75.3376
R14571 vbn.n9 vbn.n145 75.3376
R14572 vbn.n9 vbn.n148 75.3376
R14573 vbn.n9 vbn.n147 75.3376
R14574 vbn.n35 vbn.n150 75.3376
R14575 vbn.n35 vbn.n149 75.3376
R14576 vbn.n36 vbn.n152 75.3376
R14577 vbn.n36 vbn.n151 75.3376
R14578 vbn.n34 vbn.n154 75.3376
R14579 vbn.n34 vbn.n153 75.3376
R14580 vbn.n32 vbn.n168 75.3376
R14581 vbn.n32 vbn.n167 75.3376
R14582 vbn.n31 vbn.n166 75.3376
R14583 vbn.n31 vbn.n165 75.3376
R14584 vbn.n30 vbn.n164 75.3376
R14585 vbn.n30 vbn.n163 75.3376
R14586 vbn.n29 vbn.n162 75.3376
R14587 vbn.n29 vbn.n161 75.3376
R14588 vbn.n28 vbn.n160 75.3376
R14589 vbn.n28 vbn.n159 75.3376
R14590 vbn.n27 vbn.n158 75.3376
R14591 vbn.n27 vbn.n157 75.3376
R14592 vbn.n26 vbn.n156 75.3376
R14593 vbn.n66 vbn.n171 75.3376
R14594 vbn.n11 vbn.n170 75.3376
R14595 vbn.n11 vbn.n173 75.3376
R14596 vbn.n11 vbn.n172 75.3376
R14597 vbn.n47 vbn.n175 75.3376
R14598 vbn.n47 vbn.n174 75.3376
R14599 vbn.n48 vbn.n177 75.3376
R14600 vbn.n48 vbn.n176 75.3376
R14601 vbn.n46 vbn.n179 75.3376
R14602 vbn.n46 vbn.n178 75.3376
R14603 vbn.n44 vbn.n193 75.3376
R14604 vbn.n44 vbn.n192 75.3376
R14605 vbn.n43 vbn.n191 75.3376
R14606 vbn.n43 vbn.n190 75.3376
R14607 vbn.n42 vbn.n189 75.3376
R14608 vbn.n42 vbn.n188 75.3376
R14609 vbn.n41 vbn.n187 75.3376
R14610 vbn.n41 vbn.n186 75.3376
R14611 vbn.n40 vbn.n185 75.3376
R14612 vbn.n40 vbn.n184 75.3376
R14613 vbn.n39 vbn.n183 75.3376
R14614 vbn.n39 vbn.n182 75.3376
R14615 vbn.n38 vbn.n181 75.3376
R14616 vbn.n67 vbn.n196 75.3376
R14617 vbn.n13 vbn.n195 75.3376
R14618 vbn.n13 vbn.n198 75.3376
R14619 vbn.n13 vbn.n197 75.3376
R14620 vbn.n59 vbn.n200 75.3376
R14621 vbn.n59 vbn.n199 75.3376
R14622 vbn.n60 vbn.n202 75.3376
R14623 vbn.n60 vbn.n201 75.3376
R14624 vbn.n58 vbn.n204 75.3376
R14625 vbn.n58 vbn.n203 75.3376
R14626 vbn.n56 vbn.n218 75.3376
R14627 vbn.n56 vbn.n217 75.3376
R14628 vbn.n55 vbn.n216 75.3376
R14629 vbn.n55 vbn.n215 75.3376
R14630 vbn.n54 vbn.n214 75.3376
R14631 vbn.n54 vbn.n213 75.3376
R14632 vbn.n53 vbn.n212 75.3376
R14633 vbn.n53 vbn.n211 75.3376
R14634 vbn.n52 vbn.n210 75.3376
R14635 vbn.n52 vbn.n209 75.3376
R14636 vbn.n51 vbn.n208 75.3376
R14637 vbn.n51 vbn.n207 75.3376
R14638 vbn.n50 vbn.n206 75.3376
R14639 vbn.n70 vbn.n68 67.183
R14640 vbn.n229 vbn.n228 67.1406
R14641 vbn.n231 vbn.n230 67.0982
R14642 vbn.n233 vbn.n232 67.0982
R14643 vbn.n236 vbn.n235 67.0982
R14644 vbn.n238 vbn.n237 67.0982
R14645 vbn.n241 vbn.n240 67.0982
R14646 vbn.n243 vbn.n242 67.0982
R14647 vbn.n246 vbn.n245 67.0982
R14648 vbn.n248 vbn.n247 67.0982
R14649 vbn.n115 vbn.n114 67.0982
R14650 vbn.n223 vbn.n222 67.0982
R14651 vbn.n221 vbn.n220 67.0982
R14652 vbn.n100 vbn.n99 67.0982
R14653 vbn.n256 vbn.n255 67.0982
R14654 vbn.n258 vbn.n257 67.0982
R14655 vbn.n96 vbn.n95 67.0982
R14656 vbn.n94 vbn.n93 67.0982
R14657 vbn.n92 vbn.n91 67.0982
R14658 vbn.n90 vbn.n89 67.0982
R14659 vbn.n88 vbn.n87 67.0982
R14660 vbn.n86 vbn.n85 67.0982
R14661 vbn.n84 vbn.n83 67.0982
R14662 vbn.n82 vbn.n81 67.0982
R14663 vbn.n80 vbn.n79 67.0982
R14664 vbn.n78 vbn.n77 67.0982
R14665 vbn.n76 vbn.n75 67.0982
R14666 vbn.n74 vbn.n73 67.0982
R14667 vbn.n72 vbn.n71 67.0982
R14668 vbn.n70 vbn.n69 67.0982
R14669 vbn.n102 vbn.t55 30.6505
R14670 vbn.n101 vbn.t7 30.6505
R14671 vbn.n110 vbn.n109 24.8505
R14672 vbn.n227 vbn.n226 24.8505
R14673 vbn.n104 vbn.n103 24.8505
R14674 vbn.n251 vbn.n250 24.8505
R14675 vbn.n106 vbn.n105 24.8505
R14676 vbn.n112 vbn.n111 24.8505
R14677 vbn.n108 vbn.n107 24.8505
R14678 vbn.n0 vbn.n118 24.8505
R14679 vbn.n4 vbn.n117 24.8505
R14680 vbn.n1 vbn.n116 24.8505
R14681 vbn.n3 vbn.n113 24.8505
R14682 vbn.n225 vbn.n219 24.8505
R14683 vbn.n2 vbn.n98 24.8505
R14684 vbn.n253 vbn.n252 24.8505
R14685 vbn.n119 vbn.t120 9.52217
R14686 vbn.n119 vbn.t213 9.52217
R14687 vbn.n121 vbn.t92 9.52217
R14688 vbn.n121 vbn.t200 9.52217
R14689 vbn.n120 vbn.t257 9.52217
R14690 vbn.n120 vbn.t75 9.52217
R14691 vbn.n123 vbn.t123 9.52217
R14692 vbn.n123 vbn.t115 9.52217
R14693 vbn.n122 vbn.t217 9.52217
R14694 vbn.n122 vbn.t133 9.52217
R14695 vbn.n125 vbn.t128 9.52217
R14696 vbn.n125 vbn.t186 9.52217
R14697 vbn.n124 vbn.t111 9.52217
R14698 vbn.n124 vbn.t247 9.52217
R14699 vbn.n127 vbn.t121 9.52217
R14700 vbn.n127 vbn.t114 9.52217
R14701 vbn.n126 vbn.t164 9.52217
R14702 vbn.n126 vbn.t227 9.52217
R14703 vbn.n129 vbn.t214 9.52217
R14704 vbn.n129 vbn.t77 9.52217
R14705 vbn.n128 vbn.t156 9.52217
R14706 vbn.n128 vbn.t245 9.52217
R14707 vbn.n143 vbn.t145 9.52217
R14708 vbn.n143 vbn.t221 9.52217
R14709 vbn.n142 vbn.t127 9.52217
R14710 vbn.n142 vbn.t196 9.52217
R14711 vbn.n141 vbn.t86 9.52217
R14712 vbn.n141 vbn.t242 9.52217
R14713 vbn.n140 vbn.t182 9.52217
R14714 vbn.n140 vbn.t85 9.52217
R14715 vbn.n139 vbn.t144 9.52217
R14716 vbn.n139 vbn.t135 9.52217
R14717 vbn.n138 vbn.t189 9.52217
R14718 vbn.n138 vbn.t185 9.52217
R14719 vbn.n137 vbn.t87 9.52217
R14720 vbn.n137 vbn.t64 9.52217
R14721 vbn.n136 vbn.t94 9.52217
R14722 vbn.n136 vbn.t84 9.52217
R14723 vbn.n135 vbn.t99 9.52217
R14724 vbn.n135 vbn.t232 9.52217
R14725 vbn.n134 vbn.t212 9.52217
R14726 vbn.n134 vbn.t105 9.52217
R14727 vbn.n133 vbn.t234 9.52217
R14728 vbn.n133 vbn.t210 9.52217
R14729 vbn.n132 vbn.t73 9.52217
R14730 vbn.n132 vbn.t91 9.52217
R14731 vbn.n131 vbn.t208 9.52217
R14732 vbn.n131 vbn.t104 9.52217
R14733 vbn.n130 vbn.t249 9.52217
R14734 vbn.n130 vbn.t256 9.52217
R14735 vbn.n144 vbn.t224 9.52217
R14736 vbn.n144 vbn.t103 9.52217
R14737 vbn.n146 vbn.t177 9.52217
R14738 vbn.n146 vbn.t109 9.52217
R14739 vbn.n145 vbn.t226 9.52217
R14740 vbn.n145 vbn.t151 9.52217
R14741 vbn.n148 vbn.t149 9.52217
R14742 vbn.n148 vbn.t241 9.52217
R14743 vbn.n147 vbn.t173 9.52217
R14744 vbn.n147 vbn.t229 9.52217
R14745 vbn.n150 vbn.t66 9.52217
R14746 vbn.n150 vbn.t238 9.52217
R14747 vbn.n149 vbn.t236 9.52217
R14748 vbn.n149 vbn.t130 9.52217
R14749 vbn.n152 vbn.t167 9.52217
R14750 vbn.n152 vbn.t170 9.52217
R14751 vbn.n151 vbn.t246 9.52217
R14752 vbn.n151 vbn.t199 9.52217
R14753 vbn.n154 vbn.t134 9.52217
R14754 vbn.n154 vbn.t166 9.52217
R14755 vbn.n153 vbn.t143 9.52217
R14756 vbn.n153 vbn.t155 9.52217
R14757 vbn.n168 vbn.t233 9.52217
R14758 vbn.n168 vbn.t204 9.52217
R14759 vbn.n167 vbn.t219 9.52217
R14760 vbn.n167 vbn.t98 9.52217
R14761 vbn.n166 vbn.t183 9.52217
R14762 vbn.n166 vbn.t184 9.52217
R14763 vbn.n165 vbn.t89 9.52217
R14764 vbn.n165 vbn.t255 9.52217
R14765 vbn.n164 vbn.t139 9.52217
R14766 vbn.n164 vbn.t259 9.52217
R14767 vbn.n163 vbn.t159 9.52217
R14768 vbn.n163 vbn.t207 9.52217
R14769 vbn.n162 vbn.t116 9.52217
R14770 vbn.n162 vbn.t71 9.52217
R14771 vbn.n161 vbn.t231 9.52217
R14772 vbn.n161 vbn.t218 9.52217
R14773 vbn.n160 vbn.t162 9.52217
R14774 vbn.n160 vbn.t63 9.52217
R14775 vbn.n159 vbn.t174 9.52217
R14776 vbn.n159 vbn.t223 9.52217
R14777 vbn.n158 vbn.t131 9.52217
R14778 vbn.n158 vbn.t154 9.52217
R14779 vbn.n157 vbn.t258 9.52217
R14780 vbn.n157 vbn.t78 9.52217
R14781 vbn.n156 vbn.t206 9.52217
R14782 vbn.n156 vbn.t122 9.52217
R14783 vbn.n155 vbn.t74 9.52217
R14784 vbn.n155 vbn.t132 9.52217
R14785 vbn.n169 vbn.t136 9.52217
R14786 vbn.n169 vbn.t230 9.52217
R14787 vbn.n171 vbn.t220 9.52217
R14788 vbn.n171 vbn.t202 9.52217
R14789 vbn.n170 vbn.t150 9.52217
R14790 vbn.n170 vbn.t117 9.52217
R14791 vbn.n173 vbn.t209 9.52217
R14792 vbn.n173 vbn.t169 9.52217
R14793 vbn.n172 vbn.t168 9.52217
R14794 vbn.n172 vbn.t197 9.52217
R14795 vbn.n175 vbn.t175 9.52217
R14796 vbn.n175 vbn.t93 9.52217
R14797 vbn.n174 vbn.t228 9.52217
R14798 vbn.n174 vbn.t180 9.52217
R14799 vbn.n177 vbn.t100 9.52217
R14800 vbn.n177 vbn.t152 9.52217
R14801 vbn.n176 vbn.t76 9.52217
R14802 vbn.n176 vbn.t72 9.52217
R14803 vbn.n179 vbn.t124 9.52217
R14804 vbn.n179 vbn.t201 9.52217
R14805 vbn.n178 vbn.t193 9.52217
R14806 vbn.n178 vbn.t110 9.52217
R14807 vbn.n193 vbn.t248 9.52217
R14808 vbn.n193 vbn.t88 9.52217
R14809 vbn.n192 vbn.t138 9.52217
R14810 vbn.n192 vbn.t190 9.52217
R14811 vbn.n191 vbn.t163 9.52217
R14812 vbn.n191 vbn.t178 9.52217
R14813 vbn.n190 vbn.t216 9.52217
R14814 vbn.n190 vbn.t67 9.52217
R14815 vbn.n189 vbn.t108 9.52217
R14816 vbn.n189 vbn.t251 9.52217
R14817 vbn.n188 vbn.t203 9.52217
R14818 vbn.n188 vbn.t129 9.52217
R14819 vbn.n187 vbn.t69 9.52217
R14820 vbn.n187 vbn.t79 9.52217
R14821 vbn.n186 vbn.t243 9.52217
R14822 vbn.n186 vbn.t82 9.52217
R14823 vbn.n185 vbn.t65 9.52217
R14824 vbn.n185 vbn.t253 9.52217
R14825 vbn.n184 vbn.t106 9.52217
R14826 vbn.n184 vbn.t61 9.52217
R14827 vbn.n183 vbn.t161 9.52217
R14828 vbn.n183 vbn.t81 9.52217
R14829 vbn.n182 vbn.t235 9.52217
R14830 vbn.n182 vbn.t237 9.52217
R14831 vbn.n181 vbn.t187 9.52217
R14832 vbn.n181 vbn.t160 9.52217
R14833 vbn.n180 vbn.t141 9.52217
R14834 vbn.n180 vbn.t147 9.52217
R14835 vbn.n194 vbn.t137 9.52217
R14836 vbn.n194 vbn.t195 9.52217
R14837 vbn.n196 vbn.t165 9.52217
R14838 vbn.n196 vbn.t240 9.52217
R14839 vbn.n195 vbn.t113 9.52217
R14840 vbn.n195 vbn.t118 9.52217
R14841 vbn.n198 vbn.t211 9.52217
R14842 vbn.n198 vbn.t171 9.52217
R14843 vbn.n197 vbn.t225 9.52217
R14844 vbn.n197 vbn.t198 9.52217
R14845 vbn.n200 vbn.t176 9.52217
R14846 vbn.n200 vbn.t96 9.52217
R14847 vbn.n199 vbn.t179 9.52217
R14848 vbn.n199 vbn.t181 9.52217
R14849 vbn.n202 vbn.t146 9.52217
R14850 vbn.n202 vbn.t153 9.52217
R14851 vbn.n201 vbn.t70 9.52217
R14852 vbn.n201 vbn.t97 9.52217
R14853 vbn.n204 vbn.t126 9.52217
R14854 vbn.n204 vbn.t239 9.52217
R14855 vbn.n203 vbn.t194 9.52217
R14856 vbn.n203 vbn.t112 9.52217
R14857 vbn.n218 vbn.t250 9.52217
R14858 vbn.n218 vbn.t158 9.52217
R14859 vbn.n217 vbn.t140 9.52217
R14860 vbn.n217 vbn.t191 9.52217
R14861 vbn.n216 vbn.t102 9.52217
R14862 vbn.n216 vbn.t95 9.52217
R14863 vbn.n215 vbn.t119 9.52217
R14864 vbn.n215 vbn.t68 9.52217
R14865 vbn.n214 vbn.t222 9.52217
R14866 vbn.n214 vbn.t252 9.52217
R14867 vbn.n213 vbn.t205 9.52217
R14868 vbn.n213 vbn.t107 9.52217
R14869 vbn.n212 vbn.t125 9.52217
R14870 vbn.n212 vbn.t80 9.52217
R14871 vbn.n211 vbn.t244 9.52217
R14872 vbn.n211 vbn.t83 9.52217
R14873 vbn.n210 vbn.t254 9.52217
R14874 vbn.n210 vbn.t215 9.52217
R14875 vbn.n209 vbn.t60 9.52217
R14876 vbn.n209 vbn.t62 9.52217
R14877 vbn.n208 vbn.t101 9.52217
R14878 vbn.n208 vbn.t90 9.52217
R14879 vbn.n207 vbn.t157 9.52217
R14880 vbn.n207 vbn.t172 9.52217
R14881 vbn.n206 vbn.t188 9.52217
R14882 vbn.n206 vbn.t192 9.52217
R14883 vbn.n205 vbn.t142 9.52217
R14884 vbn.n205 vbn.t148 9.52217
R14885 vbn.n109 vbn.t29 5.8005
R14886 vbn.n109 vbn.t21 5.8005
R14887 vbn.n226 vbn.t45 5.8005
R14888 vbn.n226 vbn.t41 5.8005
R14889 vbn.n103 vbn.t13 5.8005
R14890 vbn.n103 vbn.t19 5.8005
R14891 vbn.n250 vbn.t25 5.8005
R14892 vbn.n250 vbn.t33 5.8005
R14893 vbn.n105 vbn.t39 5.8005
R14894 vbn.n105 vbn.t49 5.8005
R14895 vbn.n111 vbn.t53 5.8005
R14896 vbn.n111 vbn.t5 5.8005
R14897 vbn.n107 vbn.t9 5.8005
R14898 vbn.n107 vbn.t15 5.8005
R14899 vbn.n118 vbn.t27 5.8005
R14900 vbn.n118 vbn.t35 5.8005
R14901 vbn.n117 vbn.t3 5.8005
R14902 vbn.n117 vbn.t23 5.8005
R14903 vbn.n116 vbn.t51 5.8005
R14904 vbn.n116 vbn.t1 5.8005
R14905 vbn.n113 vbn.t43 5.8005
R14906 vbn.n113 vbn.t47 5.8005
R14907 vbn.n219 vbn.t31 5.8005
R14908 vbn.n219 vbn.t37 5.8005
R14909 vbn.n98 vbn.t11 5.8005
R14910 vbn.n98 vbn.t17 5.8005
R14911 vbn.n252 vbn.t57 5.8005
R14912 vbn.n252 vbn.t59 5.8005
R14913 vbn.n5 vbn.n102 1.07649
R14914 vbn.n5 vbn.n101 1.07649
R14915 vbn.n5 vbn.n104 0.974786
R14916 vbn.n5 vbn.n251 0.974786
R14917 vbn.n5 vbn.n106 0.974786
R14918 vbn.n5 vbn.n112 0.974786
R14919 vbn.n5 vbn.n108 0.974786
R14920 vbn.n5 vbn.n0 0.974786
R14921 vbn.n5 vbn.n4 0.974786
R14922 vbn.n5 vbn.n1 0.974786
R14923 vbn.n5 vbn.n3 0.974786
R14924 vbn.n5 vbn.n225 0.974786
R14925 vbn.n5 vbn.n2 0.974786
R14926 vbn.n227 vbn.n5 0.974786
R14927 vbn.n5 vbn.n110 0.974786
R14928 vbn.n253 vbn.n5 0.974786
R14929 vbn.n224 vbn.n104 0.71925
R14930 vbn.n251 vbn.n249 0.71925
R14931 vbn.n244 vbn.n106 0.71925
R14932 vbn.n239 vbn.n112 0.71925
R14933 vbn.n234 vbn.n108 0.71925
R14934 vbn.n234 vbn.n0 0.71925
R14935 vbn.n239 vbn.n4 0.71925
R14936 vbn.n244 vbn.n1 0.71925
R14937 vbn.n249 vbn.n3 0.71925
R14938 vbn.n225 vbn.n224 0.71925
R14939 vbn.n254 vbn.n2 0.71925
R14940 vbn.n102 vbn.n97 0.71925
R14941 vbn.n101 vbn.n97 0.71925
R14942 vbn.n229 vbn.n227 0.71925
R14943 vbn.n229 vbn.n110 0.71925
R14944 vbn.n254 vbn.n253 0.71925
R14945 vbn.n63 vbn.n57 0.111521
R14946 vbn.n57 vbn.n60 0.0192606
R14947 vbn.n63 vbn.n61 0.111521
R14948 vbn.n61 vbn.n13 0.0192606
R14949 vbn.n63 vbn.n12 0.113704
R14950 vbn.n12 vbn.n67 0.0148932
R14951 vbn.n63 vbn.n45 0.111521
R14952 vbn.n45 vbn.n48 0.0192606
R14953 vbn.n63 vbn.n49 0.111521
R14954 vbn.n49 vbn.n11 0.0192606
R14955 vbn.n63 vbn.n10 0.113704
R14956 vbn.n10 vbn.n66 0.0148932
R14957 vbn.n62 vbn.n33 0.111521
R14958 vbn.n33 vbn.n36 0.0192606
R14959 vbn.n62 vbn.n37 0.111521
R14960 vbn.n37 vbn.n9 0.0192606
R14961 vbn.n62 vbn.n8 0.113704
R14962 vbn.n8 vbn.n65 0.0148932
R14963 vbn.n62 vbn.n21 0.111521
R14964 vbn.n21 vbn.n24 0.0192606
R14965 vbn.n62 vbn.n25 0.111521
R14966 vbn.n25 vbn.n7 0.0192606
R14967 vbn.n62 vbn.n6 0.113704
R14968 vbn.n6 vbn.n64 0.0148932
R14969 vbn.n97 vbn.n96 0.206678
R14970 vbn.n5 vbn.n63 0.18421
R14971 vbn.n72 vbn.n70 0.0852701
R14972 vbn.n74 vbn.n72 0.0852701
R14973 vbn.n76 vbn.n74 0.0852701
R14974 vbn.n78 vbn.n76 0.0852701
R14975 vbn.n80 vbn.n78 0.0852701
R14976 vbn.n82 vbn.n80 0.0852701
R14977 vbn.n84 vbn.n82 0.0852701
R14978 vbn.n86 vbn.n84 0.0852701
R14979 vbn.n88 vbn.n86 0.0852701
R14980 vbn.n90 vbn.n88 0.0852701
R14981 vbn.n92 vbn.n90 0.0852701
R14982 vbn.n94 vbn.n92 0.0852701
R14983 vbn.n96 vbn.n94 0.0852701
R14984 vbn.n258 vbn.n256 0.0852701
R14985 vbn.n221 vbn.n100 0.0852701
R14986 vbn.n223 vbn.n115 0.0852701
R14987 vbn.n248 vbn.n246 0.0852701
R14988 vbn.n243 vbn.n241 0.0852701
R14989 vbn.n238 vbn.n236 0.0852701
R14990 vbn.n233 vbn.n231 0.0852701
R14991 vbn.n63 vbn.n62 0.0483793
R14992 vbn.n256 vbn.n254 0.0428851
R14993 vbn.n254 vbn.n100 0.0428851
R14994 vbn.n224 vbn.n221 0.0428851
R14995 vbn.n224 vbn.n223 0.0428851
R14996 vbn.n249 vbn.n115 0.0428851
R14997 vbn.n249 vbn.n248 0.0428851
R14998 vbn.n246 vbn.n244 0.0428851
R14999 vbn.n244 vbn.n243 0.0428851
R15000 vbn.n241 vbn.n239 0.0428851
R15001 vbn.n239 vbn.n238 0.0428851
R15002 vbn.n236 vbn.n234 0.0428851
R15003 vbn.n234 vbn.n233 0.0428851
R15004 vbn.n231 vbn.n229 0.0428851
R15005 vbn.n258 vbn.n97 0.0428851
R15006 vbn.n59 vbn.n61 0.0192606
R15007 vbn.n60 vbn.n59 0.0400382
R15008 vbn.n58 vbn.n57 0.0192606
R15009 vbn.n58 vbn.n56 0.0400382
R15010 vbn.n47 vbn.n49 0.0192606
R15011 vbn.n48 vbn.n47 0.0400382
R15012 vbn.n46 vbn.n45 0.0192606
R15013 vbn.n46 vbn.n44 0.0400382
R15014 vbn.n35 vbn.n37 0.0192606
R15015 vbn.n36 vbn.n35 0.0400382
R15016 vbn.n34 vbn.n33 0.0192606
R15017 vbn.n34 vbn.n32 0.0400382
R15018 vbn.n23 vbn.n25 0.0192606
R15019 vbn.n24 vbn.n23 0.0400382
R15020 vbn.n22 vbn.n21 0.0192606
R15021 vbn.n22 vbn.n20 0.0400382
R15022 vbn.n56 vbn.n55 0.0394193
R15023 vbn.n55 vbn.n54 0.0394193
R15024 vbn.n54 vbn.n53 0.0394193
R15025 vbn.n53 vbn.n52 0.0394193
R15026 vbn.n52 vbn.n51 0.0394193
R15027 vbn.n51 vbn.n50 0.0394193
R15028 vbn.n44 vbn.n43 0.0394193
R15029 vbn.n43 vbn.n42 0.0394193
R15030 vbn.n42 vbn.n41 0.0394193
R15031 vbn.n41 vbn.n40 0.0394193
R15032 vbn.n40 vbn.n39 0.0394193
R15033 vbn.n39 vbn.n38 0.0394193
R15034 vbn.n32 vbn.n31 0.0394193
R15035 vbn.n31 vbn.n30 0.0394193
R15036 vbn.n30 vbn.n29 0.0394193
R15037 vbn.n29 vbn.n28 0.0394193
R15038 vbn.n28 vbn.n27 0.0394193
R15039 vbn.n27 vbn.n26 0.0394193
R15040 vbn.n20 vbn.n19 0.0394193
R15041 vbn.n19 vbn.n18 0.0394193
R15042 vbn.n18 vbn.n17 0.0394193
R15043 vbn.n17 vbn.n16 0.0394193
R15044 vbn.n16 vbn.n15 0.0394193
R15045 vbn.n15 vbn.n14 0.0394193
R15046 vbn.n13 vbn.n12 0.0349718
R15047 vbn.n11 vbn.n10 0.0349718
R15048 vbn.n9 vbn.n8 0.0349718
R15049 vbn.n7 vbn.n6 0.0349718
R15050 w_4660_n6791.n1763 w_4660_n6791.n110 13874.1
R15051 w_4660_n6791.n2650 w_4660_n6791.n110 13874.1
R15052 w_4660_n6791.n1763 w_4660_n6791.n111 13874.1
R15053 w_4660_n6791.n2650 w_4660_n6791.n111 13874.1
R15054 w_4660_n6791.n452 w_4660_n6791.n238 13874.1
R15055 w_4660_n6791.n238 w_4660_n6791.n112 13874.1
R15056 w_4660_n6791.n452 w_4660_n6791.n239 13874.1
R15057 w_4660_n6791.n239 w_4660_n6791.n112 13874.1
R15058 w_4660_n6791.n1761 w_4660_n6791.n114 13874.1
R15059 w_4660_n6791.n2648 w_4660_n6791.n114 13874.1
R15060 w_4660_n6791.n1761 w_4660_n6791.n115 13874.1
R15061 w_4660_n6791.n2648 w_4660_n6791.n115 13874.1
R15062 w_4660_n6791.n2521 w_4660_n6791.n246 13874.1
R15063 w_4660_n6791.n2521 w_4660_n6791.n113 13874.1
R15064 w_4660_n6791.n246 w_4660_n6791.n244 13874.1
R15065 w_4660_n6791.n244 w_4660_n6791.n113 13874.1
R15066 w_4660_n6791.n1760 w_4660_n6791.n1520 1479.91
R15067 w_4660_n6791.n937 w_4660_n6791.n936 1479.91
R15068 w_4660_n6791.n2520 w_4660_n6791.n247 1479.91
R15069 w_4660_n6791.n1520 w_4660_n6791.n1519 1147.11
R15070 w_4660_n6791.n1421 w_4660_n6791.n937 1147.11
R15071 w_4660_n6791.n2520 w_4660_n6791.n2519 1147.11
R15072 w_4660_n6791.n1760 w_4660_n6791.n1759 356.519
R15073 w_4660_n6791.n1765 w_4660_n6791.n1764 356.519
R15074 w_4660_n6791.n936 w_4660_n6791.n935 353.507
R15075 w_4660_n6791.n1764 w_4660_n6791.n451 353.507
R15076 w_4660_n6791.n2286 w_4660_n6791.n247 332.827
R15077 w_4660_n6791.n2614 w_4660_n6791.t434 85.6582
R15078 w_4660_n6791.n427 w_4660_n6791.t159 85.6582
R15079 w_4660_n6791.n759 w_4660_n6791.t447 85.6582
R15080 w_4660_n6791.n428 w_4660_n6791.t463 85.6582
R15081 w_4660_n6791.n1190 w_4660_n6791.t254 85.6558
R15082 w_4660_n6791.n429 w_4660_n6791.t220 85.6558
R15083 w_4660_n6791.n43 w_4660_n6791.t346 85.4034
R15084 w_4660_n6791.n2266 w_4660_n6791.t349 85.4034
R15085 w_4660_n6791.n2459 w_4660_n6791.t425 85.4034
R15086 w_4660_n6791.n2614 w_4660_n6791.t78 85.4034
R15087 w_4660_n6791.n427 w_4660_n6791.t123 85.4034
R15088 w_4660_n6791.n1190 w_4660_n6791.t239 85.4034
R15089 w_4660_n6791.n429 w_4660_n6791.t273 85.4034
R15090 w_4660_n6791.n2277 w_4660_n6791.t136 85.4034
R15091 w_4660_n6791.n759 w_4660_n6791.t257 85.401
R15092 w_4660_n6791.n428 w_4660_n6791.t221 85.401
R15093 w_4660_n6791.n35 w_4660_n6791.t468 85.3454
R15094 w_4660_n6791.n1959 w_4660_n6791.t460 85.3454
R15095 w_4660_n6791.n2613 w_4660_n6791.n148 76.1366
R15096 w_4660_n6791.n152 w_4660_n6791.n150 76.1366
R15097 w_4660_n6791.n1662 w_4660_n6791.n1660 76.1366
R15098 w_4660_n6791.n1663 w_4660_n6791.n1658 76.1366
R15099 w_4660_n6791.n1664 w_4660_n6791.n1656 76.1366
R15100 w_4660_n6791.n1665 w_4660_n6791.n1654 76.1366
R15101 w_4660_n6791.n1666 w_4660_n6791.n1652 76.1366
R15102 w_4660_n6791.n1667 w_4660_n6791.n1650 76.1366
R15103 w_4660_n6791.n1668 w_4660_n6791.n1648 76.1366
R15104 w_4660_n6791.n1669 w_4660_n6791.n1646 76.1366
R15105 w_4660_n6791.n1670 w_4660_n6791.n1644 76.1366
R15106 w_4660_n6791.n1671 w_4660_n6791.n1642 76.1366
R15107 w_4660_n6791.n1672 w_4660_n6791.n1607 76.1366
R15108 w_4660_n6791.n1641 w_4660_n6791.n1609 76.1366
R15109 w_4660_n6791.n1640 w_4660_n6791.n1611 76.1366
R15110 w_4660_n6791.n1639 w_4660_n6791.n1613 76.1366
R15111 w_4660_n6791.n1638 w_4660_n6791.n1615 76.1366
R15112 w_4660_n6791.n1637 w_4660_n6791.n1617 76.1366
R15113 w_4660_n6791.n1636 w_4660_n6791.n1619 76.1366
R15114 w_4660_n6791.n1635 w_4660_n6791.n1621 76.1366
R15115 w_4660_n6791.n1634 w_4660_n6791.n1623 76.1366
R15116 w_4660_n6791.n1633 w_4660_n6791.n1625 76.1366
R15117 w_4660_n6791.n1632 w_4660_n6791.n1627 76.1366
R15118 w_4660_n6791.n1631 w_4660_n6791.n1629 76.1366
R15119 w_4660_n6791.n758 w_4660_n6791.n687 76.1366
R15120 w_4660_n6791.n757 w_4660_n6791.n689 76.1366
R15121 w_4660_n6791.n756 w_4660_n6791.n691 76.1366
R15122 w_4660_n6791.n755 w_4660_n6791.n693 76.1366
R15123 w_4660_n6791.n754 w_4660_n6791.n695 76.1366
R15124 w_4660_n6791.n753 w_4660_n6791.n697 76.1366
R15125 w_4660_n6791.n752 w_4660_n6791.n699 76.1366
R15126 w_4660_n6791.n751 w_4660_n6791.n701 76.1366
R15127 w_4660_n6791.n750 w_4660_n6791.n703 76.1366
R15128 w_4660_n6791.n749 w_4660_n6791.n705 76.1366
R15129 w_4660_n6791.n748 w_4660_n6791.n707 76.1366
R15130 w_4660_n6791.n747 w_4660_n6791.n709 76.1366
R15131 w_4660_n6791.n746 w_4660_n6791.n711 76.1366
R15132 w_4660_n6791.n745 w_4660_n6791.n713 76.1366
R15133 w_4660_n6791.n744 w_4660_n6791.n715 76.1366
R15134 w_4660_n6791.n743 w_4660_n6791.n717 76.1366
R15135 w_4660_n6791.n742 w_4660_n6791.n719 76.1366
R15136 w_4660_n6791.n741 w_4660_n6791.n721 76.1366
R15137 w_4660_n6791.n740 w_4660_n6791.n723 76.1366
R15138 w_4660_n6791.n739 w_4660_n6791.n725 76.1366
R15139 w_4660_n6791.n738 w_4660_n6791.n727 76.1366
R15140 w_4660_n6791.n737 w_4660_n6791.n729 76.1366
R15141 w_4660_n6791.n736 w_4660_n6791.n731 76.1366
R15142 w_4660_n6791.n735 w_4660_n6791.n733 76.1366
R15143 w_4660_n6791.n1191 w_4660_n6791.n1188 76.1342
R15144 w_4660_n6791.n1192 w_4660_n6791.n1186 76.1342
R15145 w_4660_n6791.n1193 w_4660_n6791.n1184 76.1342
R15146 w_4660_n6791.n1194 w_4660_n6791.n1182 76.1342
R15147 w_4660_n6791.n1195 w_4660_n6791.n1180 76.1342
R15148 w_4660_n6791.n1196 w_4660_n6791.n1178 76.1342
R15149 w_4660_n6791.n1197 w_4660_n6791.n1176 76.1342
R15150 w_4660_n6791.n1198 w_4660_n6791.n1174 76.1342
R15151 w_4660_n6791.n1199 w_4660_n6791.n1172 76.1342
R15152 w_4660_n6791.n1200 w_4660_n6791.n1170 76.1342
R15153 w_4660_n6791.n1201 w_4660_n6791.n1168 76.1342
R15154 w_4660_n6791.n1202 w_4660_n6791.n1166 76.1342
R15155 w_4660_n6791.n1203 w_4660_n6791.n1164 76.1342
R15156 w_4660_n6791.n1204 w_4660_n6791.n1162 76.1342
R15157 w_4660_n6791.n1205 w_4660_n6791.n1160 76.1342
R15158 w_4660_n6791.n1206 w_4660_n6791.n1158 76.1342
R15159 w_4660_n6791.n1207 w_4660_n6791.n1156 76.1342
R15160 w_4660_n6791.n1208 w_4660_n6791.n1154 76.1342
R15161 w_4660_n6791.n1209 w_4660_n6791.n1152 76.1342
R15162 w_4660_n6791.n1210 w_4660_n6791.n1150 76.1342
R15163 w_4660_n6791.n1211 w_4660_n6791.n1148 76.1342
R15164 w_4660_n6791.n1212 w_4660_n6791.n1146 76.1342
R15165 w_4660_n6791.n1213 w_4660_n6791.n1144 76.1342
R15166 w_4660_n6791.n1214 w_4660_n6791.n1142 76.1342
R15167 w_4660_n6791.n2697 w_4660_n6791.n45 75.8817
R15168 w_4660_n6791.n2111 w_4660_n6791.n1921 75.8817
R15169 w_4660_n6791.n2103 w_4660_n6791.n1924 75.8817
R15170 w_4660_n6791.n2097 w_4660_n6791.n1927 75.8817
R15171 w_4660_n6791.n2090 w_4660_n6791.n2089 75.8817
R15172 w_4660_n6791.n1931 w_4660_n6791.n1930 75.8817
R15173 w_4660_n6791.n1934 w_4660_n6791.n1933 75.8817
R15174 w_4660_n6791.n37 w_4660_n6791.n1935 75.8817
R15175 w_4660_n6791.n2073 w_4660_n6791.n1937 75.8817
R15176 w_4660_n6791.n2065 w_4660_n6791.n1941 75.8817
R15177 w_4660_n6791.n2059 w_4660_n6791.n1945 75.8817
R15178 w_4660_n6791.n2053 w_4660_n6791.n1949 75.8817
R15179 w_4660_n6791.n2047 w_4660_n6791.n1953 75.8817
R15180 w_4660_n6791.n2041 w_4660_n6791.n1957 75.8817
R15181 w_4660_n6791.n2035 w_4660_n6791.n1960 75.8817
R15182 w_4660_n6791.n2029 w_4660_n6791.n1963 75.8817
R15183 w_4660_n6791.n2020 w_4660_n6791.n2019 75.8817
R15184 w_4660_n6791.n2013 w_4660_n6791.n2012 75.8817
R15185 w_4660_n6791.n1971 w_4660_n6791.n1970 75.8817
R15186 w_4660_n6791.n1975 w_4660_n6791.n1974 75.8817
R15187 w_4660_n6791.n1978 w_4660_n6791.n1977 75.8817
R15188 w_4660_n6791.n1980 w_4660_n6791.n1979 75.8817
R15189 w_4660_n6791.n1982 w_4660_n6791.n1981 75.8817
R15190 w_4660_n6791.n2460 w_4660_n6791.n310 75.8817
R15191 w_4660_n6791.n2458 w_4660_n6791.n311 75.8817
R15192 w_4660_n6791.n313 w_4660_n6791.n312 75.8817
R15193 w_4660_n6791.n2433 w_4660_n6791.n2432 75.8817
R15194 w_4660_n6791.n2434 w_4660_n6791.n331 75.8817
R15195 w_4660_n6791.n2431 w_4660_n6791.n332 75.8817
R15196 w_4660_n6791.n334 w_4660_n6791.n333 75.8817
R15197 w_4660_n6791.n2394 w_4660_n6791.n2393 75.8817
R15198 w_4660_n6791.n2395 w_4660_n6791.n2392 75.8817
R15199 w_4660_n6791.n2396 w_4660_n6791.n357 75.8817
R15200 w_4660_n6791.n2391 w_4660_n6791.n358 75.8817
R15201 w_4660_n6791.n360 w_4660_n6791.n359 75.8817
R15202 w_4660_n6791.n2355 w_4660_n6791.n2354 75.8817
R15203 w_4660_n6791.n2356 w_4660_n6791.n2353 75.8817
R15204 w_4660_n6791.n2357 w_4660_n6791.n382 75.8817
R15205 w_4660_n6791.n2352 w_4660_n6791.n383 75.8817
R15206 w_4660_n6791.n385 w_4660_n6791.n384 75.8817
R15207 w_4660_n6791.n2327 w_4660_n6791.n2326 75.8817
R15208 w_4660_n6791.n2328 w_4660_n6791.n404 75.8817
R15209 w_4660_n6791.n2325 w_4660_n6791.n405 75.8817
R15210 w_4660_n6791.n407 w_4660_n6791.n406 75.8817
R15211 w_4660_n6791.n2300 w_4660_n6791.n2299 75.8817
R15212 w_4660_n6791.n2301 w_4660_n6791.n425 75.8817
R15213 w_4660_n6791.n2298 w_4660_n6791.n426 75.8817
R15214 w_4660_n6791.n2613 w_4660_n6791.n149 75.8817
R15215 w_4660_n6791.n152 w_4660_n6791.n151 75.8817
R15216 w_4660_n6791.n1662 w_4660_n6791.n1661 75.8817
R15217 w_4660_n6791.n1663 w_4660_n6791.n1659 75.8817
R15218 w_4660_n6791.n1664 w_4660_n6791.n1657 75.8817
R15219 w_4660_n6791.n1665 w_4660_n6791.n1655 75.8817
R15220 w_4660_n6791.n1666 w_4660_n6791.n1653 75.8817
R15221 w_4660_n6791.n1667 w_4660_n6791.n1651 75.8817
R15222 w_4660_n6791.n1668 w_4660_n6791.n1649 75.8817
R15223 w_4660_n6791.n1669 w_4660_n6791.n1647 75.8817
R15224 w_4660_n6791.n1670 w_4660_n6791.n1645 75.8817
R15225 w_4660_n6791.n1671 w_4660_n6791.n1643 75.8817
R15226 w_4660_n6791.n1672 w_4660_n6791.n1608 75.8817
R15227 w_4660_n6791.n1641 w_4660_n6791.n1610 75.8817
R15228 w_4660_n6791.n1640 w_4660_n6791.n1612 75.8817
R15229 w_4660_n6791.n1639 w_4660_n6791.n1614 75.8817
R15230 w_4660_n6791.n1638 w_4660_n6791.n1616 75.8817
R15231 w_4660_n6791.n1637 w_4660_n6791.n1618 75.8817
R15232 w_4660_n6791.n1636 w_4660_n6791.n1620 75.8817
R15233 w_4660_n6791.n1635 w_4660_n6791.n1622 75.8817
R15234 w_4660_n6791.n1634 w_4660_n6791.n1624 75.8817
R15235 w_4660_n6791.n1633 w_4660_n6791.n1626 75.8817
R15236 w_4660_n6791.n1632 w_4660_n6791.n1628 75.8817
R15237 w_4660_n6791.n1631 w_4660_n6791.n1630 75.8817
R15238 w_4660_n6791.n1191 w_4660_n6791.n1189 75.8817
R15239 w_4660_n6791.n1192 w_4660_n6791.n1187 75.8817
R15240 w_4660_n6791.n1193 w_4660_n6791.n1185 75.8817
R15241 w_4660_n6791.n1194 w_4660_n6791.n1183 75.8817
R15242 w_4660_n6791.n1195 w_4660_n6791.n1181 75.8817
R15243 w_4660_n6791.n1196 w_4660_n6791.n1179 75.8817
R15244 w_4660_n6791.n1197 w_4660_n6791.n1177 75.8817
R15245 w_4660_n6791.n1198 w_4660_n6791.n1175 75.8817
R15246 w_4660_n6791.n1199 w_4660_n6791.n1173 75.8817
R15247 w_4660_n6791.n1200 w_4660_n6791.n1171 75.8817
R15248 w_4660_n6791.n1201 w_4660_n6791.n1169 75.8817
R15249 w_4660_n6791.n1202 w_4660_n6791.n1167 75.8817
R15250 w_4660_n6791.n1203 w_4660_n6791.n1165 75.8817
R15251 w_4660_n6791.n1204 w_4660_n6791.n1163 75.8817
R15252 w_4660_n6791.n1205 w_4660_n6791.n1161 75.8817
R15253 w_4660_n6791.n1206 w_4660_n6791.n1159 75.8817
R15254 w_4660_n6791.n1207 w_4660_n6791.n1157 75.8817
R15255 w_4660_n6791.n1208 w_4660_n6791.n1155 75.8817
R15256 w_4660_n6791.n1209 w_4660_n6791.n1153 75.8817
R15257 w_4660_n6791.n1210 w_4660_n6791.n1151 75.8817
R15258 w_4660_n6791.n1211 w_4660_n6791.n1149 75.8817
R15259 w_4660_n6791.n1212 w_4660_n6791.n1147 75.8817
R15260 w_4660_n6791.n1213 w_4660_n6791.n1145 75.8817
R15261 w_4660_n6791.n1214 w_4660_n6791.n1143 75.8817
R15262 w_4660_n6791.n2704 w_4660_n6791.n2703 75.8817
R15263 w_4660_n6791.n758 w_4660_n6791.n688 75.8793
R15264 w_4660_n6791.n757 w_4660_n6791.n690 75.8793
R15265 w_4660_n6791.n756 w_4660_n6791.n692 75.8793
R15266 w_4660_n6791.n755 w_4660_n6791.n694 75.8793
R15267 w_4660_n6791.n754 w_4660_n6791.n696 75.8793
R15268 w_4660_n6791.n753 w_4660_n6791.n698 75.8793
R15269 w_4660_n6791.n752 w_4660_n6791.n700 75.8793
R15270 w_4660_n6791.n751 w_4660_n6791.n702 75.8793
R15271 w_4660_n6791.n750 w_4660_n6791.n704 75.8793
R15272 w_4660_n6791.n749 w_4660_n6791.n706 75.8793
R15273 w_4660_n6791.n748 w_4660_n6791.n708 75.8793
R15274 w_4660_n6791.n747 w_4660_n6791.n710 75.8793
R15275 w_4660_n6791.n746 w_4660_n6791.n712 75.8793
R15276 w_4660_n6791.n745 w_4660_n6791.n714 75.8793
R15277 w_4660_n6791.n744 w_4660_n6791.n716 75.8793
R15278 w_4660_n6791.n743 w_4660_n6791.n718 75.8793
R15279 w_4660_n6791.n742 w_4660_n6791.n720 75.8793
R15280 w_4660_n6791.n741 w_4660_n6791.n722 75.8793
R15281 w_4660_n6791.n740 w_4660_n6791.n724 75.8793
R15282 w_4660_n6791.n739 w_4660_n6791.n726 75.8793
R15283 w_4660_n6791.n738 w_4660_n6791.n728 75.8793
R15284 w_4660_n6791.n737 w_4660_n6791.n730 75.8793
R15285 w_4660_n6791.n736 w_4660_n6791.n732 75.8793
R15286 w_4660_n6791.n735 w_4660_n6791.n734 75.8793
R15287 w_4660_n6791.n38 w_4660_n6791.n1986 75.8237
R15288 w_4660_n6791.n0 w_4660_n6791.n1992 75.8237
R15289 w_4660_n6791.n1999 w_4660_n6791.n1998 75.8237
R15290 w_4660_n6791.n1973 w_4660_n6791.n1972 75.8237
R15291 w_4660_n6791.n1969 w_4660_n6791.n1968 75.8237
R15292 w_4660_n6791.n1966 w_4660_n6791.n1965 75.8237
R15293 w_4660_n6791.n2025 w_4660_n6791.n2024 75.8237
R15294 w_4660_n6791.n1956 w_4660_n6791.n1955 75.8237
R15295 w_4660_n6791.n1952 w_4660_n6791.n1951 75.8237
R15296 w_4660_n6791.n1948 w_4660_n6791.n1947 75.8237
R15297 w_4660_n6791.n1944 w_4660_n6791.n1943 75.8237
R15298 w_4660_n6791.n1940 w_4660_n6791.n1939 75.8237
R15299 w_4660_n6791.n2070 w_4660_n6791.n2069 75.8237
R15300 w_4660_n6791.n4 w_4660_n6791.n2077 75.8237
R15301 w_4660_n6791.n2471 w_4660_n6791.n2470 57.4714
R15302 w_4660_n6791.n450 w_4660_n6791.n447 36.4064
R15303 w_4660_n6791.n71 w_4660_n6791.n69 36.4064
R15304 w_4660_n6791.n301 w_4660_n6791.n299 36.4064
R15305 w_4660_n6791.n75 w_4660_n6791.n69 36.4064
R15306 w_4660_n6791.n448 w_4660_n6791.n447 36.4064
R15307 w_4660_n6791.n1222 w_4660_n6791.n1216 36.4064
R15308 w_4660_n6791.n1220 w_4660_n6791.n1216 36.4064
R15309 w_4660_n6791.n934 w_4660_n6791.n506 36.4064
R15310 w_4660_n6791.n934 w_4660_n6791.n933 36.4064
R15311 w_4660_n6791.n2288 w_4660_n6791.n2287 36.4064
R15312 w_4660_n6791.n2469 w_4660_n6791.n2468 36.4064
R15313 w_4660_n6791.n1758 w_4660_n6791.n1522 36.4064
R15314 w_4660_n6791.n1758 w_4660_n6791.n1757 36.4064
R15315 w_4660_n6791.n73 w_4660_n6791.n72 34.5085
R15316 w_4660_n6791.n2475 w_4660_n6791.n2474 34.5085
R15317 w_4660_n6791.n1475 w_4660_n6791.n1474 34.3446
R15318 w_4660_n6791.n1476 w_4660_n6791.n1475 34.3446
R15319 w_4660_n6791.n1472 w_4660_n6791.n1471 34.3446
R15320 w_4660_n6791.n1471 w_4660_n6791.n1470 34.3446
R15321 w_4660_n6791.n1418 w_4660_n6791.n1417 34.032
R15322 w_4660_n6791.n253 w_4660_n6791.n252 34.032
R15323 w_4660_n6791.n944 w_4660_n6791.n941 34.032
R15324 w_4660_n6791.n257 w_4660_n6791.n256 34.032
R15325 w_4660_n6791.n1417 w_4660_n6791.n1416 34.0311
R15326 w_4660_n6791.n253 w_4660_n6791.n138 34.0311
R15327 w_4660_n6791.n945 w_4660_n6791.n944 34.0311
R15328 w_4660_n6791.n256 w_4660_n6791.n255 34.0311
R15329 w_4660_n6791.n2286 w_4660_n6791.n2283 33.0027
R15330 w_4660_n6791.n991 w_4660_n6791.n990 30.4946
R15331 w_4660_n6791.n1410 w_4660_n6791.n938 30.4946
R15332 w_4660_n6791.n766 w_4660_n6791.n684 30.4946
R15333 w_4660_n6791.n770 w_4660_n6791.n761 30.4946
R15334 w_4660_n6791.n83 w_4660_n6791.n82 27.4829
R15335 w_4660_n6791.n2620 w_4660_n6791.n144 27.4829
R15336 w_4660_n6791.n2618 w_4660_n6791.n2617 27.4829
R15337 w_4660_n6791.n1759 w_4660_n6791.n1521 27.1064
R15338 w_4660_n6791.n1754 w_4660_n6791.n1521 27.1064
R15339 w_4660_n6791.n1754 w_4660_n6791.n1753 27.1064
R15340 w_4660_n6791.n1753 w_4660_n6791.n1752 27.1064
R15341 w_4660_n6791.n1752 w_4660_n6791.n1527 27.1064
R15342 w_4660_n6791.n1746 w_4660_n6791.n1527 27.1064
R15343 w_4660_n6791.n1746 w_4660_n6791.n1745 27.1064
R15344 w_4660_n6791.n1745 w_4660_n6791.n1744 27.1064
R15345 w_4660_n6791.n1744 w_4660_n6791.n1535 27.1064
R15346 w_4660_n6791.n1738 w_4660_n6791.n1535 27.1064
R15347 w_4660_n6791.n1738 w_4660_n6791.n1737 27.1064
R15348 w_4660_n6791.n1737 w_4660_n6791.n1543 27.1064
R15349 w_4660_n6791.n1552 w_4660_n6791.n1543 27.1064
R15350 w_4660_n6791.n1730 w_4660_n6791.n1552 27.1064
R15351 w_4660_n6791.n1730 w_4660_n6791.n1729 27.1064
R15352 w_4660_n6791.n1729 w_4660_n6791.n1728 27.1064
R15353 w_4660_n6791.n1728 w_4660_n6791.n1553 27.1064
R15354 w_4660_n6791.n1722 w_4660_n6791.n1553 27.1064
R15355 w_4660_n6791.n1722 w_4660_n6791.n1721 27.1064
R15356 w_4660_n6791.n1721 w_4660_n6791.n1720 27.1064
R15357 w_4660_n6791.n1720 w_4660_n6791.n1561 27.1064
R15358 w_4660_n6791.n1714 w_4660_n6791.n1561 27.1064
R15359 w_4660_n6791.n1714 w_4660_n6791.n1713 27.1064
R15360 w_4660_n6791.n1713 w_4660_n6791.n1712 27.1064
R15361 w_4660_n6791.n1712 w_4660_n6791.n1570 27.1064
R15362 w_4660_n6791.n1706 w_4660_n6791.n1570 27.1064
R15363 w_4660_n6791.n1706 w_4660_n6791.n1705 27.1064
R15364 w_4660_n6791.n1705 w_4660_n6791.n1580 27.1064
R15365 w_4660_n6791.n1587 w_4660_n6791.n1580 27.1064
R15366 w_4660_n6791.n1699 w_4660_n6791.n1587 27.1064
R15367 w_4660_n6791.n1699 w_4660_n6791.n1698 27.1064
R15368 w_4660_n6791.n1698 w_4660_n6791.n1697 27.1064
R15369 w_4660_n6791.n1697 w_4660_n6791.n1588 27.1064
R15370 w_4660_n6791.n1691 w_4660_n6791.n1588 27.1064
R15371 w_4660_n6791.n1691 w_4660_n6791.n1690 27.1064
R15372 w_4660_n6791.n1690 w_4660_n6791.n1689 27.1064
R15373 w_4660_n6791.n1689 w_4660_n6791.n1597 27.1064
R15374 w_4660_n6791.n1683 w_4660_n6791.n1597 27.1064
R15375 w_4660_n6791.n1683 w_4660_n6791.n1682 27.1064
R15376 w_4660_n6791.n1682 w_4660_n6791.n1681 27.1064
R15377 w_4660_n6791.n1681 w_4660_n6791.n1606 27.1064
R15378 w_4660_n6791.n2527 w_4660_n6791.n232 27.1064
R15379 w_4660_n6791.n2528 w_4660_n6791.n2527 27.1064
R15380 w_4660_n6791.n2528 w_4660_n6791.n226 27.1064
R15381 w_4660_n6791.n2534 w_4660_n6791.n226 27.1064
R15382 w_4660_n6791.n2535 w_4660_n6791.n2534 27.1064
R15383 w_4660_n6791.n2535 w_4660_n6791.n220 27.1064
R15384 w_4660_n6791.n2541 w_4660_n6791.n220 27.1064
R15385 w_4660_n6791.n2542 w_4660_n6791.n2541 27.1064
R15386 w_4660_n6791.n2542 w_4660_n6791.n211 27.1064
R15387 w_4660_n6791.n2548 w_4660_n6791.n211 27.1064
R15388 w_4660_n6791.n2549 w_4660_n6791.n2548 27.1064
R15389 w_4660_n6791.n2550 w_4660_n6791.n2549 27.1064
R15390 w_4660_n6791.n2550 w_4660_n6791.n205 27.1064
R15391 w_4660_n6791.n2556 w_4660_n6791.n205 27.1064
R15392 w_4660_n6791.n2557 w_4660_n6791.n2556 27.1064
R15393 w_4660_n6791.n2557 w_4660_n6791.n199 27.1064
R15394 w_4660_n6791.n2563 w_4660_n6791.n199 27.1064
R15395 w_4660_n6791.n2564 w_4660_n6791.n2563 27.1064
R15396 w_4660_n6791.n2564 w_4660_n6791.n190 27.1064
R15397 w_4660_n6791.n2570 w_4660_n6791.n190 27.1064
R15398 w_4660_n6791.n2571 w_4660_n6791.n2570 27.1064
R15399 w_4660_n6791.n2572 w_4660_n6791.n2571 27.1064
R15400 w_4660_n6791.n2572 w_4660_n6791.n184 27.1064
R15401 w_4660_n6791.n2577 w_4660_n6791.n184 27.1064
R15402 w_4660_n6791.n2578 w_4660_n6791.n2577 27.1064
R15403 w_4660_n6791.n2578 w_4660_n6791.n180 27.1064
R15404 w_4660_n6791.n2584 w_4660_n6791.n180 27.1064
R15405 w_4660_n6791.n2585 w_4660_n6791.n2584 27.1064
R15406 w_4660_n6791.n2585 w_4660_n6791.n174 27.1064
R15407 w_4660_n6791.n2591 w_4660_n6791.n174 27.1064
R15408 w_4660_n6791.n2592 w_4660_n6791.n2591 27.1064
R15409 w_4660_n6791.n2592 w_4660_n6791.n168 27.1064
R15410 w_4660_n6791.n2598 w_4660_n6791.n168 27.1064
R15411 w_4660_n6791.n2599 w_4660_n6791.n2598 27.1064
R15412 w_4660_n6791.n2599 w_4660_n6791.n160 27.1064
R15413 w_4660_n6791.n2606 w_4660_n6791.n160 27.1064
R15414 w_4660_n6791.n2607 w_4660_n6791.n2606 27.1064
R15415 w_4660_n6791.n2610 w_4660_n6791.n2607 27.1064
R15416 w_4660_n6791.n2610 w_4660_n6791.n2609 27.1064
R15417 w_4660_n6791.n2609 w_4660_n6791.n2608 27.1064
R15418 w_4660_n6791.n2608 w_4660_n6791.n142 27.1064
R15419 w_4660_n6791.n935 w_4660_n6791.n504 27.1064
R15420 w_4660_n6791.n508 w_4660_n6791.n504 27.1064
R15421 w_4660_n6791.n512 w_4660_n6791.n508 27.1064
R15422 w_4660_n6791.n513 w_4660_n6791.n512 27.1064
R15423 w_4660_n6791.n517 w_4660_n6791.n513 27.1064
R15424 w_4660_n6791.n518 w_4660_n6791.n517 27.1064
R15425 w_4660_n6791.n522 w_4660_n6791.n518 27.1064
R15426 w_4660_n6791.n523 w_4660_n6791.n522 27.1064
R15427 w_4660_n6791.n526 w_4660_n6791.n523 27.1064
R15428 w_4660_n6791.n527 w_4660_n6791.n526 27.1064
R15429 w_4660_n6791.n530 w_4660_n6791.n527 27.1064
R15430 w_4660_n6791.n531 w_4660_n6791.n530 27.1064
R15431 w_4660_n6791.n535 w_4660_n6791.n531 27.1064
R15432 w_4660_n6791.n536 w_4660_n6791.n535 27.1064
R15433 w_4660_n6791.n539 w_4660_n6791.n536 27.1064
R15434 w_4660_n6791.n540 w_4660_n6791.n539 27.1064
R15435 w_4660_n6791.n542 w_4660_n6791.n540 27.1064
R15436 w_4660_n6791.n543 w_4660_n6791.n542 27.1064
R15437 w_4660_n6791.n546 w_4660_n6791.n543 27.1064
R15438 w_4660_n6791.n547 w_4660_n6791.n546 27.1064
R15439 w_4660_n6791.n551 w_4660_n6791.n547 27.1064
R15440 w_4660_n6791.n552 w_4660_n6791.n551 27.1064
R15441 w_4660_n6791.n556 w_4660_n6791.n552 27.1064
R15442 w_4660_n6791.n557 w_4660_n6791.n556 27.1064
R15443 w_4660_n6791.n561 w_4660_n6791.n557 27.1064
R15444 w_4660_n6791.n562 w_4660_n6791.n561 27.1064
R15445 w_4660_n6791.n565 w_4660_n6791.n562 27.1064
R15446 w_4660_n6791.n566 w_4660_n6791.n565 27.1064
R15447 w_4660_n6791.n569 w_4660_n6791.n566 27.1064
R15448 w_4660_n6791.n570 w_4660_n6791.n569 27.1064
R15449 w_4660_n6791.n574 w_4660_n6791.n570 27.1064
R15450 w_4660_n6791.n575 w_4660_n6791.n574 27.1064
R15451 w_4660_n6791.n579 w_4660_n6791.n575 27.1064
R15452 w_4660_n6791.n580 w_4660_n6791.n579 27.1064
R15453 w_4660_n6791.n584 w_4660_n6791.n580 27.1064
R15454 w_4660_n6791.n585 w_4660_n6791.n584 27.1064
R15455 w_4660_n6791.n588 w_4660_n6791.n585 27.1064
R15456 w_4660_n6791.n589 w_4660_n6791.n588 27.1064
R15457 w_4660_n6791.n593 w_4660_n6791.n589 27.1064
R15458 w_4660_n6791.n594 w_4660_n6791.n593 27.1064
R15459 w_4660_n6791.n595 w_4660_n6791.n594 27.1064
R15460 w_4660_n6791.n602 w_4660_n6791.n597 27.1064
R15461 w_4660_n6791.n603 w_4660_n6791.n602 27.1064
R15462 w_4660_n6791.n607 w_4660_n6791.n603 27.1064
R15463 w_4660_n6791.n608 w_4660_n6791.n607 27.1064
R15464 w_4660_n6791.n611 w_4660_n6791.n608 27.1064
R15465 w_4660_n6791.n612 w_4660_n6791.n611 27.1064
R15466 w_4660_n6791.n616 w_4660_n6791.n612 27.1064
R15467 w_4660_n6791.n617 w_4660_n6791.n616 27.1064
R15468 w_4660_n6791.n620 w_4660_n6791.n617 27.1064
R15469 w_4660_n6791.n621 w_4660_n6791.n620 27.1064
R15470 w_4660_n6791.n623 w_4660_n6791.n621 27.1064
R15471 w_4660_n6791.n624 w_4660_n6791.n623 27.1064
R15472 w_4660_n6791.n627 w_4660_n6791.n624 27.1064
R15473 w_4660_n6791.n628 w_4660_n6791.n627 27.1064
R15474 w_4660_n6791.n631 w_4660_n6791.n628 27.1064
R15475 w_4660_n6791.n632 w_4660_n6791.n631 27.1064
R15476 w_4660_n6791.n636 w_4660_n6791.n632 27.1064
R15477 w_4660_n6791.n637 w_4660_n6791.n636 27.1064
R15478 w_4660_n6791.n641 w_4660_n6791.n637 27.1064
R15479 w_4660_n6791.n642 w_4660_n6791.n641 27.1064
R15480 w_4660_n6791.n645 w_4660_n6791.n642 27.1064
R15481 w_4660_n6791.n646 w_4660_n6791.n645 27.1064
R15482 w_4660_n6791.n649 w_4660_n6791.n646 27.1064
R15483 w_4660_n6791.n650 w_4660_n6791.n649 27.1064
R15484 w_4660_n6791.n654 w_4660_n6791.n650 27.1064
R15485 w_4660_n6791.n655 w_4660_n6791.n654 27.1064
R15486 w_4660_n6791.n659 w_4660_n6791.n655 27.1064
R15487 w_4660_n6791.n660 w_4660_n6791.n659 27.1064
R15488 w_4660_n6791.n664 w_4660_n6791.n660 27.1064
R15489 w_4660_n6791.n665 w_4660_n6791.n664 27.1064
R15490 w_4660_n6791.n668 w_4660_n6791.n665 27.1064
R15491 w_4660_n6791.n669 w_4660_n6791.n668 27.1064
R15492 w_4660_n6791.n671 w_4660_n6791.n669 27.1064
R15493 w_4660_n6791.n672 w_4660_n6791.n671 27.1064
R15494 w_4660_n6791.n676 w_4660_n6791.n672 27.1064
R15495 w_4660_n6791.n677 w_4660_n6791.n676 27.1064
R15496 w_4660_n6791.n681 w_4660_n6791.n677 27.1064
R15497 w_4660_n6791.n682 w_4660_n6791.n681 27.1064
R15498 w_4660_n6791.n685 w_4660_n6791.n682 27.1064
R15499 w_4660_n6791.n686 w_4660_n6791.n685 27.1064
R15500 w_4660_n6791.n762 w_4660_n6791.n686 27.1064
R15501 w_4660_n6791.n1770 w_4660_n6791.n450 27.1064
R15502 w_4660_n6791.n2259 w_4660_n6791.n1770 27.1064
R15503 w_4660_n6791.n2259 w_4660_n6791.n2258 27.1064
R15504 w_4660_n6791.n2258 w_4660_n6791.n1771 27.1064
R15505 w_4660_n6791.n1777 w_4660_n6791.n1771 27.1064
R15506 w_4660_n6791.n2252 w_4660_n6791.n1777 27.1064
R15507 w_4660_n6791.n2252 w_4660_n6791.n2251 27.1064
R15508 w_4660_n6791.n2251 w_4660_n6791.n1778 27.1064
R15509 w_4660_n6791.n1787 w_4660_n6791.n1778 27.1064
R15510 w_4660_n6791.n2244 w_4660_n6791.n1787 27.1064
R15511 w_4660_n6791.n2244 w_4660_n6791.n2243 27.1064
R15512 w_4660_n6791.n2243 w_4660_n6791.n2242 27.1064
R15513 w_4660_n6791.n2242 w_4660_n6791.n1788 27.1064
R15514 w_4660_n6791.n2236 w_4660_n6791.n1788 27.1064
R15515 w_4660_n6791.n2236 w_4660_n6791.n2235 27.1064
R15516 w_4660_n6791.n2235 w_4660_n6791.n2234 27.1064
R15517 w_4660_n6791.n2234 w_4660_n6791.n1796 27.1064
R15518 w_4660_n6791.n2228 w_4660_n6791.n1796 27.1064
R15519 w_4660_n6791.n2228 w_4660_n6791.n2227 27.1064
R15520 w_4660_n6791.n2227 w_4660_n6791.n2226 27.1064
R15521 w_4660_n6791.n2226 w_4660_n6791.n1806 27.1064
R15522 w_4660_n6791.n2220 w_4660_n6791.n1806 27.1064
R15523 w_4660_n6791.n2220 w_4660_n6791.n2219 27.1064
R15524 w_4660_n6791.n2219 w_4660_n6791.n1815 27.1064
R15525 w_4660_n6791.n1824 w_4660_n6791.n1815 27.1064
R15526 w_4660_n6791.n2212 w_4660_n6791.n1824 27.1064
R15527 w_4660_n6791.n2212 w_4660_n6791.n2211 27.1064
R15528 w_4660_n6791.n2211 w_4660_n6791.n2210 27.1064
R15529 w_4660_n6791.n2210 w_4660_n6791.n7 27.1064
R15530 w_4660_n6791.n2205 w_4660_n6791.n7 27.1064
R15531 w_4660_n6791.n2205 w_4660_n6791.n2204 27.1064
R15532 w_4660_n6791.n2204 w_4660_n6791.n2203 27.1064
R15533 w_4660_n6791.n2203 w_4660_n6791.n1831 27.1064
R15534 w_4660_n6791.n2197 w_4660_n6791.n1831 27.1064
R15535 w_4660_n6791.n2197 w_4660_n6791.n2196 27.1064
R15536 w_4660_n6791.n2196 w_4660_n6791.n2195 27.1064
R15537 w_4660_n6791.n2195 w_4660_n6791.n1840 27.1064
R15538 w_4660_n6791.n2189 w_4660_n6791.n1840 27.1064
R15539 w_4660_n6791.n2189 w_4660_n6791.n2188 27.1064
R15540 w_4660_n6791.n2188 w_4660_n6791.n1850 27.1064
R15541 w_4660_n6791.n1858 w_4660_n6791.n1850 27.1064
R15542 w_4660_n6791.n2180 w_4660_n6791.n1858 27.1064
R15543 w_4660_n6791.n2180 w_4660_n6791.n2179 27.1064
R15544 w_4660_n6791.n2179 w_4660_n6791.n1859 27.1064
R15545 w_4660_n6791.n1868 w_4660_n6791.n1859 27.1064
R15546 w_4660_n6791.n2172 w_4660_n6791.n1868 27.1064
R15547 w_4660_n6791.n2172 w_4660_n6791.n2171 27.1064
R15548 w_4660_n6791.n2171 w_4660_n6791.n2170 27.1064
R15549 w_4660_n6791.n2170 w_4660_n6791.n1869 27.1064
R15550 w_4660_n6791.n2164 w_4660_n6791.n1869 27.1064
R15551 w_4660_n6791.n2164 w_4660_n6791.n2163 27.1064
R15552 w_4660_n6791.n2163 w_4660_n6791.n2162 27.1064
R15553 w_4660_n6791.n2162 w_4660_n6791.n1877 27.1064
R15554 w_4660_n6791.n2156 w_4660_n6791.n1877 27.1064
R15555 w_4660_n6791.n2156 w_4660_n6791.n2155 27.1064
R15556 w_4660_n6791.n2155 w_4660_n6791.n2154 27.1064
R15557 w_4660_n6791.n2154 w_4660_n6791.n1886 27.1064
R15558 w_4660_n6791.n2148 w_4660_n6791.n1886 27.1064
R15559 w_4660_n6791.n2148 w_4660_n6791.n2147 27.1064
R15560 w_4660_n6791.n2147 w_4660_n6791.n1895 27.1064
R15561 w_4660_n6791.n1904 w_4660_n6791.n1895 27.1064
R15562 w_4660_n6791.n2140 w_4660_n6791.n1904 27.1064
R15563 w_4660_n6791.n2140 w_4660_n6791.n2139 27.1064
R15564 w_4660_n6791.n2139 w_4660_n6791.n2138 27.1064
R15565 w_4660_n6791.n2138 w_4660_n6791.n9 27.1064
R15566 w_4660_n6791.n2132 w_4660_n6791.n9 27.1064
R15567 w_4660_n6791.n2132 w_4660_n6791.n2131 27.1064
R15568 w_4660_n6791.n2131 w_4660_n6791.n2130 27.1064
R15569 w_4660_n6791.n2130 w_4660_n6791.n1911 27.1064
R15570 w_4660_n6791.n2124 w_4660_n6791.n1911 27.1064
R15571 w_4660_n6791.n2124 w_4660_n6791.n2123 27.1064
R15572 w_4660_n6791.n2123 w_4660_n6791.n2122 27.1064
R15573 w_4660_n6791.n2122 w_4660_n6791.n1920 27.1064
R15574 w_4660_n6791.n1920 w_4660_n6791.n1919 27.1064
R15575 w_4660_n6791.n1919 w_4660_n6791.n50 27.1064
R15576 w_4660_n6791.n56 w_4660_n6791.n50 27.1064
R15577 w_4660_n6791.n2690 w_4660_n6791.n56 27.1064
R15578 w_4660_n6791.n2690 w_4660_n6791.n2689 27.1064
R15579 w_4660_n6791.n2689 w_4660_n6791.n2688 27.1064
R15580 w_4660_n6791.n2688 w_4660_n6791.n57 27.1064
R15581 w_4660_n6791.n2682 w_4660_n6791.n57 27.1064
R15582 w_4660_n6791.n2682 w_4660_n6791.n2 32.6532
R15583 w_4660_n6791.n71 w_4660_n6791.n70 27.1064
R15584 w_4660_n6791.n70 w_4660_n6791.n67 27.1064
R15585 w_4660_n6791.n79 w_4660_n6791.n67 27.1064
R15586 w_4660_n6791.n80 w_4660_n6791.n79 27.1064
R15587 w_4660_n6791.n85 w_4660_n6791.n80 27.1064
R15588 w_4660_n6791.n86 w_4660_n6791.n85 27.1064
R15589 w_4660_n6791.n89 w_4660_n6791.n86 27.1064
R15590 w_4660_n6791.n90 w_4660_n6791.n89 27.1064
R15591 w_4660_n6791.n94 w_4660_n6791.n90 27.1064
R15592 w_4660_n6791.n95 w_4660_n6791.n94 27.1064
R15593 w_4660_n6791.n98 w_4660_n6791.n95 27.1064
R15594 w_4660_n6791.n99 w_4660_n6791.n98 27.1064
R15595 w_4660_n6791.n102 w_4660_n6791.n99 27.1064
R15596 w_4660_n6791.n103 w_4660_n6791.n102 27.1064
R15597 w_4660_n6791.n106 w_4660_n6791.n103 27.1064
R15598 w_4660_n6791.n107 w_4660_n6791.n106 27.1064
R15599 w_4660_n6791.n961 w_4660_n6791.n107 27.1064
R15600 w_4660_n6791.n963 w_4660_n6791.n961 27.1064
R15601 w_4660_n6791.n963 w_4660_n6791.n962 27.1064
R15602 w_4660_n6791.n962 w_4660_n6791.n960 27.1064
R15603 w_4660_n6791.n960 w_4660_n6791.n959 27.1064
R15604 w_4660_n6791.n959 w_4660_n6791.n956 27.1064
R15605 w_4660_n6791.n956 w_4660_n6791.n955 27.1064
R15606 w_4660_n6791.n955 w_4660_n6791.n952 27.1064
R15607 w_4660_n6791.n952 w_4660_n6791.n951 27.1064
R15608 w_4660_n6791.n951 w_4660_n6791.n948 27.1064
R15609 w_4660_n6791.n948 w_4660_n6791.n942 27.1064
R15610 w_4660_n6791.n1416 w_4660_n6791.n942 27.1064
R15611 w_4660_n6791.n1418 w_4660_n6791.n500 27.1064
R15612 w_4660_n6791.n1425 w_4660_n6791.n500 27.1064
R15613 w_4660_n6791.n1426 w_4660_n6791.n1425 27.1064
R15614 w_4660_n6791.n1427 w_4660_n6791.n1426 27.1064
R15615 w_4660_n6791.n1427 w_4660_n6791.n492 27.1064
R15616 w_4660_n6791.n1433 w_4660_n6791.n492 27.1064
R15617 w_4660_n6791.n1434 w_4660_n6791.n1433 27.1064
R15618 w_4660_n6791.n1435 w_4660_n6791.n1434 27.1064
R15619 w_4660_n6791.n1435 w_4660_n6791.n484 27.1064
R15620 w_4660_n6791.n1441 w_4660_n6791.n484 27.1064
R15621 w_4660_n6791.n1442 w_4660_n6791.n1441 27.1064
R15622 w_4660_n6791.n1443 w_4660_n6791.n1442 27.1064
R15623 w_4660_n6791.n1443 w_4660_n6791.n476 27.1064
R15624 w_4660_n6791.n1450 w_4660_n6791.n476 27.1064
R15625 w_4660_n6791.n1451 w_4660_n6791.n1450 27.1064
R15626 w_4660_n6791.n1452 w_4660_n6791.n1451 27.1064
R15627 w_4660_n6791.n1452 w_4660_n6791.n468 27.1064
R15628 w_4660_n6791.n1458 w_4660_n6791.n468 27.1064
R15629 w_4660_n6791.n1459 w_4660_n6791.n1458 27.1064
R15630 w_4660_n6791.n1461 w_4660_n6791.n1459 27.1064
R15631 w_4660_n6791.n1461 w_4660_n6791.n1460 27.1064
R15632 w_4660_n6791.n1460 w_4660_n6791.n464 27.1064
R15633 w_4660_n6791.n464 w_4660_n6791.n459 27.1064
R15634 w_4660_n6791.n1474 w_4660_n6791.n459 27.1064
R15635 w_4660_n6791.n1516 w_4660_n6791.n1476 27.1064
R15636 w_4660_n6791.n1516 w_4660_n6791.n1515 27.1064
R15637 w_4660_n6791.n1515 w_4660_n6791.n1514 27.1064
R15638 w_4660_n6791.n1514 w_4660_n6791.n1477 27.1064
R15639 w_4660_n6791.n1508 w_4660_n6791.n1477 27.1064
R15640 w_4660_n6791.n1508 w_4660_n6791.n1507 27.1064
R15641 w_4660_n6791.n1507 w_4660_n6791.n1506 27.1064
R15642 w_4660_n6791.n1506 w_4660_n6791.n1485 27.1064
R15643 w_4660_n6791.n1500 w_4660_n6791.n1485 27.1064
R15644 w_4660_n6791.n1500 w_4660_n6791.n1499 27.1064
R15645 w_4660_n6791.n1499 w_4660_n6791.n1498 27.1064
R15646 w_4660_n6791.n1498 w_4660_n6791.n121 27.1064
R15647 w_4660_n6791.n2644 w_4660_n6791.n121 27.1064
R15648 w_4660_n6791.n2644 w_4660_n6791.n2643 27.1064
R15649 w_4660_n6791.n2643 w_4660_n6791.n2642 27.1064
R15650 w_4660_n6791.n2642 w_4660_n6791.n122 27.1064
R15651 w_4660_n6791.n2636 w_4660_n6791.n122 27.1064
R15652 w_4660_n6791.n2636 w_4660_n6791.n2635 27.1064
R15653 w_4660_n6791.n2635 w_4660_n6791.n2634 27.1064
R15654 w_4660_n6791.n2634 w_4660_n6791.n130 27.1064
R15655 w_4660_n6791.n2628 w_4660_n6791.n130 27.1064
R15656 w_4660_n6791.n2628 w_4660_n6791.n2627 27.1064
R15657 w_4660_n6791.n2627 w_4660_n6791.n2626 27.1064
R15658 w_4660_n6791.n2626 w_4660_n6791.n138 27.1064
R15659 w_4660_n6791.n252 w_4660_n6791.n250 27.1064
R15660 w_4660_n6791.n259 w_4660_n6791.n250 27.1064
R15661 w_4660_n6791.n260 w_4660_n6791.n259 27.1064
R15662 w_4660_n6791.n263 w_4660_n6791.n260 27.1064
R15663 w_4660_n6791.n264 w_4660_n6791.n263 27.1064
R15664 w_4660_n6791.n267 w_4660_n6791.n264 27.1064
R15665 w_4660_n6791.n268 w_4660_n6791.n267 27.1064
R15666 w_4660_n6791.n271 w_4660_n6791.n268 27.1064
R15667 w_4660_n6791.n272 w_4660_n6791.n271 27.1064
R15668 w_4660_n6791.n275 w_4660_n6791.n272 27.1064
R15669 w_4660_n6791.n276 w_4660_n6791.n275 27.1064
R15670 w_4660_n6791.n279 w_4660_n6791.n276 27.1064
R15671 w_4660_n6791.n280 w_4660_n6791.n279 27.1064
R15672 w_4660_n6791.n283 w_4660_n6791.n280 27.1064
R15673 w_4660_n6791.n284 w_4660_n6791.n283 27.1064
R15674 w_4660_n6791.n288 w_4660_n6791.n284 27.1064
R15675 w_4660_n6791.n289 w_4660_n6791.n288 27.1064
R15676 w_4660_n6791.n292 w_4660_n6791.n289 27.1064
R15677 w_4660_n6791.n293 w_4660_n6791.n292 27.1064
R15678 w_4660_n6791.n296 w_4660_n6791.n293 27.1064
R15679 w_4660_n6791.n297 w_4660_n6791.n296 27.1064
R15680 w_4660_n6791.n300 w_4660_n6791.n297 27.1064
R15681 w_4660_n6791.n301 w_4660_n6791.n300 27.1064
R15682 w_4660_n6791.n76 w_4660_n6791.n75 27.1064
R15683 w_4660_n6791.n2681 w_4660_n6791.n76 27.1064
R15684 w_4660_n6791.n2681 w_4660_n6791.n2680 27.1064
R15685 w_4660_n6791.n2680 w_4660_n6791.n2679 27.1064
R15686 w_4660_n6791.n2679 w_4660_n6791.n77 27.1064
R15687 w_4660_n6791.n2672 w_4660_n6791.n77 27.1064
R15688 w_4660_n6791.n2672 w_4660_n6791.n2671 27.1064
R15689 w_4660_n6791.n2671 w_4660_n6791.n2670 27.1064
R15690 w_4660_n6791.n2670 w_4660_n6791.n88 27.1064
R15691 w_4660_n6791.n2664 w_4660_n6791.n88 27.1064
R15692 w_4660_n6791.n2664 w_4660_n6791.n2663 27.1064
R15693 w_4660_n6791.n2663 w_4660_n6791.n2662 27.1064
R15694 w_4660_n6791.n2662 w_4660_n6791.n97 27.1064
R15695 w_4660_n6791.n2656 w_4660_n6791.n97 27.1064
R15696 w_4660_n6791.n2656 w_4660_n6791.n2655 27.1064
R15697 w_4660_n6791.n2655 w_4660_n6791.n2654 27.1064
R15698 w_4660_n6791.n2654 w_4660_n6791.n105 27.1064
R15699 w_4660_n6791.n964 w_4660_n6791.n105 27.1064
R15700 w_4660_n6791.n964 w_4660_n6791.n957 27.1064
R15701 w_4660_n6791.n970 w_4660_n6791.n957 27.1064
R15702 w_4660_n6791.n971 w_4660_n6791.n970 27.1064
R15703 w_4660_n6791.n972 w_4660_n6791.n971 27.1064
R15704 w_4660_n6791.n972 w_4660_n6791.n949 27.1064
R15705 w_4660_n6791.n978 w_4660_n6791.n949 27.1064
R15706 w_4660_n6791.n979 w_4660_n6791.n978 27.1064
R15707 w_4660_n6791.n981 w_4660_n6791.n979 27.1064
R15708 w_4660_n6791.n981 w_4660_n6791.n980 27.1064
R15709 w_4660_n6791.n980 w_4660_n6791.n945 27.1064
R15710 w_4660_n6791.n941 w_4660_n6791.n940 27.1064
R15711 w_4660_n6791.n940 w_4660_n6791.n503 27.1064
R15712 w_4660_n6791.n503 w_4660_n6791.n502 27.1064
R15713 w_4660_n6791.n502 w_4660_n6791.n499 27.1064
R15714 w_4660_n6791.n499 w_4660_n6791.n498 27.1064
R15715 w_4660_n6791.n498 w_4660_n6791.n495 27.1064
R15716 w_4660_n6791.n495 w_4660_n6791.n494 27.1064
R15717 w_4660_n6791.n494 w_4660_n6791.n491 27.1064
R15718 w_4660_n6791.n491 w_4660_n6791.n490 27.1064
R15719 w_4660_n6791.n490 w_4660_n6791.n487 27.1064
R15720 w_4660_n6791.n487 w_4660_n6791.n486 27.1064
R15721 w_4660_n6791.n486 w_4660_n6791.n483 27.1064
R15722 w_4660_n6791.n483 w_4660_n6791.n482 27.1064
R15723 w_4660_n6791.n482 w_4660_n6791.n479 27.1064
R15724 w_4660_n6791.n479 w_4660_n6791.n478 27.1064
R15725 w_4660_n6791.n478 w_4660_n6791.n475 27.1064
R15726 w_4660_n6791.n475 w_4660_n6791.n474 27.1064
R15727 w_4660_n6791.n474 w_4660_n6791.n471 27.1064
R15728 w_4660_n6791.n471 w_4660_n6791.n470 27.1064
R15729 w_4660_n6791.n470 w_4660_n6791.n467 27.1064
R15730 w_4660_n6791.n467 w_4660_n6791.n462 27.1064
R15731 w_4660_n6791.n1468 w_4660_n6791.n462 27.1064
R15732 w_4660_n6791.n1469 w_4660_n6791.n1468 27.1064
R15733 w_4660_n6791.n1472 w_4660_n6791.n1469 27.1064
R15734 w_4660_n6791.n1470 w_4660_n6791.n456 27.1064
R15735 w_4660_n6791.n1478 w_4660_n6791.n456 27.1064
R15736 w_4660_n6791.n1479 w_4660_n6791.n1478 27.1064
R15737 w_4660_n6791.n1482 w_4660_n6791.n1479 27.1064
R15738 w_4660_n6791.n1483 w_4660_n6791.n1482 27.1064
R15739 w_4660_n6791.n1486 w_4660_n6791.n1483 27.1064
R15740 w_4660_n6791.n1487 w_4660_n6791.n1486 27.1064
R15741 w_4660_n6791.n1490 w_4660_n6791.n1487 27.1064
R15742 w_4660_n6791.n1491 w_4660_n6791.n1490 27.1064
R15743 w_4660_n6791.n1493 w_4660_n6791.n1491 27.1064
R15744 w_4660_n6791.n1495 w_4660_n6791.n1493 27.1064
R15745 w_4660_n6791.n1495 w_4660_n6791.n1494 27.1064
R15746 w_4660_n6791.n1494 w_4660_n6791.n119 27.1064
R15747 w_4660_n6791.n123 w_4660_n6791.n119 27.1064
R15748 w_4660_n6791.n124 w_4660_n6791.n123 27.1064
R15749 w_4660_n6791.n127 w_4660_n6791.n124 27.1064
R15750 w_4660_n6791.n128 w_4660_n6791.n127 27.1064
R15751 w_4660_n6791.n131 w_4660_n6791.n128 27.1064
R15752 w_4660_n6791.n132 w_4660_n6791.n131 27.1064
R15753 w_4660_n6791.n135 w_4660_n6791.n132 27.1064
R15754 w_4660_n6791.n136 w_4660_n6791.n135 27.1064
R15755 w_4660_n6791.n139 w_4660_n6791.n136 27.1064
R15756 w_4660_n6791.n140 w_4660_n6791.n139 27.1064
R15757 w_4660_n6791.n255 w_4660_n6791.n140 27.1064
R15758 w_4660_n6791.n2516 w_4660_n6791.n257 27.1064
R15759 w_4660_n6791.n2516 w_4660_n6791.n2515 27.1064
R15760 w_4660_n6791.n2515 w_4660_n6791.n2514 27.1064
R15761 w_4660_n6791.n2514 w_4660_n6791.n258 27.1064
R15762 w_4660_n6791.n2508 w_4660_n6791.n258 27.1064
R15763 w_4660_n6791.n2508 w_4660_n6791.n2507 27.1064
R15764 w_4660_n6791.n2507 w_4660_n6791.n2506 27.1064
R15765 w_4660_n6791.n2506 w_4660_n6791.n266 27.1064
R15766 w_4660_n6791.n2500 w_4660_n6791.n266 27.1064
R15767 w_4660_n6791.n2500 w_4660_n6791.n2499 27.1064
R15768 w_4660_n6791.n2499 w_4660_n6791.n2498 27.1064
R15769 w_4660_n6791.n2498 w_4660_n6791.n274 27.1064
R15770 w_4660_n6791.n2492 w_4660_n6791.n274 27.1064
R15771 w_4660_n6791.n2492 w_4660_n6791.n2491 27.1064
R15772 w_4660_n6791.n2491 w_4660_n6791.n2490 27.1064
R15773 w_4660_n6791.n2490 w_4660_n6791.n282 27.1064
R15774 w_4660_n6791.n2484 w_4660_n6791.n282 27.1064
R15775 w_4660_n6791.n2484 w_4660_n6791.n2483 27.1064
R15776 w_4660_n6791.n2483 w_4660_n6791.n2482 27.1064
R15777 w_4660_n6791.n2482 w_4660_n6791.n291 27.1064
R15778 w_4660_n6791.n2476 w_4660_n6791.n291 27.1064
R15779 w_4660_n6791.n2476 w_4660_n6791.n2475 27.1064
R15780 w_4660_n6791.n1767 w_4660_n6791.n448 27.1064
R15781 w_4660_n6791.n1768 w_4660_n6791.n1767 27.1064
R15782 w_4660_n6791.n1772 w_4660_n6791.n1768 27.1064
R15783 w_4660_n6791.n1773 w_4660_n6791.n1772 27.1064
R15784 w_4660_n6791.n1775 w_4660_n6791.n1773 27.1064
R15785 w_4660_n6791.n1776 w_4660_n6791.n1775 27.1064
R15786 w_4660_n6791.n1779 w_4660_n6791.n1776 27.1064
R15787 w_4660_n6791.n1780 w_4660_n6791.n1779 27.1064
R15788 w_4660_n6791.n1784 w_4660_n6791.n1780 27.1064
R15789 w_4660_n6791.n1785 w_4660_n6791.n1784 27.1064
R15790 w_4660_n6791.n1789 w_4660_n6791.n1785 27.1064
R15791 w_4660_n6791.n1790 w_4660_n6791.n1789 27.1064
R15792 w_4660_n6791.n1793 w_4660_n6791.n1790 27.1064
R15793 w_4660_n6791.n1794 w_4660_n6791.n1793 27.1064
R15794 w_4660_n6791.n1798 w_4660_n6791.n1794 27.1064
R15795 w_4660_n6791.n1799 w_4660_n6791.n1798 27.1064
R15796 w_4660_n6791.n1803 w_4660_n6791.n1799 27.1064
R15797 w_4660_n6791.n1804 w_4660_n6791.n1803 27.1064
R15798 w_4660_n6791.n1808 w_4660_n6791.n1804 27.1064
R15799 w_4660_n6791.n1809 w_4660_n6791.n1808 27.1064
R15800 w_4660_n6791.n1812 w_4660_n6791.n1809 27.1064
R15801 w_4660_n6791.n1813 w_4660_n6791.n1812 27.1064
R15802 w_4660_n6791.n1816 w_4660_n6791.n1813 27.1064
R15803 w_4660_n6791.n1817 w_4660_n6791.n1816 27.1064
R15804 w_4660_n6791.n1821 w_4660_n6791.n1817 27.1064
R15805 w_4660_n6791.n1822 w_4660_n6791.n1821 27.1064
R15806 w_4660_n6791.n1825 w_4660_n6791.n1822 27.1064
R15807 w_4660_n6791.n1826 w_4660_n6791.n1825 27.1064
R15808 w_4660_n6791.n1828 w_4660_n6791.n1826 27.1064
R15809 w_4660_n6791.n1829 w_4660_n6791.n1828 27.1064
R15810 w_4660_n6791.n1832 w_4660_n6791.n1829 27.1064
R15811 w_4660_n6791.n1833 w_4660_n6791.n1832 27.1064
R15812 w_4660_n6791.n1837 w_4660_n6791.n1833 27.1064
R15813 w_4660_n6791.n1838 w_4660_n6791.n1837 27.1064
R15814 w_4660_n6791.n1842 w_4660_n6791.n1838 27.1064
R15815 w_4660_n6791.n1843 w_4660_n6791.n1842 27.1064
R15816 w_4660_n6791.n1847 w_4660_n6791.n1843 27.1064
R15817 w_4660_n6791.n1848 w_4660_n6791.n1847 27.1064
R15818 w_4660_n6791.n1851 w_4660_n6791.n1848 27.1064
R15819 w_4660_n6791.n1852 w_4660_n6791.n1851 27.1064
R15820 w_4660_n6791.n1856 w_4660_n6791.n1855 27.1064
R15821 w_4660_n6791.n1860 w_4660_n6791.n1856 27.1064
R15822 w_4660_n6791.n1861 w_4660_n6791.n1860 27.1064
R15823 w_4660_n6791.n1865 w_4660_n6791.n1861 27.1064
R15824 w_4660_n6791.n1866 w_4660_n6791.n1865 27.1064
R15825 w_4660_n6791.n1870 w_4660_n6791.n1866 27.1064
R15826 w_4660_n6791.n1871 w_4660_n6791.n1870 27.1064
R15827 w_4660_n6791.n1874 w_4660_n6791.n1871 27.1064
R15828 w_4660_n6791.n1875 w_4660_n6791.n1874 27.1064
R15829 w_4660_n6791.n1878 w_4660_n6791.n1875 27.1064
R15830 w_4660_n6791.n1879 w_4660_n6791.n1878 27.1064
R15831 w_4660_n6791.n1883 w_4660_n6791.n1879 27.1064
R15832 w_4660_n6791.n1884 w_4660_n6791.n1883 27.1064
R15833 w_4660_n6791.n1888 w_4660_n6791.n1884 27.1064
R15834 w_4660_n6791.n1889 w_4660_n6791.n1888 27.1064
R15835 w_4660_n6791.n1892 w_4660_n6791.n1889 27.1064
R15836 w_4660_n6791.n1893 w_4660_n6791.n1892 27.1064
R15837 w_4660_n6791.n1896 w_4660_n6791.n1893 27.1064
R15838 w_4660_n6791.n1897 w_4660_n6791.n1896 27.1064
R15839 w_4660_n6791.n1901 w_4660_n6791.n1897 27.1064
R15840 w_4660_n6791.n1902 w_4660_n6791.n1901 27.1064
R15841 w_4660_n6791.n1905 w_4660_n6791.n1902 27.1064
R15842 w_4660_n6791.n1906 w_4660_n6791.n1905 27.1064
R15843 w_4660_n6791.n1908 w_4660_n6791.n1906 27.1064
R15844 w_4660_n6791.n1909 w_4660_n6791.n1908 27.1064
R15845 w_4660_n6791.n1912 w_4660_n6791.n1909 27.1064
R15846 w_4660_n6791.n1913 w_4660_n6791.n1912 27.1064
R15847 w_4660_n6791.n1916 w_4660_n6791.n1913 27.1064
R15848 w_4660_n6791.n1917 w_4660_n6791.n1916 27.1064
R15849 w_4660_n6791.n2113 w_4660_n6791.n1917 27.1064
R15850 w_4660_n6791.n2114 w_4660_n6791.n2113 27.1064
R15851 w_4660_n6791.n2116 w_4660_n6791.n2114 27.1064
R15852 w_4660_n6791.n2116 w_4660_n6791.n2115 27.1064
R15853 w_4660_n6791.n2115 w_4660_n6791.n48 27.1064
R15854 w_4660_n6791.n53 w_4660_n6791.n48 27.1064
R15855 w_4660_n6791.n54 w_4660_n6791.n53 27.1064
R15856 w_4660_n6791.n58 w_4660_n6791.n54 27.1064
R15857 w_4660_n6791.n59 w_4660_n6791.n58 27.1064
R15858 w_4660_n6791.n62 w_4660_n6791.n59 27.1064
R15859 w_4660_n6791.n63 w_4660_n6791.n62 27.1064
R15860 w_4660_n6791.n82 w_4660_n6791.n63 27.1064
R15861 w_4660_n6791.n2263 w_4660_n6791.n1765 27.1064
R15862 w_4660_n6791.n2263 w_4660_n6791.n2262 27.1064
R15863 w_4660_n6791.n2262 w_4660_n6791.n2261 27.1064
R15864 w_4660_n6791.n2261 w_4660_n6791.n1766 27.1064
R15865 w_4660_n6791.n2255 w_4660_n6791.n1766 27.1064
R15866 w_4660_n6791.n2255 w_4660_n6791.n2254 27.1064
R15867 w_4660_n6791.n2254 w_4660_n6791.n2253 27.1064
R15868 w_4660_n6791.n2253 w_4660_n6791.n1774 27.1064
R15869 w_4660_n6791.n2248 w_4660_n6791.n1774 27.1064
R15870 w_4660_n6791.n2248 w_4660_n6791.n2247 27.1064
R15871 w_4660_n6791.n2247 w_4660_n6791.n2246 27.1064
R15872 w_4660_n6791.n2246 w_4660_n6791.n1782 27.1064
R15873 w_4660_n6791.n2240 w_4660_n6791.n1782 27.1064
R15874 w_4660_n6791.n2240 w_4660_n6791.n2239 27.1064
R15875 w_4660_n6791.n2239 w_4660_n6791.n1792 27.1064
R15876 w_4660_n6791.n1801 w_4660_n6791.n1792 27.1064
R15877 w_4660_n6791.n2232 w_4660_n6791.n1801 27.1064
R15878 w_4660_n6791.n2232 w_4660_n6791.n2231 27.1064
R15879 w_4660_n6791.n2231 w_4660_n6791.n2230 27.1064
R15880 w_4660_n6791.n2230 w_4660_n6791.n1802 27.1064
R15881 w_4660_n6791.n2224 w_4660_n6791.n1802 27.1064
R15882 w_4660_n6791.n2224 w_4660_n6791.n2223 27.1064
R15883 w_4660_n6791.n2223 w_4660_n6791.n2222 27.1064
R15884 w_4660_n6791.n2222 w_4660_n6791.n1811 27.1064
R15885 w_4660_n6791.n2216 w_4660_n6791.n1811 27.1064
R15886 w_4660_n6791.n2216 w_4660_n6791.n2215 27.1064
R15887 w_4660_n6791.n2215 w_4660_n6791.n2214 27.1064
R15888 w_4660_n6791.n2214 w_4660_n6791.n1819 27.1064
R15889 w_4660_n6791.n2208 w_4660_n6791.n1819 27.1064
R15890 w_4660_n6791.n2208 w_4660_n6791.n2207 27.1064
R15891 w_4660_n6791.n2207 w_4660_n6791.n1827 27.1064
R15892 w_4660_n6791.n1835 w_4660_n6791.n1827 27.1064
R15893 w_4660_n6791.n2201 w_4660_n6791.n1835 27.1064
R15894 w_4660_n6791.n2201 w_4660_n6791.n2200 27.1064
R15895 w_4660_n6791.n2200 w_4660_n6791.n1836 27.1064
R15896 w_4660_n6791.n1845 w_4660_n6791.n1836 27.1064
R15897 w_4660_n6791.n2193 w_4660_n6791.n1845 27.1064
R15898 w_4660_n6791.n2193 w_4660_n6791.n2192 27.1064
R15899 w_4660_n6791.n2192 w_4660_n6791.n2191 27.1064
R15900 w_4660_n6791.n2191 w_4660_n6791.n1846 27.1064
R15901 w_4660_n6791.n2185 w_4660_n6791.n1846 27.1064
R15902 w_4660_n6791.n2183 w_4660_n6791.n2182 27.1064
R15903 w_4660_n6791.n2182 w_4660_n6791.n1854 27.1064
R15904 w_4660_n6791.n2176 w_4660_n6791.n1854 27.1064
R15905 w_4660_n6791.n2176 w_4660_n6791.n2175 27.1064
R15906 w_4660_n6791.n2175 w_4660_n6791.n2174 27.1064
R15907 w_4660_n6791.n2174 w_4660_n6791.n1863 27.1064
R15908 w_4660_n6791.n2168 w_4660_n6791.n1863 27.1064
R15909 w_4660_n6791.n2168 w_4660_n6791.n2167 27.1064
R15910 w_4660_n6791.n2167 w_4660_n6791.n1873 27.1064
R15911 w_4660_n6791.n1881 w_4660_n6791.n1873 27.1064
R15912 w_4660_n6791.n2160 w_4660_n6791.n1881 27.1064
R15913 w_4660_n6791.n2160 w_4660_n6791.n2159 27.1064
R15914 w_4660_n6791.n2159 w_4660_n6791.n2158 27.1064
R15915 w_4660_n6791.n2158 w_4660_n6791.n1882 27.1064
R15916 w_4660_n6791.n2152 w_4660_n6791.n1882 27.1064
R15917 w_4660_n6791.n2152 w_4660_n6791.n2151 27.1064
R15918 w_4660_n6791.n2151 w_4660_n6791.n2150 27.1064
R15919 w_4660_n6791.n2150 w_4660_n6791.n1891 27.1064
R15920 w_4660_n6791.n2144 w_4660_n6791.n1891 27.1064
R15921 w_4660_n6791.n2144 w_4660_n6791.n2143 27.1064
R15922 w_4660_n6791.n2143 w_4660_n6791.n2142 27.1064
R15923 w_4660_n6791.n2142 w_4660_n6791.n1899 27.1064
R15924 w_4660_n6791.n2136 w_4660_n6791.n1899 27.1064
R15925 w_4660_n6791.n2136 w_4660_n6791.n2135 27.1064
R15926 w_4660_n6791.n2135 w_4660_n6791.n2134 27.1064
R15927 w_4660_n6791.n2134 w_4660_n6791.n1907 27.1064
R15928 w_4660_n6791.n2128 w_4660_n6791.n1907 27.1064
R15929 w_4660_n6791.n2128 w_4660_n6791.n2127 27.1064
R15930 w_4660_n6791.n2127 w_4660_n6791.n1915 27.1064
R15931 w_4660_n6791.n2118 w_4660_n6791.n1915 27.1064
R15932 w_4660_n6791.n2120 w_4660_n6791.n2118 27.1064
R15933 w_4660_n6791.n2120 w_4660_n6791.n2119 27.1064
R15934 w_4660_n6791.n2119 w_4660_n6791.n51 27.1064
R15935 w_4660_n6791.n2694 w_4660_n6791.n51 27.1064
R15936 w_4660_n6791.n2694 w_4660_n6791.n2693 27.1064
R15937 w_4660_n6791.n2693 w_4660_n6791.n2692 27.1064
R15938 w_4660_n6791.n2692 w_4660_n6791.n52 27.1064
R15939 w_4660_n6791.n2686 w_4660_n6791.n52 27.1064
R15940 w_4660_n6791.n2686 w_4660_n6791.n2685 27.1064
R15941 w_4660_n6791.n2685 w_4660_n6791.n2684 27.1064
R15942 w_4660_n6791.n2684 w_4660_n6791.n61 27.1064
R15943 w_4660_n6791.n1219 w_4660_n6791.n451 27.1064
R15944 w_4660_n6791.n1219 w_4660_n6791.n1218 27.1064
R15945 w_4660_n6791.n1218 w_4660_n6791.n1141 27.1064
R15946 w_4660_n6791.n1141 w_4660_n6791.n1135 27.1064
R15947 w_4660_n6791.n1231 w_4660_n6791.n1135 27.1064
R15948 w_4660_n6791.n1232 w_4660_n6791.n1231 27.1064
R15949 w_4660_n6791.n1233 w_4660_n6791.n1232 27.1064
R15950 w_4660_n6791.n1233 w_4660_n6791.n1132 27.1064
R15951 w_4660_n6791.n1132 w_4660_n6791.n1131 27.1064
R15952 w_4660_n6791.n1131 w_4660_n6791.n1123 27.1064
R15953 w_4660_n6791.n1245 w_4660_n6791.n1123 27.1064
R15954 w_4660_n6791.n1246 w_4660_n6791.n1245 27.1064
R15955 w_4660_n6791.n1247 w_4660_n6791.n1246 27.1064
R15956 w_4660_n6791.n1247 w_4660_n6791.n1120 27.1064
R15957 w_4660_n6791.n1120 w_4660_n6791.n1119 27.1064
R15958 w_4660_n6791.n1119 w_4660_n6791.n1116 27.1064
R15959 w_4660_n6791.n1116 w_4660_n6791.n1115 27.1064
R15960 w_4660_n6791.n1115 w_4660_n6791.n1112 27.1064
R15961 w_4660_n6791.n1112 w_4660_n6791.n1111 27.1064
R15962 w_4660_n6791.n1111 w_4660_n6791.n1105 27.1064
R15963 w_4660_n6791.n1267 w_4660_n6791.n1105 27.1064
R15964 w_4660_n6791.n1268 w_4660_n6791.n1267 27.1064
R15965 w_4660_n6791.n1269 w_4660_n6791.n1268 27.1064
R15966 w_4660_n6791.n1269 w_4660_n6791.n1102 27.1064
R15967 w_4660_n6791.n1102 w_4660_n6791.n1101 27.1064
R15968 w_4660_n6791.n1101 w_4660_n6791.n1097 27.1064
R15969 w_4660_n6791.n1097 w_4660_n6791.n1091 27.1064
R15970 w_4660_n6791.n1283 w_4660_n6791.n1091 27.1064
R15971 w_4660_n6791.n1284 w_4660_n6791.n1283 27.1064
R15972 w_4660_n6791.n1285 w_4660_n6791.n1284 27.1064
R15973 w_4660_n6791.n1285 w_4660_n6791.n1088 27.1064
R15974 w_4660_n6791.n1088 w_4660_n6791.n1087 27.1064
R15975 w_4660_n6791.n1087 w_4660_n6791.n1079 27.1064
R15976 w_4660_n6791.n1297 w_4660_n6791.n1079 27.1064
R15977 w_4660_n6791.n1298 w_4660_n6791.n1297 27.1064
R15978 w_4660_n6791.n1299 w_4660_n6791.n1298 27.1064
R15979 w_4660_n6791.n1299 w_4660_n6791.n1076 27.1064
R15980 w_4660_n6791.n1076 w_4660_n6791.n1075 27.1064
R15981 w_4660_n6791.n1075 w_4660_n6791.n1067 27.1064
R15982 w_4660_n6791.n1312 w_4660_n6791.n1067 27.1064
R15983 w_4660_n6791.n1313 w_4660_n6791.n1312 27.1064
R15984 w_4660_n6791.n1315 w_4660_n6791.n1061 27.1064
R15985 w_4660_n6791.n1323 w_4660_n6791.n1061 27.1064
R15986 w_4660_n6791.n1324 w_4660_n6791.n1323 27.1064
R15987 w_4660_n6791.n1325 w_4660_n6791.n1324 27.1064
R15988 w_4660_n6791.n1325 w_4660_n6791.n1058 27.1064
R15989 w_4660_n6791.n1058 w_4660_n6791.n1057 27.1064
R15990 w_4660_n6791.n1057 w_4660_n6791.n1053 27.1064
R15991 w_4660_n6791.n1053 w_4660_n6791.n1047 27.1064
R15992 w_4660_n6791.n1339 w_4660_n6791.n1047 27.1064
R15993 w_4660_n6791.n1340 w_4660_n6791.n1339 27.1064
R15994 w_4660_n6791.n1341 w_4660_n6791.n1340 27.1064
R15995 w_4660_n6791.n1341 w_4660_n6791.n1044 27.1064
R15996 w_4660_n6791.n1044 w_4660_n6791.n1043 27.1064
R15997 w_4660_n6791.n1043 w_4660_n6791.n1037 27.1064
R15998 w_4660_n6791.n1352 w_4660_n6791.n1037 27.1064
R15999 w_4660_n6791.n1353 w_4660_n6791.n1352 27.1064
R16000 w_4660_n6791.n1354 w_4660_n6791.n1353 27.1064
R16001 w_4660_n6791.n1354 w_4660_n6791.n1034 27.1064
R16002 w_4660_n6791.n1034 w_4660_n6791.n1033 27.1064
R16003 w_4660_n6791.n1033 w_4660_n6791.n1029 27.1064
R16004 w_4660_n6791.n1029 w_4660_n6791.n1023 27.1064
R16005 w_4660_n6791.n1368 w_4660_n6791.n1023 27.1064
R16006 w_4660_n6791.n1369 w_4660_n6791.n1368 27.1064
R16007 w_4660_n6791.n1370 w_4660_n6791.n1369 27.1064
R16008 w_4660_n6791.n1370 w_4660_n6791.n1020 27.1064
R16009 w_4660_n6791.n1020 w_4660_n6791.n1019 27.1064
R16010 w_4660_n6791.n1019 w_4660_n6791.n1011 27.1064
R16011 w_4660_n6791.n1382 w_4660_n6791.n1011 27.1064
R16012 w_4660_n6791.n1383 w_4660_n6791.n1382 27.1064
R16013 w_4660_n6791.n1384 w_4660_n6791.n1383 27.1064
R16014 w_4660_n6791.n1384 w_4660_n6791.n1008 27.1064
R16015 w_4660_n6791.n1008 w_4660_n6791.n1007 27.1064
R16016 w_4660_n6791.n1007 w_4660_n6791.n1004 27.1064
R16017 w_4660_n6791.n1004 w_4660_n6791.n15 27.1064
R16018 w_4660_n6791.n1398 w_4660_n6791.n15 27.1064
R16019 w_4660_n6791.n1399 w_4660_n6791.n1398 27.1064
R16020 w_4660_n6791.n1400 w_4660_n6791.n1399 27.1064
R16021 w_4660_n6791.n1400 w_4660_n6791.n997 27.1064
R16022 w_4660_n6791.n997 w_4660_n6791.n996 27.1064
R16023 w_4660_n6791.n996 w_4660_n6791.n986 27.1064
R16024 w_4660_n6791.n1412 w_4660_n6791.n986 27.1064
R16025 w_4660_n6791.n1223 w_4660_n6791.n1222 27.1064
R16026 w_4660_n6791.n1225 w_4660_n6791.n1223 27.1064
R16027 w_4660_n6791.n1225 w_4660_n6791.n1224 27.1064
R16028 w_4660_n6791.n1224 w_4660_n6791.n1138 27.1064
R16029 w_4660_n6791.n1138 w_4660_n6791.n1137 27.1064
R16030 w_4660_n6791.n1137 w_4660_n6791.n1129 27.1064
R16031 w_4660_n6791.n1238 w_4660_n6791.n1129 27.1064
R16032 w_4660_n6791.n1239 w_4660_n6791.n1238 27.1064
R16033 w_4660_n6791.n1240 w_4660_n6791.n1239 27.1064
R16034 w_4660_n6791.n1240 w_4660_n6791.n1126 27.1064
R16035 w_4660_n6791.n1126 w_4660_n6791.n1125 27.1064
R16036 w_4660_n6791.n1125 w_4660_n6791.n1117 27.1064
R16037 w_4660_n6791.n1252 w_4660_n6791.n1117 27.1064
R16038 w_4660_n6791.n1253 w_4660_n6791.n1252 27.1064
R16039 w_4660_n6791.n1254 w_4660_n6791.n1253 27.1064
R16040 w_4660_n6791.n1254 w_4660_n6791.n11 27.1064
R16041 w_4660_n6791.n1260 w_4660_n6791.n11 27.1064
R16042 w_4660_n6791.n1261 w_4660_n6791.n1260 27.1064
R16043 w_4660_n6791.n1262 w_4660_n6791.n1261 27.1064
R16044 w_4660_n6791.n1262 w_4660_n6791.n1108 27.1064
R16045 w_4660_n6791.n1108 w_4660_n6791.n1107 27.1064
R16046 w_4660_n6791.n1107 w_4660_n6791.n1099 27.1064
R16047 w_4660_n6791.n1274 w_4660_n6791.n1099 27.1064
R16048 w_4660_n6791.n1275 w_4660_n6791.n1274 27.1064
R16049 w_4660_n6791.n1277 w_4660_n6791.n1275 27.1064
R16050 w_4660_n6791.n1277 w_4660_n6791.n1276 27.1064
R16051 w_4660_n6791.n1276 w_4660_n6791.n1094 27.1064
R16052 w_4660_n6791.n1094 w_4660_n6791.n1093 27.1064
R16053 w_4660_n6791.n1093 w_4660_n6791.n1085 27.1064
R16054 w_4660_n6791.n1290 w_4660_n6791.n1085 27.1064
R16055 w_4660_n6791.n1291 w_4660_n6791.n1290 27.1064
R16056 w_4660_n6791.n1292 w_4660_n6791.n1291 27.1064
R16057 w_4660_n6791.n1292 w_4660_n6791.n1082 27.1064
R16058 w_4660_n6791.n1082 w_4660_n6791.n1081 27.1064
R16059 w_4660_n6791.n1081 w_4660_n6791.n1073 27.1064
R16060 w_4660_n6791.n1304 w_4660_n6791.n1073 27.1064
R16061 w_4660_n6791.n1305 w_4660_n6791.n1304 27.1064
R16062 w_4660_n6791.n1306 w_4660_n6791.n1305 27.1064
R16063 w_4660_n6791.n1306 w_4660_n6791.n1070 27.1064
R16064 w_4660_n6791.n1070 w_4660_n6791.n1069 27.1064
R16065 w_4660_n6791.n1318 w_4660_n6791.n1317 27.1064
R16066 w_4660_n6791.n1318 w_4660_n6791.n1064 27.1064
R16067 w_4660_n6791.n1064 w_4660_n6791.n1063 27.1064
R16068 w_4660_n6791.n1063 w_4660_n6791.n1055 27.1064
R16069 w_4660_n6791.n1330 w_4660_n6791.n1055 27.1064
R16070 w_4660_n6791.n1331 w_4660_n6791.n1330 27.1064
R16071 w_4660_n6791.n1333 w_4660_n6791.n1331 27.1064
R16072 w_4660_n6791.n1333 w_4660_n6791.n1332 27.1064
R16073 w_4660_n6791.n1332 w_4660_n6791.n1050 27.1064
R16074 w_4660_n6791.n1050 w_4660_n6791.n1049 27.1064
R16075 w_4660_n6791.n1049 w_4660_n6791.n13 27.1064
R16076 w_4660_n6791.n1345 w_4660_n6791.n13 27.1064
R16077 w_4660_n6791.n1346 w_4660_n6791.n1345 27.1064
R16078 w_4660_n6791.n1347 w_4660_n6791.n1346 27.1064
R16079 w_4660_n6791.n1347 w_4660_n6791.n1040 27.1064
R16080 w_4660_n6791.n1040 w_4660_n6791.n1039 27.1064
R16081 w_4660_n6791.n1039 w_4660_n6791.n1031 27.1064
R16082 w_4660_n6791.n1359 w_4660_n6791.n1031 27.1064
R16083 w_4660_n6791.n1360 w_4660_n6791.n1359 27.1064
R16084 w_4660_n6791.n1362 w_4660_n6791.n1360 27.1064
R16085 w_4660_n6791.n1362 w_4660_n6791.n1361 27.1064
R16086 w_4660_n6791.n1361 w_4660_n6791.n1026 27.1064
R16087 w_4660_n6791.n1026 w_4660_n6791.n1025 27.1064
R16088 w_4660_n6791.n1025 w_4660_n6791.n1017 27.1064
R16089 w_4660_n6791.n1375 w_4660_n6791.n1017 27.1064
R16090 w_4660_n6791.n1376 w_4660_n6791.n1375 27.1064
R16091 w_4660_n6791.n1377 w_4660_n6791.n1376 27.1064
R16092 w_4660_n6791.n1377 w_4660_n6791.n1014 27.1064
R16093 w_4660_n6791.n1014 w_4660_n6791.n1013 27.1064
R16094 w_4660_n6791.n1013 w_4660_n6791.n1005 27.1064
R16095 w_4660_n6791.n1389 w_4660_n6791.n1005 27.1064
R16096 w_4660_n6791.n1390 w_4660_n6791.n1389 27.1064
R16097 w_4660_n6791.n1392 w_4660_n6791.n1390 27.1064
R16098 w_4660_n6791.n1392 w_4660_n6791.n1391 27.1064
R16099 w_4660_n6791.n1391 w_4660_n6791.n1001 27.1064
R16100 w_4660_n6791.n1001 w_4660_n6791.n1000 27.1064
R16101 w_4660_n6791.n1000 w_4660_n6791.n994 27.1064
R16102 w_4660_n6791.n1405 w_4660_n6791.n994 27.1064
R16103 w_4660_n6791.n1406 w_4660_n6791.n1405 27.1064
R16104 w_4660_n6791.n1407 w_4660_n6791.n1406 27.1064
R16105 w_4660_n6791.n1407 w_4660_n6791.n991 27.1064
R16106 w_4660_n6791.n1220 w_4660_n6791.n1139 27.1064
R16107 w_4660_n6791.n1227 w_4660_n6791.n1139 27.1064
R16108 w_4660_n6791.n1228 w_4660_n6791.n1227 27.1064
R16109 w_4660_n6791.n1229 w_4660_n6791.n1228 27.1064
R16110 w_4660_n6791.n1229 w_4660_n6791.n1133 27.1064
R16111 w_4660_n6791.n1235 w_4660_n6791.n1133 27.1064
R16112 w_4660_n6791.n1236 w_4660_n6791.n1235 27.1064
R16113 w_4660_n6791.n1236 w_4660_n6791.n1127 27.1064
R16114 w_4660_n6791.n1242 w_4660_n6791.n1127 27.1064
R16115 w_4660_n6791.n1243 w_4660_n6791.n1242 27.1064
R16116 w_4660_n6791.n1243 w_4660_n6791.n1121 27.1064
R16117 w_4660_n6791.n1249 w_4660_n6791.n1121 27.1064
R16118 w_4660_n6791.n1250 w_4660_n6791.n1249 27.1064
R16119 w_4660_n6791.n1250 w_4660_n6791.n1113 27.1064
R16120 w_4660_n6791.n1256 w_4660_n6791.n1113 27.1064
R16121 w_4660_n6791.n1257 w_4660_n6791.n1256 27.1064
R16122 w_4660_n6791.n1258 w_4660_n6791.n1257 27.1064
R16123 w_4660_n6791.n1258 w_4660_n6791.n1109 27.1064
R16124 w_4660_n6791.n1264 w_4660_n6791.n1109 27.1064
R16125 w_4660_n6791.n1265 w_4660_n6791.n1264 27.1064
R16126 w_4660_n6791.n1265 w_4660_n6791.n1103 27.1064
R16127 w_4660_n6791.n1271 w_4660_n6791.n1103 27.1064
R16128 w_4660_n6791.n1272 w_4660_n6791.n1271 27.1064
R16129 w_4660_n6791.n1272 w_4660_n6791.n1095 27.1064
R16130 w_4660_n6791.n1279 w_4660_n6791.n1095 27.1064
R16131 w_4660_n6791.n1280 w_4660_n6791.n1279 27.1064
R16132 w_4660_n6791.n1281 w_4660_n6791.n1280 27.1064
R16133 w_4660_n6791.n1281 w_4660_n6791.n1089 27.1064
R16134 w_4660_n6791.n1287 w_4660_n6791.n1089 27.1064
R16135 w_4660_n6791.n1288 w_4660_n6791.n1287 27.1064
R16136 w_4660_n6791.n1288 w_4660_n6791.n1083 27.1064
R16137 w_4660_n6791.n1294 w_4660_n6791.n1083 27.1064
R16138 w_4660_n6791.n1295 w_4660_n6791.n1294 27.1064
R16139 w_4660_n6791.n1295 w_4660_n6791.n1077 27.1064
R16140 w_4660_n6791.n1301 w_4660_n6791.n1077 27.1064
R16141 w_4660_n6791.n1302 w_4660_n6791.n1301 27.1064
R16142 w_4660_n6791.n1302 w_4660_n6791.n1071 27.1064
R16143 w_4660_n6791.n1308 w_4660_n6791.n1071 27.1064
R16144 w_4660_n6791.n1310 w_4660_n6791.n1308 27.1064
R16145 w_4660_n6791.n1310 w_4660_n6791.n1309 27.1064
R16146 w_4660_n6791.n1320 w_4660_n6791.n1065 27.1064
R16147 w_4660_n6791.n1321 w_4660_n6791.n1320 27.1064
R16148 w_4660_n6791.n1321 w_4660_n6791.n1059 27.1064
R16149 w_4660_n6791.n1327 w_4660_n6791.n1059 27.1064
R16150 w_4660_n6791.n1328 w_4660_n6791.n1327 27.1064
R16151 w_4660_n6791.n1328 w_4660_n6791.n1051 27.1064
R16152 w_4660_n6791.n1335 w_4660_n6791.n1051 27.1064
R16153 w_4660_n6791.n1336 w_4660_n6791.n1335 27.1064
R16154 w_4660_n6791.n1337 w_4660_n6791.n1336 27.1064
R16155 w_4660_n6791.n1337 w_4660_n6791.n1045 27.1064
R16156 w_4660_n6791.n1342 w_4660_n6791.n1045 27.1064
R16157 w_4660_n6791.n1343 w_4660_n6791.n1342 27.1064
R16158 w_4660_n6791.n1343 w_4660_n6791.n1041 27.1064
R16159 w_4660_n6791.n1349 w_4660_n6791.n1041 27.1064
R16160 w_4660_n6791.n1350 w_4660_n6791.n1349 27.1064
R16161 w_4660_n6791.n1350 w_4660_n6791.n1035 27.1064
R16162 w_4660_n6791.n1356 w_4660_n6791.n1035 27.1064
R16163 w_4660_n6791.n1357 w_4660_n6791.n1356 27.1064
R16164 w_4660_n6791.n1357 w_4660_n6791.n1027 27.1064
R16165 w_4660_n6791.n1364 w_4660_n6791.n1027 27.1064
R16166 w_4660_n6791.n1365 w_4660_n6791.n1364 27.1064
R16167 w_4660_n6791.n1366 w_4660_n6791.n1365 27.1064
R16168 w_4660_n6791.n1366 w_4660_n6791.n1021 27.1064
R16169 w_4660_n6791.n1372 w_4660_n6791.n1021 27.1064
R16170 w_4660_n6791.n1373 w_4660_n6791.n1372 27.1064
R16171 w_4660_n6791.n1373 w_4660_n6791.n1015 27.1064
R16172 w_4660_n6791.n1379 w_4660_n6791.n1015 27.1064
R16173 w_4660_n6791.n1380 w_4660_n6791.n1379 27.1064
R16174 w_4660_n6791.n1380 w_4660_n6791.n1009 27.1064
R16175 w_4660_n6791.n1386 w_4660_n6791.n1009 27.1064
R16176 w_4660_n6791.n1387 w_4660_n6791.n1386 27.1064
R16177 w_4660_n6791.n1387 w_4660_n6791.n1002 27.1064
R16178 w_4660_n6791.n1394 w_4660_n6791.n1002 27.1064
R16179 w_4660_n6791.n1395 w_4660_n6791.n1394 27.1064
R16180 w_4660_n6791.n1396 w_4660_n6791.n1395 27.1064
R16181 w_4660_n6791.n1396 w_4660_n6791.n998 27.1064
R16182 w_4660_n6791.n1402 w_4660_n6791.n998 27.1064
R16183 w_4660_n6791.n1403 w_4660_n6791.n1402 27.1064
R16184 w_4660_n6791.n1403 w_4660_n6791.n992 27.1064
R16185 w_4660_n6791.n1409 w_4660_n6791.n992 27.1064
R16186 w_4660_n6791.n1410 w_4660_n6791.n1409 27.1064
R16187 w_4660_n6791.n930 w_4660_n6791.n506 27.1064
R16188 w_4660_n6791.n930 w_4660_n6791.n929 27.1064
R16189 w_4660_n6791.n929 w_4660_n6791.n928 27.1064
R16190 w_4660_n6791.n928 w_4660_n6791.n510 27.1064
R16191 w_4660_n6791.n922 w_4660_n6791.n510 27.1064
R16192 w_4660_n6791.n922 w_4660_n6791.n921 27.1064
R16193 w_4660_n6791.n921 w_4660_n6791.n920 27.1064
R16194 w_4660_n6791.n920 w_4660_n6791.n520 27.1064
R16195 w_4660_n6791.n914 w_4660_n6791.n520 27.1064
R16196 w_4660_n6791.n914 w_4660_n6791.n913 27.1064
R16197 w_4660_n6791.n913 w_4660_n6791.n529 27.1064
R16198 w_4660_n6791.n538 w_4660_n6791.n529 27.1064
R16199 w_4660_n6791.n906 w_4660_n6791.n538 27.1064
R16200 w_4660_n6791.n906 w_4660_n6791.n905 27.1064
R16201 w_4660_n6791.n905 w_4660_n6791.n904 27.1064
R16202 w_4660_n6791.n904 w_4660_n6791.n17 27.1064
R16203 w_4660_n6791.n899 w_4660_n6791.n17 27.1064
R16204 w_4660_n6791.n899 w_4660_n6791.n898 27.1064
R16205 w_4660_n6791.n898 w_4660_n6791.n897 27.1064
R16206 w_4660_n6791.n897 w_4660_n6791.n545 27.1064
R16207 w_4660_n6791.n891 w_4660_n6791.n545 27.1064
R16208 w_4660_n6791.n891 w_4660_n6791.n890 27.1064
R16209 w_4660_n6791.n890 w_4660_n6791.n889 27.1064
R16210 w_4660_n6791.n889 w_4660_n6791.n554 27.1064
R16211 w_4660_n6791.n883 w_4660_n6791.n554 27.1064
R16212 w_4660_n6791.n883 w_4660_n6791.n882 27.1064
R16213 w_4660_n6791.n882 w_4660_n6791.n564 27.1064
R16214 w_4660_n6791.n572 w_4660_n6791.n564 27.1064
R16215 w_4660_n6791.n875 w_4660_n6791.n572 27.1064
R16216 w_4660_n6791.n875 w_4660_n6791.n874 27.1064
R16217 w_4660_n6791.n874 w_4660_n6791.n573 27.1064
R16218 w_4660_n6791.n582 w_4660_n6791.n573 27.1064
R16219 w_4660_n6791.n867 w_4660_n6791.n582 27.1064
R16220 w_4660_n6791.n867 w_4660_n6791.n866 27.1064
R16221 w_4660_n6791.n866 w_4660_n6791.n865 27.1064
R16222 w_4660_n6791.n865 w_4660_n6791.n583 27.1064
R16223 w_4660_n6791.n859 w_4660_n6791.n583 27.1064
R16224 w_4660_n6791.n859 w_4660_n6791.n858 27.1064
R16225 w_4660_n6791.n858 w_4660_n6791.n857 27.1064
R16226 w_4660_n6791.n857 w_4660_n6791.n591 27.1064
R16227 w_4660_n6791.n605 w_4660_n6791.n599 27.1064
R16228 w_4660_n6791.n846 w_4660_n6791.n605 27.1064
R16229 w_4660_n6791.n846 w_4660_n6791.n845 27.1064
R16230 w_4660_n6791.n845 w_4660_n6791.n844 27.1064
R16231 w_4660_n6791.n844 w_4660_n6791.n606 27.1064
R16232 w_4660_n6791.n838 w_4660_n6791.n606 27.1064
R16233 w_4660_n6791.n838 w_4660_n6791.n837 27.1064
R16234 w_4660_n6791.n837 w_4660_n6791.n836 27.1064
R16235 w_4660_n6791.n836 w_4660_n6791.n614 27.1064
R16236 w_4660_n6791.n830 w_4660_n6791.n614 27.1064
R16237 w_4660_n6791.n830 w_4660_n6791.n829 27.1064
R16238 w_4660_n6791.n829 w_4660_n6791.n828 27.1064
R16239 w_4660_n6791.n828 w_4660_n6791.n622 27.1064
R16240 w_4660_n6791.n822 w_4660_n6791.n622 27.1064
R16241 w_4660_n6791.n822 w_4660_n6791.n821 27.1064
R16242 w_4660_n6791.n821 w_4660_n6791.n630 27.1064
R16243 w_4660_n6791.n639 w_4660_n6791.n630 27.1064
R16244 w_4660_n6791.n814 w_4660_n6791.n639 27.1064
R16245 w_4660_n6791.n814 w_4660_n6791.n813 27.1064
R16246 w_4660_n6791.n813 w_4660_n6791.n812 27.1064
R16247 w_4660_n6791.n812 w_4660_n6791.n640 27.1064
R16248 w_4660_n6791.n806 w_4660_n6791.n640 27.1064
R16249 w_4660_n6791.n806 w_4660_n6791.n805 27.1064
R16250 w_4660_n6791.n805 w_4660_n6791.n804 27.1064
R16251 w_4660_n6791.n804 w_4660_n6791.n648 27.1064
R16252 w_4660_n6791.n798 w_4660_n6791.n648 27.1064
R16253 w_4660_n6791.n798 w_4660_n6791.n797 27.1064
R16254 w_4660_n6791.n797 w_4660_n6791.n796 27.1064
R16255 w_4660_n6791.n796 w_4660_n6791.n657 27.1064
R16256 w_4660_n6791.n790 w_4660_n6791.n657 27.1064
R16257 w_4660_n6791.n790 w_4660_n6791.n789 27.1064
R16258 w_4660_n6791.n789 w_4660_n6791.n667 27.1064
R16259 w_4660_n6791.n674 w_4660_n6791.n667 27.1064
R16260 w_4660_n6791.n783 w_4660_n6791.n674 27.1064
R16261 w_4660_n6791.n783 w_4660_n6791.n782 27.1064
R16262 w_4660_n6791.n782 w_4660_n6791.n781 27.1064
R16263 w_4660_n6791.n781 w_4660_n6791.n675 27.1064
R16264 w_4660_n6791.n775 w_4660_n6791.n675 27.1064
R16265 w_4660_n6791.n775 w_4660_n6791.n774 27.1064
R16266 w_4660_n6791.n774 w_4660_n6791.n773 27.1064
R16267 w_4660_n6791.n773 w_4660_n6791.n684 27.1064
R16268 w_4660_n6791.n933 w_4660_n6791.n507 27.1064
R16269 w_4660_n6791.n515 w_4660_n6791.n507 27.1064
R16270 w_4660_n6791.n926 w_4660_n6791.n515 27.1064
R16271 w_4660_n6791.n926 w_4660_n6791.n925 27.1064
R16272 w_4660_n6791.n925 w_4660_n6791.n924 27.1064
R16273 w_4660_n6791.n924 w_4660_n6791.n516 27.1064
R16274 w_4660_n6791.n918 w_4660_n6791.n516 27.1064
R16275 w_4660_n6791.n918 w_4660_n6791.n917 27.1064
R16276 w_4660_n6791.n917 w_4660_n6791.n916 27.1064
R16277 w_4660_n6791.n916 w_4660_n6791.n525 27.1064
R16278 w_4660_n6791.n910 w_4660_n6791.n525 27.1064
R16279 w_4660_n6791.n910 w_4660_n6791.n909 27.1064
R16280 w_4660_n6791.n909 w_4660_n6791.n908 27.1064
R16281 w_4660_n6791.n908 w_4660_n6791.n533 27.1064
R16282 w_4660_n6791.n902 w_4660_n6791.n533 27.1064
R16283 w_4660_n6791.n902 w_4660_n6791.n901 27.1064
R16284 w_4660_n6791.n901 w_4660_n6791.n541 27.1064
R16285 w_4660_n6791.n549 w_4660_n6791.n541 27.1064
R16286 w_4660_n6791.n895 w_4660_n6791.n549 27.1064
R16287 w_4660_n6791.n895 w_4660_n6791.n894 27.1064
R16288 w_4660_n6791.n894 w_4660_n6791.n550 27.1064
R16289 w_4660_n6791.n559 w_4660_n6791.n550 27.1064
R16290 w_4660_n6791.n887 w_4660_n6791.n559 27.1064
R16291 w_4660_n6791.n887 w_4660_n6791.n886 27.1064
R16292 w_4660_n6791.n886 w_4660_n6791.n885 27.1064
R16293 w_4660_n6791.n885 w_4660_n6791.n560 27.1064
R16294 w_4660_n6791.n879 w_4660_n6791.n560 27.1064
R16295 w_4660_n6791.n879 w_4660_n6791.n878 27.1064
R16296 w_4660_n6791.n878 w_4660_n6791.n877 27.1064
R16297 w_4660_n6791.n877 w_4660_n6791.n568 27.1064
R16298 w_4660_n6791.n871 w_4660_n6791.n568 27.1064
R16299 w_4660_n6791.n871 w_4660_n6791.n870 27.1064
R16300 w_4660_n6791.n870 w_4660_n6791.n869 27.1064
R16301 w_4660_n6791.n869 w_4660_n6791.n577 27.1064
R16302 w_4660_n6791.n863 w_4660_n6791.n577 27.1064
R16303 w_4660_n6791.n863 w_4660_n6791.n862 27.1064
R16304 w_4660_n6791.n862 w_4660_n6791.n587 27.1064
R16305 w_4660_n6791.n853 w_4660_n6791.n587 27.1064
R16306 w_4660_n6791.n855 w_4660_n6791.n853 27.1064
R16307 w_4660_n6791.n855 w_4660_n6791.n854 27.1064
R16308 w_4660_n6791.n850 w_4660_n6791.n849 27.1064
R16309 w_4660_n6791.n849 w_4660_n6791.n848 27.1064
R16310 w_4660_n6791.n848 w_4660_n6791.n600 27.1064
R16311 w_4660_n6791.n842 w_4660_n6791.n600 27.1064
R16312 w_4660_n6791.n842 w_4660_n6791.n841 27.1064
R16313 w_4660_n6791.n841 w_4660_n6791.n610 27.1064
R16314 w_4660_n6791.n619 w_4660_n6791.n610 27.1064
R16315 w_4660_n6791.n834 w_4660_n6791.n619 27.1064
R16316 w_4660_n6791.n834 w_4660_n6791.n833 27.1064
R16317 w_4660_n6791.n833 w_4660_n6791.n832 27.1064
R16318 w_4660_n6791.n832 w_4660_n6791.n19 27.1064
R16319 w_4660_n6791.n826 w_4660_n6791.n19 27.1064
R16320 w_4660_n6791.n826 w_4660_n6791.n825 27.1064
R16321 w_4660_n6791.n825 w_4660_n6791.n824 27.1064
R16322 w_4660_n6791.n824 w_4660_n6791.n626 27.1064
R16323 w_4660_n6791.n818 w_4660_n6791.n626 27.1064
R16324 w_4660_n6791.n818 w_4660_n6791.n817 27.1064
R16325 w_4660_n6791.n817 w_4660_n6791.n816 27.1064
R16326 w_4660_n6791.n816 w_4660_n6791.n634 27.1064
R16327 w_4660_n6791.n810 w_4660_n6791.n634 27.1064
R16328 w_4660_n6791.n810 w_4660_n6791.n809 27.1064
R16329 w_4660_n6791.n809 w_4660_n6791.n644 27.1064
R16330 w_4660_n6791.n652 w_4660_n6791.n644 27.1064
R16331 w_4660_n6791.n802 w_4660_n6791.n652 27.1064
R16332 w_4660_n6791.n802 w_4660_n6791.n801 27.1064
R16333 w_4660_n6791.n801 w_4660_n6791.n653 27.1064
R16334 w_4660_n6791.n662 w_4660_n6791.n653 27.1064
R16335 w_4660_n6791.n794 w_4660_n6791.n662 27.1064
R16336 w_4660_n6791.n794 w_4660_n6791.n793 27.1064
R16337 w_4660_n6791.n793 w_4660_n6791.n792 27.1064
R16338 w_4660_n6791.n792 w_4660_n6791.n663 27.1064
R16339 w_4660_n6791.n786 w_4660_n6791.n663 27.1064
R16340 w_4660_n6791.n786 w_4660_n6791.n785 27.1064
R16341 w_4660_n6791.n785 w_4660_n6791.n784 27.1064
R16342 w_4660_n6791.n784 w_4660_n6791.n670 27.1064
R16343 w_4660_n6791.n779 w_4660_n6791.n670 27.1064
R16344 w_4660_n6791.n779 w_4660_n6791.n778 27.1064
R16345 w_4660_n6791.n778 w_4660_n6791.n777 27.1064
R16346 w_4660_n6791.n777 w_4660_n6791.n679 27.1064
R16347 w_4660_n6791.n771 w_4660_n6791.n679 27.1064
R16348 w_4660_n6791.n771 w_4660_n6791.n770 27.1064
R16349 w_4660_n6791.n2292 w_4660_n6791.n2283 27.1064
R16350 w_4660_n6791.n2293 w_4660_n6791.n2292 27.1064
R16351 w_4660_n6791.n2295 w_4660_n6791.n2293 27.1064
R16352 w_4660_n6791.n2295 w_4660_n6791.n2294 27.1064
R16353 w_4660_n6791.n2294 w_4660_n6791.n421 27.1064
R16354 w_4660_n6791.n2302 w_4660_n6791.n421 27.1064
R16355 w_4660_n6791.n2303 w_4660_n6791.n2302 27.1064
R16356 w_4660_n6791.n2304 w_4660_n6791.n2303 27.1064
R16357 w_4660_n6791.n2304 w_4660_n6791.n418 27.1064
R16358 w_4660_n6791.n2310 w_4660_n6791.n418 27.1064
R16359 w_4660_n6791.n2311 w_4660_n6791.n2310 27.1064
R16360 w_4660_n6791.n2312 w_4660_n6791.n2311 27.1064
R16361 w_4660_n6791.n2312 w_4660_n6791.n413 27.1064
R16362 w_4660_n6791.n2319 w_4660_n6791.n413 27.1064
R16363 w_4660_n6791.n2320 w_4660_n6791.n2319 27.1064
R16364 w_4660_n6791.n2322 w_4660_n6791.n2320 27.1064
R16365 w_4660_n6791.n2322 w_4660_n6791.n2321 27.1064
R16366 w_4660_n6791.n2321 w_4660_n6791.n400 27.1064
R16367 w_4660_n6791.n2331 w_4660_n6791.n400 27.1064
R16368 w_4660_n6791.n2332 w_4660_n6791.n2331 27.1064
R16369 w_4660_n6791.n2333 w_4660_n6791.n2332 27.1064
R16370 w_4660_n6791.n2333 w_4660_n6791.n396 27.1064
R16371 w_4660_n6791.n2339 w_4660_n6791.n396 27.1064
R16372 w_4660_n6791.n2340 w_4660_n6791.n2339 27.1064
R16373 w_4660_n6791.n2341 w_4660_n6791.n2340 27.1064
R16374 w_4660_n6791.n2341 w_4660_n6791.n391 27.1064
R16375 w_4660_n6791.n2348 w_4660_n6791.n391 27.1064
R16376 w_4660_n6791.n2349 w_4660_n6791.n2348 27.1064
R16377 w_4660_n6791.n2351 w_4660_n6791.n2349 27.1064
R16378 w_4660_n6791.n2351 w_4660_n6791.n2350 27.1064
R16379 w_4660_n6791.n2350 w_4660_n6791.n378 27.1064
R16380 w_4660_n6791.n2360 w_4660_n6791.n378 27.1064
R16381 w_4660_n6791.n2361 w_4660_n6791.n2360 27.1064
R16382 w_4660_n6791.n2362 w_4660_n6791.n2361 27.1064
R16383 w_4660_n6791.n2362 w_4660_n6791.n374 27.1064
R16384 w_4660_n6791.n2368 w_4660_n6791.n374 27.1064
R16385 w_4660_n6791.n2369 w_4660_n6791.n2368 27.1064
R16386 w_4660_n6791.n2370 w_4660_n6791.n2369 27.1064
R16387 w_4660_n6791.n2370 w_4660_n6791.n369 27.1064
R16388 w_4660_n6791.n2376 w_4660_n6791.n369 27.1064
R16389 w_4660_n6791.n2379 w_4660_n6791.n2378 27.1064
R16390 w_4660_n6791.n2379 w_4660_n6791.n364 27.1064
R16391 w_4660_n6791.n2386 w_4660_n6791.n364 27.1064
R16392 w_4660_n6791.n2387 w_4660_n6791.n2386 27.1064
R16393 w_4660_n6791.n2388 w_4660_n6791.n2387 27.1064
R16394 w_4660_n6791.n2388 w_4660_n6791.n353 27.1064
R16395 w_4660_n6791.n2399 w_4660_n6791.n353 27.1064
R16396 w_4660_n6791.n2400 w_4660_n6791.n2399 27.1064
R16397 w_4660_n6791.n2401 w_4660_n6791.n2400 27.1064
R16398 w_4660_n6791.n2401 w_4660_n6791.n349 27.1064
R16399 w_4660_n6791.n2408 w_4660_n6791.n349 27.1064
R16400 w_4660_n6791.n2409 w_4660_n6791.n2408 27.1064
R16401 w_4660_n6791.n2410 w_4660_n6791.n2409 27.1064
R16402 w_4660_n6791.n2410 w_4660_n6791.n345 27.1064
R16403 w_4660_n6791.n2416 w_4660_n6791.n345 27.1064
R16404 w_4660_n6791.n2417 w_4660_n6791.n2416 27.1064
R16405 w_4660_n6791.n2418 w_4660_n6791.n2417 27.1064
R16406 w_4660_n6791.n2418 w_4660_n6791.n340 27.1064
R16407 w_4660_n6791.n2425 w_4660_n6791.n340 27.1064
R16408 w_4660_n6791.n2426 w_4660_n6791.n2425 27.1064
R16409 w_4660_n6791.n2428 w_4660_n6791.n2426 27.1064
R16410 w_4660_n6791.n2428 w_4660_n6791.n2427 27.1064
R16411 w_4660_n6791.n2427 w_4660_n6791.n327 27.1064
R16412 w_4660_n6791.n2435 w_4660_n6791.n327 27.1064
R16413 w_4660_n6791.n2436 w_4660_n6791.n2435 27.1064
R16414 w_4660_n6791.n2437 w_4660_n6791.n2436 27.1064
R16415 w_4660_n6791.n2437 w_4660_n6791.n324 27.1064
R16416 w_4660_n6791.n2443 w_4660_n6791.n324 27.1064
R16417 w_4660_n6791.n2444 w_4660_n6791.n2443 27.1064
R16418 w_4660_n6791.n2445 w_4660_n6791.n2444 27.1064
R16419 w_4660_n6791.n2445 w_4660_n6791.n319 27.1064
R16420 w_4660_n6791.n2452 w_4660_n6791.n319 27.1064
R16421 w_4660_n6791.n2453 w_4660_n6791.n2452 27.1064
R16422 w_4660_n6791.n2455 w_4660_n6791.n2453 27.1064
R16423 w_4660_n6791.n2455 w_4660_n6791.n2454 27.1064
R16424 w_4660_n6791.n2454 w_4660_n6791.n306 27.1064
R16425 w_4660_n6791.n2463 w_4660_n6791.n306 27.1064
R16426 w_4660_n6791.n2464 w_4660_n6791.n2463 27.1064
R16427 w_4660_n6791.n2465 w_4660_n6791.n2464 27.1064
R16428 w_4660_n6791.n2465 w_4660_n6791.n302 27.1064
R16429 w_4660_n6791.n2470 w_4660_n6791.n302 27.1064
R16430 w_4660_n6791.n2290 w_4660_n6791.n2288 27.1064
R16431 w_4660_n6791.n2290 w_4660_n6791.n2289 27.1064
R16432 w_4660_n6791.n2289 w_4660_n6791.n2279 27.1064
R16433 w_4660_n6791.n2281 w_4660_n6791.n2279 27.1064
R16434 w_4660_n6791.n2281 w_4660_n6791.n2280 27.1064
R16435 w_4660_n6791.n2280 w_4660_n6791.n424 27.1064
R16436 w_4660_n6791.n424 w_4660_n6791.n423 27.1064
R16437 w_4660_n6791.n423 w_4660_n6791.n420 27.1064
R16438 w_4660_n6791.n2307 w_4660_n6791.n420 27.1064
R16439 w_4660_n6791.n2308 w_4660_n6791.n2307 27.1064
R16440 w_4660_n6791.n2308 w_4660_n6791.n415 27.1064
R16441 w_4660_n6791.n2314 w_4660_n6791.n415 27.1064
R16442 w_4660_n6791.n2315 w_4660_n6791.n2314 27.1064
R16443 w_4660_n6791.n2317 w_4660_n6791.n2315 27.1064
R16444 w_4660_n6791.n2317 w_4660_n6791.n2316 27.1064
R16445 w_4660_n6791.n2316 w_4660_n6791.n409 27.1064
R16446 w_4660_n6791.n411 w_4660_n6791.n409 27.1064
R16447 w_4660_n6791.n411 w_4660_n6791.n410 27.1064
R16448 w_4660_n6791.n410 w_4660_n6791.n403 27.1064
R16449 w_4660_n6791.n403 w_4660_n6791.n402 27.1064
R16450 w_4660_n6791.n402 w_4660_n6791.n398 27.1064
R16451 w_4660_n6791.n2336 w_4660_n6791.n398 27.1064
R16452 w_4660_n6791.n2337 w_4660_n6791.n2336 27.1064
R16453 w_4660_n6791.n2337 w_4660_n6791.n393 27.1064
R16454 w_4660_n6791.n2343 w_4660_n6791.n393 27.1064
R16455 w_4660_n6791.n2344 w_4660_n6791.n2343 27.1064
R16456 w_4660_n6791.n2346 w_4660_n6791.n2344 27.1064
R16457 w_4660_n6791.n2346 w_4660_n6791.n2345 27.1064
R16458 w_4660_n6791.n2345 w_4660_n6791.n387 27.1064
R16459 w_4660_n6791.n389 w_4660_n6791.n387 27.1064
R16460 w_4660_n6791.n389 w_4660_n6791.n388 27.1064
R16461 w_4660_n6791.n388 w_4660_n6791.n381 27.1064
R16462 w_4660_n6791.n381 w_4660_n6791.n380 27.1064
R16463 w_4660_n6791.n380 w_4660_n6791.n376 27.1064
R16464 w_4660_n6791.n2365 w_4660_n6791.n376 27.1064
R16465 w_4660_n6791.n2366 w_4660_n6791.n2365 27.1064
R16466 w_4660_n6791.n2366 w_4660_n6791.n371 27.1064
R16467 w_4660_n6791.n2372 w_4660_n6791.n371 27.1064
R16468 w_4660_n6791.n2373 w_4660_n6791.n2372 27.1064
R16469 w_4660_n6791.n2374 w_4660_n6791.n2373 27.1064
R16470 w_4660_n6791.n2381 w_4660_n6791.n366 27.1064
R16471 w_4660_n6791.n2382 w_4660_n6791.n2381 27.1064
R16472 w_4660_n6791.n2384 w_4660_n6791.n2382 27.1064
R16473 w_4660_n6791.n2384 w_4660_n6791.n2383 27.1064
R16474 w_4660_n6791.n2383 w_4660_n6791.n363 27.1064
R16475 w_4660_n6791.n363 w_4660_n6791.n362 27.1064
R16476 w_4660_n6791.n362 w_4660_n6791.n356 27.1064
R16477 w_4660_n6791.n356 w_4660_n6791.n355 27.1064
R16478 w_4660_n6791.n355 w_4660_n6791.n351 27.1064
R16479 w_4660_n6791.n2404 w_4660_n6791.n351 27.1064
R16480 w_4660_n6791.n2406 w_4660_n6791.n2404 27.1064
R16481 w_4660_n6791.n2406 w_4660_n6791.n2405 27.1064
R16482 w_4660_n6791.n2405 w_4660_n6791.n347 27.1064
R16483 w_4660_n6791.n2413 w_4660_n6791.n347 27.1064
R16484 w_4660_n6791.n2414 w_4660_n6791.n2413 27.1064
R16485 w_4660_n6791.n2414 w_4660_n6791.n342 27.1064
R16486 w_4660_n6791.n2420 w_4660_n6791.n342 27.1064
R16487 w_4660_n6791.n2421 w_4660_n6791.n2420 27.1064
R16488 w_4660_n6791.n2423 w_4660_n6791.n2421 27.1064
R16489 w_4660_n6791.n2423 w_4660_n6791.n2422 27.1064
R16490 w_4660_n6791.n2422 w_4660_n6791.n336 27.1064
R16491 w_4660_n6791.n338 w_4660_n6791.n336 27.1064
R16492 w_4660_n6791.n338 w_4660_n6791.n337 27.1064
R16493 w_4660_n6791.n337 w_4660_n6791.n330 27.1064
R16494 w_4660_n6791.n330 w_4660_n6791.n329 27.1064
R16495 w_4660_n6791.n329 w_4660_n6791.n326 27.1064
R16496 w_4660_n6791.n2440 w_4660_n6791.n326 27.1064
R16497 w_4660_n6791.n2441 w_4660_n6791.n2440 27.1064
R16498 w_4660_n6791.n2441 w_4660_n6791.n321 27.1064
R16499 w_4660_n6791.n2447 w_4660_n6791.n321 27.1064
R16500 w_4660_n6791.n2448 w_4660_n6791.n2447 27.1064
R16501 w_4660_n6791.n2450 w_4660_n6791.n2448 27.1064
R16502 w_4660_n6791.n2450 w_4660_n6791.n2449 27.1064
R16503 w_4660_n6791.n2449 w_4660_n6791.n315 27.1064
R16504 w_4660_n6791.n317 w_4660_n6791.n315 27.1064
R16505 w_4660_n6791.n317 w_4660_n6791.n316 27.1064
R16506 w_4660_n6791.n316 w_4660_n6791.n309 27.1064
R16507 w_4660_n6791.n309 w_4660_n6791.n308 27.1064
R16508 w_4660_n6791.n308 w_4660_n6791.n304 27.1064
R16509 w_4660_n6791.n2468 w_4660_n6791.n304 27.1064
R16510 w_4660_n6791.n1525 w_4660_n6791.n1522 27.1064
R16511 w_4660_n6791.n1529 w_4660_n6791.n1525 27.1064
R16512 w_4660_n6791.n1530 w_4660_n6791.n1529 27.1064
R16513 w_4660_n6791.n1533 w_4660_n6791.n1530 27.1064
R16514 w_4660_n6791.n1534 w_4660_n6791.n1533 27.1064
R16515 w_4660_n6791.n1536 w_4660_n6791.n1534 27.1064
R16516 w_4660_n6791.n1537 w_4660_n6791.n1536 27.1064
R16517 w_4660_n6791.n1540 w_4660_n6791.n1537 27.1064
R16518 w_4660_n6791.n1541 w_4660_n6791.n1540 27.1064
R16519 w_4660_n6791.n1544 w_4660_n6791.n1541 27.1064
R16520 w_4660_n6791.n1545 w_4660_n6791.n1544 27.1064
R16521 w_4660_n6791.n1549 w_4660_n6791.n1545 27.1064
R16522 w_4660_n6791.n1550 w_4660_n6791.n1549 27.1064
R16523 w_4660_n6791.n1554 w_4660_n6791.n1550 27.1064
R16524 w_4660_n6791.n1555 w_4660_n6791.n1554 27.1064
R16525 w_4660_n6791.n1558 w_4660_n6791.n1555 27.1064
R16526 w_4660_n6791.n1559 w_4660_n6791.n1558 27.1064
R16527 w_4660_n6791.n1562 w_4660_n6791.n1559 27.1064
R16528 w_4660_n6791.n1563 w_4660_n6791.n1562 27.1064
R16529 w_4660_n6791.n1567 w_4660_n6791.n1563 27.1064
R16530 w_4660_n6791.n1568 w_4660_n6791.n1567 27.1064
R16531 w_4660_n6791.n1572 w_4660_n6791.n1568 27.1064
R16532 w_4660_n6791.n1573 w_4660_n6791.n1572 27.1064
R16533 w_4660_n6791.n1577 w_4660_n6791.n1573 27.1064
R16534 w_4660_n6791.n1578 w_4660_n6791.n1577 27.1064
R16535 w_4660_n6791.n1581 w_4660_n6791.n1578 27.1064
R16536 w_4660_n6791.n1582 w_4660_n6791.n1581 27.1064
R16537 w_4660_n6791.n1584 w_4660_n6791.n1582 27.1064
R16538 w_4660_n6791.n1585 w_4660_n6791.n1584 27.1064
R16539 w_4660_n6791.n1589 w_4660_n6791.n1585 27.1064
R16540 w_4660_n6791.n1590 w_4660_n6791.n1589 27.1064
R16541 w_4660_n6791.n1594 w_4660_n6791.n1590 27.1064
R16542 w_4660_n6791.n1595 w_4660_n6791.n1594 27.1064
R16543 w_4660_n6791.n1598 w_4660_n6791.n1595 27.1064
R16544 w_4660_n6791.n1599 w_4660_n6791.n1598 27.1064
R16545 w_4660_n6791.n1602 w_4660_n6791.n1599 27.1064
R16546 w_4660_n6791.n1603 w_4660_n6791.n1602 27.1064
R16547 w_4660_n6791.n1674 w_4660_n6791.n1603 27.1064
R16548 w_4660_n6791.n1675 w_4660_n6791.n1674 27.1064
R16549 w_4660_n6791.n1675 w_4660_n6791.n234 27.1064
R16550 w_4660_n6791.n2525 w_4660_n6791.n2524 27.1064
R16551 w_4660_n6791.n2525 w_4660_n6791.n231 27.1064
R16552 w_4660_n6791.n231 w_4660_n6791.n230 27.1064
R16553 w_4660_n6791.n230 w_4660_n6791.n222 27.1064
R16554 w_4660_n6791.n2537 w_4660_n6791.n222 27.1064
R16555 w_4660_n6791.n2538 w_4660_n6791.n2537 27.1064
R16556 w_4660_n6791.n2539 w_4660_n6791.n2538 27.1064
R16557 w_4660_n6791.n2539 w_4660_n6791.n219 27.1064
R16558 w_4660_n6791.n219 w_4660_n6791.n218 27.1064
R16559 w_4660_n6791.n218 w_4660_n6791.n214 27.1064
R16560 w_4660_n6791.n214 w_4660_n6791.n213 27.1064
R16561 w_4660_n6791.n213 w_4660_n6791.n210 27.1064
R16562 w_4660_n6791.n210 w_4660_n6791.n209 27.1064
R16563 w_4660_n6791.n209 w_4660_n6791.n201 27.1064
R16564 w_4660_n6791.n2559 w_4660_n6791.n201 27.1064
R16565 w_4660_n6791.n2560 w_4660_n6791.n2559 27.1064
R16566 w_4660_n6791.n2561 w_4660_n6791.n2560 27.1064
R16567 w_4660_n6791.n2561 w_4660_n6791.n198 27.1064
R16568 w_4660_n6791.n198 w_4660_n6791.n197 27.1064
R16569 w_4660_n6791.n197 w_4660_n6791.n193 27.1064
R16570 w_4660_n6791.n193 w_4660_n6791.n192 27.1064
R16571 w_4660_n6791.n192 w_4660_n6791.n189 27.1064
R16572 w_4660_n6791.n189 w_4660_n6791.n188 27.1064
R16573 w_4660_n6791.n188 w_4660_n6791.n27 27.1064
R16574 w_4660_n6791.n2580 w_4660_n6791.n27 27.1064
R16575 w_4660_n6791.n2581 w_4660_n6791.n2580 27.1064
R16576 w_4660_n6791.n2582 w_4660_n6791.n2581 27.1064
R16577 w_4660_n6791.n2582 w_4660_n6791.n179 27.1064
R16578 w_4660_n6791.n179 w_4660_n6791.n178 27.1064
R16579 w_4660_n6791.n178 w_4660_n6791.n170 27.1064
R16580 w_4660_n6791.n2594 w_4660_n6791.n170 27.1064
R16581 w_4660_n6791.n2595 w_4660_n6791.n2594 27.1064
R16582 w_4660_n6791.n2596 w_4660_n6791.n2595 27.1064
R16583 w_4660_n6791.n2596 w_4660_n6791.n167 27.1064
R16584 w_4660_n6791.n167 w_4660_n6791.n166 27.1064
R16585 w_4660_n6791.n166 w_4660_n6791.n163 27.1064
R16586 w_4660_n6791.n163 w_4660_n6791.n162 27.1064
R16587 w_4660_n6791.n162 w_4660_n6791.n154 27.1064
R16588 w_4660_n6791.n156 w_4660_n6791.n154 27.1064
R16589 w_4660_n6791.n156 w_4660_n6791.n155 27.1064
R16590 w_4660_n6791.n155 w_4660_n6791.n144 27.1064
R16591 w_4660_n6791.n1757 w_4660_n6791.n1524 27.1064
R16592 w_4660_n6791.n1532 w_4660_n6791.n1524 27.1064
R16593 w_4660_n6791.n1750 w_4660_n6791.n1532 27.1064
R16594 w_4660_n6791.n1750 w_4660_n6791.n1749 27.1064
R16595 w_4660_n6791.n1749 w_4660_n6791.n1748 27.1064
R16596 w_4660_n6791.n1748 w_4660_n6791.n23 27.1064
R16597 w_4660_n6791.n1742 w_4660_n6791.n23 27.1064
R16598 w_4660_n6791.n1742 w_4660_n6791.n1741 27.1064
R16599 w_4660_n6791.n1741 w_4660_n6791.n1740 27.1064
R16600 w_4660_n6791.n1740 w_4660_n6791.n1539 27.1064
R16601 w_4660_n6791.n1734 w_4660_n6791.n1539 27.1064
R16602 w_4660_n6791.n1734 w_4660_n6791.n1733 27.1064
R16603 w_4660_n6791.n1733 w_4660_n6791.n1732 27.1064
R16604 w_4660_n6791.n1732 w_4660_n6791.n1547 27.1064
R16605 w_4660_n6791.n1726 w_4660_n6791.n1547 27.1064
R16606 w_4660_n6791.n1726 w_4660_n6791.n1725 27.1064
R16607 w_4660_n6791.n1725 w_4660_n6791.n1557 27.1064
R16608 w_4660_n6791.n1565 w_4660_n6791.n1557 27.1064
R16609 w_4660_n6791.n1718 w_4660_n6791.n1565 27.1064
R16610 w_4660_n6791.n1718 w_4660_n6791.n1717 27.1064
R16611 w_4660_n6791.n1717 w_4660_n6791.n1566 27.1064
R16612 w_4660_n6791.n1575 w_4660_n6791.n1566 27.1064
R16613 w_4660_n6791.n1710 w_4660_n6791.n1575 27.1064
R16614 w_4660_n6791.n1710 w_4660_n6791.n1709 27.1064
R16615 w_4660_n6791.n1709 w_4660_n6791.n1708 27.1064
R16616 w_4660_n6791.n1708 w_4660_n6791.n1576 27.1064
R16617 w_4660_n6791.n1702 w_4660_n6791.n1576 27.1064
R16618 w_4660_n6791.n1702 w_4660_n6791.n1701 27.1064
R16619 w_4660_n6791.n1701 w_4660_n6791.n1700 27.1064
R16620 w_4660_n6791.n1700 w_4660_n6791.n1583 27.1064
R16621 w_4660_n6791.n1695 w_4660_n6791.n1583 27.1064
R16622 w_4660_n6791.n1695 w_4660_n6791.n1694 27.1064
R16623 w_4660_n6791.n1694 w_4660_n6791.n1693 27.1064
R16624 w_4660_n6791.n1693 w_4660_n6791.n1592 27.1064
R16625 w_4660_n6791.n1687 w_4660_n6791.n1592 27.1064
R16626 w_4660_n6791.n1687 w_4660_n6791.n1686 27.1064
R16627 w_4660_n6791.n1686 w_4660_n6791.n1601 27.1064
R16628 w_4660_n6791.n1677 w_4660_n6791.n1601 27.1064
R16629 w_4660_n6791.n1679 w_4660_n6791.n1677 27.1064
R16630 w_4660_n6791.n1679 w_4660_n6791.n1678 27.1064
R16631 w_4660_n6791.n242 w_4660_n6791.n228 27.1064
R16632 w_4660_n6791.n2530 w_4660_n6791.n228 27.1064
R16633 w_4660_n6791.n2531 w_4660_n6791.n2530 27.1064
R16634 w_4660_n6791.n2532 w_4660_n6791.n2531 27.1064
R16635 w_4660_n6791.n2532 w_4660_n6791.n225 27.1064
R16636 w_4660_n6791.n225 w_4660_n6791.n224 27.1064
R16637 w_4660_n6791.n224 w_4660_n6791.n216 27.1064
R16638 w_4660_n6791.n2544 w_4660_n6791.n216 27.1064
R16639 w_4660_n6791.n2545 w_4660_n6791.n2544 27.1064
R16640 w_4660_n6791.n2546 w_4660_n6791.n2545 27.1064
R16641 w_4660_n6791.n2546 w_4660_n6791.n207 27.1064
R16642 w_4660_n6791.n2552 w_4660_n6791.n207 27.1064
R16643 w_4660_n6791.n2553 w_4660_n6791.n2552 27.1064
R16644 w_4660_n6791.n2554 w_4660_n6791.n2553 27.1064
R16645 w_4660_n6791.n2554 w_4660_n6791.n204 27.1064
R16646 w_4660_n6791.n204 w_4660_n6791.n203 27.1064
R16647 w_4660_n6791.n203 w_4660_n6791.n195 27.1064
R16648 w_4660_n6791.n2566 w_4660_n6791.n195 27.1064
R16649 w_4660_n6791.n2567 w_4660_n6791.n2566 27.1064
R16650 w_4660_n6791.n2568 w_4660_n6791.n2567 27.1064
R16651 w_4660_n6791.n2568 w_4660_n6791.n186 27.1064
R16652 w_4660_n6791.n2574 w_4660_n6791.n186 27.1064
R16653 w_4660_n6791.n2575 w_4660_n6791.n2574 27.1064
R16654 w_4660_n6791.n2576 w_4660_n6791.n2575 27.1064
R16655 w_4660_n6791.n2576 w_4660_n6791.n183 27.1064
R16656 w_4660_n6791.n183 w_4660_n6791.n182 27.1064
R16657 w_4660_n6791.n182 w_4660_n6791.n176 27.1064
R16658 w_4660_n6791.n2587 w_4660_n6791.n176 27.1064
R16659 w_4660_n6791.n2588 w_4660_n6791.n2587 27.1064
R16660 w_4660_n6791.n2589 w_4660_n6791.n2588 27.1064
R16661 w_4660_n6791.n2589 w_4660_n6791.n173 27.1064
R16662 w_4660_n6791.n173 w_4660_n6791.n172 27.1064
R16663 w_4660_n6791.n172 w_4660_n6791.n164 27.1064
R16664 w_4660_n6791.n2601 w_4660_n6791.n164 27.1064
R16665 w_4660_n6791.n2602 w_4660_n6791.n2601 27.1064
R16666 w_4660_n6791.n2604 w_4660_n6791.n2602 27.1064
R16667 w_4660_n6791.n2604 w_4660_n6791.n2603 27.1064
R16668 w_4660_n6791.n2603 w_4660_n6791.n159 27.1064
R16669 w_4660_n6791.n159 w_4660_n6791.n158 27.1064
R16670 w_4660_n6791.n158 w_4660_n6791.n146 27.1064
R16671 w_4660_n6791.n2617 w_4660_n6791.n146 27.1064
R16672 w_4660_n6791.n2675 w_4660_n6791.n84 26.3319
R16673 w_4660_n6791.n92 w_4660_n6791.n84 26.3319
R16674 w_4660_n6791.n2668 w_4660_n6791.n92 26.3319
R16675 w_4660_n6791.n2668 w_4660_n6791.n2667 26.3319
R16676 w_4660_n6791.n2667 w_4660_n6791.n2666 26.3319
R16677 w_4660_n6791.n2666 w_4660_n6791.n93 26.3319
R16678 w_4660_n6791.n2660 w_4660_n6791.n93 26.3319
R16679 w_4660_n6791.n2660 w_4660_n6791.n2659 26.3319
R16680 w_4660_n6791.n2659 w_4660_n6791.n2658 26.3319
R16681 w_4660_n6791.n2658 w_4660_n6791.n101 26.3319
R16682 w_4660_n6791.n2652 w_4660_n6791.n101 26.3319
R16683 w_4660_n6791.n966 w_4660_n6791.n109 26.3319
R16684 w_4660_n6791.n967 w_4660_n6791.n966 26.3319
R16685 w_4660_n6791.n968 w_4660_n6791.n967 26.3319
R16686 w_4660_n6791.n968 w_4660_n6791.n953 26.3319
R16687 w_4660_n6791.n974 w_4660_n6791.n953 26.3319
R16688 w_4660_n6791.n975 w_4660_n6791.n974 26.3319
R16689 w_4660_n6791.n976 w_4660_n6791.n975 26.3319
R16690 w_4660_n6791.n976 w_4660_n6791.n946 26.3319
R16691 w_4660_n6791.n983 w_4660_n6791.n946 26.3319
R16692 w_4660_n6791.n984 w_4660_n6791.n983 26.3319
R16693 w_4660_n6791.n1414 w_4660_n6791.n984 26.3319
R16694 w_4660_n6791.n1423 w_4660_n6791.n1422 26.3319
R16695 w_4660_n6791.n1423 w_4660_n6791.n496 26.3319
R16696 w_4660_n6791.n1429 w_4660_n6791.n496 26.3319
R16697 w_4660_n6791.n1430 w_4660_n6791.n1429 26.3319
R16698 w_4660_n6791.n1431 w_4660_n6791.n1430 26.3319
R16699 w_4660_n6791.n1431 w_4660_n6791.n488 26.3319
R16700 w_4660_n6791.n1437 w_4660_n6791.n488 26.3319
R16701 w_4660_n6791.n1438 w_4660_n6791.n1437 26.3319
R16702 w_4660_n6791.n1439 w_4660_n6791.n1438 26.3319
R16703 w_4660_n6791.n1439 w_4660_n6791.n480 26.3319
R16704 w_4660_n6791.n1445 w_4660_n6791.n480 26.3319
R16705 w_4660_n6791.n1446 w_4660_n6791.n1445 26.3319
R16706 w_4660_n6791.n1448 w_4660_n6791.n472 26.3319
R16707 w_4660_n6791.n1454 w_4660_n6791.n472 26.3319
R16708 w_4660_n6791.n1455 w_4660_n6791.n1454 26.3319
R16709 w_4660_n6791.n1456 w_4660_n6791.n1455 26.3319
R16710 w_4660_n6791.n1456 w_4660_n6791.n465 26.3319
R16711 w_4660_n6791.n1463 w_4660_n6791.n465 26.3319
R16712 w_4660_n6791.n1464 w_4660_n6791.n1463 26.3319
R16713 w_4660_n6791.n1466 w_4660_n6791.n1464 26.3319
R16714 w_4660_n6791.n1466 w_4660_n6791.n1465 26.3319
R16715 w_4660_n6791.n1465 w_4660_n6791.n461 26.3319
R16716 w_4660_n6791.n765 w_4660_n6791.n461 26.3319
R16717 w_4660_n6791.n1518 w_4660_n6791.n454 26.3319
R16718 w_4660_n6791.n1512 w_4660_n6791.n454 26.3319
R16719 w_4660_n6791.n1512 w_4660_n6791.n1511 26.3319
R16720 w_4660_n6791.n1511 w_4660_n6791.n1510 26.3319
R16721 w_4660_n6791.n1510 w_4660_n6791.n1481 26.3319
R16722 w_4660_n6791.n1504 w_4660_n6791.n1481 26.3319
R16723 w_4660_n6791.n1504 w_4660_n6791.n1503 26.3319
R16724 w_4660_n6791.n1503 w_4660_n6791.n1502 26.3319
R16725 w_4660_n6791.n1502 w_4660_n6791.n1489 26.3319
R16726 w_4660_n6791.n1496 w_4660_n6791.n1489 26.3319
R16727 w_4660_n6791.n1496 w_4660_n6791.n116 26.3319
R16728 w_4660_n6791.n2646 w_4660_n6791.n117 26.3319
R16729 w_4660_n6791.n2640 w_4660_n6791.n117 26.3319
R16730 w_4660_n6791.n2640 w_4660_n6791.n2639 26.3319
R16731 w_4660_n6791.n2639 w_4660_n6791.n2638 26.3319
R16732 w_4660_n6791.n2638 w_4660_n6791.n126 26.3319
R16733 w_4660_n6791.n2632 w_4660_n6791.n126 26.3319
R16734 w_4660_n6791.n2632 w_4660_n6791.n2631 26.3319
R16735 w_4660_n6791.n2631 w_4660_n6791.n2630 26.3319
R16736 w_4660_n6791.n2630 w_4660_n6791.n134 26.3319
R16737 w_4660_n6791.n2624 w_4660_n6791.n134 26.3319
R16738 w_4660_n6791.n2624 w_4660_n6791.n2623 26.3319
R16739 w_4660_n6791.n2518 w_4660_n6791.n248 26.3319
R16740 w_4660_n6791.n2512 w_4660_n6791.n248 26.3319
R16741 w_4660_n6791.n2512 w_4660_n6791.n2511 26.3319
R16742 w_4660_n6791.n2511 w_4660_n6791.n2510 26.3319
R16743 w_4660_n6791.n2510 w_4660_n6791.n262 26.3319
R16744 w_4660_n6791.n2504 w_4660_n6791.n262 26.3319
R16745 w_4660_n6791.n2504 w_4660_n6791.n2503 26.3319
R16746 w_4660_n6791.n2503 w_4660_n6791.n2502 26.3319
R16747 w_4660_n6791.n2502 w_4660_n6791.n270 26.3319
R16748 w_4660_n6791.n2496 w_4660_n6791.n270 26.3319
R16749 w_4660_n6791.n2496 w_4660_n6791.n2495 26.3319
R16750 w_4660_n6791.n2495 w_4660_n6791.n2494 26.3319
R16751 w_4660_n6791.n2488 w_4660_n6791.n286 26.3319
R16752 w_4660_n6791.n2488 w_4660_n6791.n2487 26.3319
R16753 w_4660_n6791.n2487 w_4660_n6791.n2486 26.3319
R16754 w_4660_n6791.n2486 w_4660_n6791.n287 26.3319
R16755 w_4660_n6791.n2480 w_4660_n6791.n287 26.3319
R16756 w_4660_n6791.n2480 w_4660_n6791.n2479 26.3319
R16757 w_4660_n6791.n2479 w_4660_n6791.n2478 26.3319
R16758 w_4660_n6791.n2478 w_4660_n6791.n295 26.3319
R16759 w_4660_n6791.n2472 w_4660_n6791.n295 26.3319
R16760 w_4660_n6791.n2472 w_4660_n6791.n2471 26.3319
R16761 w_4660_n6791.n990 w_4660_n6791.n985 25.4499
R16762 w_4660_n6791.n1414 w_4660_n6791.n1413 25.2348
R16763 w_4660_n6791.n761 w_4660_n6791.n453 24.0946
R16764 w_4660_n6791.n2623 w_4660_n6791.n2622 23.7719
R16765 w_4660_n6791.n286 w_4660_n6791.n278 23.7719
R16766 w_4660_n6791.n764 w_4660_n6791.n762 23.7181
R16767 w_4660_n6791.n1413 w_4660_n6791.n1412 23.7181
R16768 w_4660_n6791.n1421 w_4660_n6791.n1420 23.5353
R16769 w_4660_n6791.n1448 w_4660_n6791.n1447 22.3091
R16770 w_4660_n6791.n2519 w_4660_n6791.n145 22.0294
R16771 w_4660_n6791.n2622 w_4660_n6791.n142 20.7064
R16772 w_4660_n6791.n2676 w_4660_n6791.n61 20.7064
R16773 w_4660_n6791.n83 w_4660_n6791.n65 20.3299
R16774 w_4660_n6791.n1762 w_4660_n6791.t122 19.6596
R16775 w_4660_n6791.n2649 w_4660_n6791.t77 19.6596
R16776 w_4660_n6791.n72 w_4660_n6791.n65 19.577
R16777 w_4660_n6791.n2652 w_4660_n6791.n2651 17.9205
R16778 w_4660_n6791.n2620 w_4660_n6791.n2619 17.3181
R16779 w_4660_n6791.n1519 w_4660_n6791.n1518 17.1891
R16780 w_4660_n6791.n2647 w_4660_n6791.n116 16.4576
R16781 w_4660_n6791.n2677 w_4660_n6791.n83 15.8123
R16782 w_4660_n6791.n2676 w_4660_n6791.n2675 15.7262
R16783 w_4660_n6791.n764 w_4660_n6791.n763 15.2529
R16784 w_4660_n6791.n1605 w_4660_n6791.n232 15.0593
R16785 w_4660_n6791.n596 w_4660_n6791.n595 15.0593
R16786 w_4660_n6791.n1855 w_4660_n6791.n235 15.0593
R16787 w_4660_n6791.n2184 w_4660_n6791.n2183 15.0593
R16788 w_4660_n6791.n1314 w_4660_n6791.n1313 15.0593
R16789 w_4660_n6791.n1069 w_4660_n6791.n236 15.0593
R16790 w_4660_n6791.n1309 w_4660_n6791.n237 15.0593
R16791 w_4660_n6791.n591 w_4660_n6791.n240 15.0593
R16792 w_4660_n6791.n854 w_4660_n6791.n241 15.0593
R16793 w_4660_n6791.n2378 w_4660_n6791.n2377 15.0593
R16794 w_4660_n6791.n366 w_4660_n6791.n245 15.0593
R16795 w_4660_n6791.n2524 w_4660_n6791.n2523 15.0593
R16796 w_4660_n6791.n243 w_4660_n6791.n242 15.0593
R16797 w_4660_n6791.t122 w_4660_n6791.t17 13.4096
R16798 w_4660_n6791.t17 w_4660_n6791.t291 13.4096
R16799 w_4660_n6791.t291 w_4660_n6791.t25 13.4096
R16800 w_4660_n6791.t25 w_4660_n6791.t166 13.4096
R16801 w_4660_n6791.t166 w_4660_n6791.t240 13.4096
R16802 w_4660_n6791.t240 w_4660_n6791.t144 13.4096
R16803 w_4660_n6791.t144 w_4660_n6791.t118 13.4096
R16804 w_4660_n6791.t118 w_4660_n6791.t60 13.4096
R16805 w_4660_n6791.t60 w_4660_n6791.t107 13.4096
R16806 w_4660_n6791.t107 w_4660_n6791.t94 13.4096
R16807 w_4660_n6791.t94 w_4660_n6791.t7 13.4096
R16808 w_4660_n6791.t7 w_4660_n6791.t33 13.4096
R16809 w_4660_n6791.t33 w_4660_n6791.t2 13.4096
R16810 w_4660_n6791.t2 w_4660_n6791.t70 13.4096
R16811 w_4660_n6791.t70 w_4660_n6791.t47 13.4096
R16812 w_4660_n6791.t47 w_4660_n6791.t30 13.4096
R16813 w_4660_n6791.t30 w_4660_n6791.t62 13.4096
R16814 w_4660_n6791.t62 w_4660_n6791.t102 13.4096
R16815 w_4660_n6791.t102 w_4660_n6791.t86 13.4096
R16816 w_4660_n6791.t86 w_4660_n6791.t37 13.4096
R16817 w_4660_n6791.t37 w_4660_n6791.t67 13.4096
R16818 w_4660_n6791.t67 w_4660_n6791.t88 13.4096
R16819 w_4660_n6791.t88 w_4660_n6791.t83 13.4096
R16820 w_4660_n6791.t83 w_4660_n6791.t79 13.4096
R16821 w_4660_n6791.t43 w_4660_n6791.t163 13.4096
R16822 w_4660_n6791.t163 w_4660_n6791.t11 13.4096
R16823 w_4660_n6791.t11 w_4660_n6791.t112 13.4096
R16824 w_4660_n6791.t112 w_4660_n6791.t168 13.4096
R16825 w_4660_n6791.t168 w_4660_n6791.t50 13.4096
R16826 w_4660_n6791.t50 w_4660_n6791.t0 13.4096
R16827 w_4660_n6791.t0 w_4660_n6791.t35 13.4096
R16828 w_4660_n6791.t35 w_4660_n6791.t72 13.4096
R16829 w_4660_n6791.t72 w_4660_n6791.t98 13.4096
R16830 w_4660_n6791.t98 w_4660_n6791.t15 13.4096
R16831 w_4660_n6791.t15 w_4660_n6791.t141 13.4096
R16832 w_4660_n6791.t141 w_4660_n6791.t41 13.4096
R16833 w_4660_n6791.t41 w_4660_n6791.t52 13.4096
R16834 w_4660_n6791.t52 w_4660_n6791.t23 13.4096
R16835 w_4660_n6791.t23 w_4660_n6791.t64 13.4096
R16836 w_4660_n6791.t64 w_4660_n6791.t5 13.4096
R16837 w_4660_n6791.t5 w_4660_n6791.t39 13.4096
R16838 w_4660_n6791.t39 w_4660_n6791.t45 13.4096
R16839 w_4660_n6791.t45 w_4660_n6791.t130 13.4096
R16840 w_4660_n6791.t130 w_4660_n6791.t13 13.4096
R16841 w_4660_n6791.t13 w_4660_n6791.t92 13.4096
R16842 w_4660_n6791.t92 w_4660_n6791.t109 13.4096
R16843 w_4660_n6791.t109 w_4660_n6791.t148 13.4096
R16844 w_4660_n6791.t148 w_4660_n6791.t77 13.4096
R16845 w_4660_n6791.n1606 w_4660_n6791.n1605 12.0476
R16846 w_4660_n6791.n597 w_4660_n6791.n596 12.0476
R16847 w_4660_n6791.n1852 w_4660_n6791.n235 12.0476
R16848 w_4660_n6791.n2185 w_4660_n6791.n2184 12.0476
R16849 w_4660_n6791.n1315 w_4660_n6791.n1314 12.0476
R16850 w_4660_n6791.n1317 w_4660_n6791.n236 12.0476
R16851 w_4660_n6791.n1065 w_4660_n6791.n237 12.0476
R16852 w_4660_n6791.n599 w_4660_n6791.n240 12.0476
R16853 w_4660_n6791.n850 w_4660_n6791.n241 12.0476
R16854 w_4660_n6791.n2377 w_4660_n6791.n2376 12.0476
R16855 w_4660_n6791.n2374 w_4660_n6791.n245 12.0476
R16856 w_4660_n6791.n2523 w_4660_n6791.n234 12.0476
R16857 w_4660_n6791.n1678 w_4660_n6791.n243 12.0476
R16858 w_4660_n6791.n765 w_4660_n6791.n764 11.3376
R16859 w_4660_n6791.n766 w_4660_n6791.n763 11.2946
R16860 w_4660_n6791.n2618 w_4660_n6791.n145 11.2946
R16861 w_4660_n6791.n2677 w_4660_n6791.n2676 10.7353
R16862 w_4660_n6791.n2647 w_4660_n6791.n2646 9.87479
R16863 w_4660_n6791.n1420 w_4660_n6791.n938 9.78874
R16864 w_4660_n6791.n45 w_4660_n6791.t274 9.52217
R16865 w_4660_n6791.n45 w_4660_n6791.t248 9.52217
R16866 w_4660_n6791.n1921 w_4660_n6791.t341 9.52217
R16867 w_4660_n6791.n1921 w_4660_n6791.t312 9.52217
R16868 w_4660_n6791.n1924 w_4660_n6791.t353 9.52217
R16869 w_4660_n6791.n1924 w_4660_n6791.t380 9.52217
R16870 w_4660_n6791.n1927 w_4660_n6791.t264 9.52217
R16871 w_4660_n6791.n1927 w_4660_n6791.t386 9.52217
R16872 w_4660_n6791.n2089 w_4660_n6791.t332 9.52217
R16873 w_4660_n6791.n2089 w_4660_n6791.t303 9.52217
R16874 w_4660_n6791.n1930 w_4660_n6791.t340 9.52217
R16875 w_4660_n6791.n1930 w_4660_n6791.t370 9.52217
R16876 w_4660_n6791.n1933 w_4660_n6791.t203 9.52217
R16877 w_4660_n6791.n1933 w_4660_n6791.t378 9.52217
R16878 w_4660_n6791.n1935 w_4660_n6791.t276 9.52217
R16879 w_4660_n6791.n1935 w_4660_n6791.t236 9.52217
R16880 w_4660_n6791.n1937 w_4660_n6791.t330 9.52217
R16881 w_4660_n6791.n1937 w_4660_n6791.t347 9.52217
R16882 w_4660_n6791.n1941 w_4660_n6791.t196 9.52217
R16883 w_4660_n6791.n1941 w_4660_n6791.t367 9.52217
R16884 w_4660_n6791.n1945 w_4660_n6791.t258 9.52217
R16885 w_4660_n6791.n1945 w_4660_n6791.t224 9.52217
R16886 w_4660_n6791.n1949 w_4660_n6791.t272 9.52217
R16887 w_4660_n6791.n1949 w_4660_n6791.t232 9.52217
R16888 w_4660_n6791.n1953 w_4660_n6791.t192 9.52217
R16889 w_4660_n6791.n1953 w_4660_n6791.t354 9.52217
R16890 w_4660_n6791.n1957 w_4660_n6791.t250 9.52217
R16891 w_4660_n6791.n1957 w_4660_n6791.t208 9.52217
R16892 w_4660_n6791.n1960 w_4660_n6791.t263 9.52217
R16893 w_4660_n6791.n1960 w_4660_n6791.t223 9.52217
R16894 w_4660_n6791.n1963 w_4660_n6791.t322 9.52217
R16895 w_4660_n6791.n1963 w_4660_n6791.t300 9.52217
R16896 w_4660_n6791.n2019 w_4660_n6791.t191 9.52217
R16897 w_4660_n6791.n2019 w_4660_n6791.t355 9.52217
R16898 w_4660_n6791.n2012 w_4660_n6791.t256 9.52217
R16899 w_4660_n6791.n2012 w_4660_n6791.t214 9.52217
R16900 w_4660_n6791.n1970 w_4660_n6791.t316 9.52217
R16901 w_4660_n6791.n1970 w_4660_n6791.t283 9.52217
R16902 w_4660_n6791.n1974 w_4660_n6791.t328 9.52217
R16903 w_4660_n6791.n1974 w_4660_n6791.t345 9.52217
R16904 w_4660_n6791.n1977 w_4660_n6791.t247 9.52217
R16905 w_4660_n6791.n1977 w_4660_n6791.t364 9.52217
R16906 w_4660_n6791.n1979 w_4660_n6791.t315 9.52217
R16907 w_4660_n6791.n1979 w_4660_n6791.t280 9.52217
R16908 w_4660_n6791.n1981 w_4660_n6791.t326 9.52217
R16909 w_4660_n6791.n1981 w_4660_n6791.t296 9.52217
R16910 w_4660_n6791.n1986 w_4660_n6791.t440 9.52217
R16911 w_4660_n6791.n1986 w_4660_n6791.t20 9.52217
R16912 w_4660_n6791.n1992 w_4660_n6791.t470 9.52217
R16913 w_4660_n6791.n1992 w_4660_n6791.t452 9.52217
R16914 w_4660_n6791.n1998 w_4660_n6791.t125 9.52217
R16915 w_4660_n6791.n1998 w_4660_n6791.t146 9.52217
R16916 w_4660_n6791.n1972 w_4660_n6791.t461 9.52217
R16917 w_4660_n6791.n1972 w_4660_n6791.t58 9.52217
R16918 w_4660_n6791.n1968 w_4660_n6791.t69 9.52217
R16919 w_4660_n6791.n1968 w_4660_n6791.t10 9.52217
R16920 w_4660_n6791.n1965 w_4660_n6791.t459 9.52217
R16921 w_4660_n6791.n1965 w_4660_n6791.t184 9.52217
R16922 w_4660_n6791.n2024 w_4660_n6791.t82 9.52217
R16923 w_4660_n6791.n2024 w_4660_n6791.t433 9.52217
R16924 w_4660_n6791.n1955 w_4660_n6791.t56 9.52217
R16925 w_4660_n6791.n1955 w_4660_n6791.t414 9.52217
R16926 w_4660_n6791.n1951 w_4660_n6791.t129 9.52217
R16927 w_4660_n6791.n1951 w_4660_n6791.t19 9.52217
R16928 w_4660_n6791.n1947 w_4660_n6791.t472 9.52217
R16929 w_4660_n6791.n1947 w_4660_n6791.t21 9.52217
R16930 w_4660_n6791.n1943 w_4660_n6791.t467 9.52217
R16931 w_4660_n6791.n1943 w_4660_n6791.t474 9.52217
R16932 w_4660_n6791.n1939 w_4660_n6791.t124 9.52217
R16933 w_4660_n6791.n1939 w_4660_n6791.t457 9.52217
R16934 w_4660_n6791.n2069 w_4660_n6791.t473 9.52217
R16935 w_4660_n6791.n2069 w_4660_n6791.t57 9.52217
R16936 w_4660_n6791.n2077 w_4660_n6791.t97 9.52217
R16937 w_4660_n6791.n2077 w_4660_n6791.t22 9.52217
R16938 w_4660_n6791.n310 w_4660_n6791.t410 9.52217
R16939 w_4660_n6791.n310 w_4660_n6791.t435 9.52217
R16940 w_4660_n6791.n311 w_4660_n6791.t14 9.52217
R16941 w_4660_n6791.n311 w_4660_n6791.t93 9.52217
R16942 w_4660_n6791.n312 w_4660_n6791.t134 9.52217
R16943 w_4660_n6791.n312 w_4660_n6791.t131 9.52217
R16944 w_4660_n6791.n2432 w_4660_n6791.t6 9.52217
R16945 w_4660_n6791.n2432 w_4660_n6791.t455 9.52217
R16946 w_4660_n6791.n331 w_4660_n6791.t143 9.52217
R16947 w_4660_n6791.n331 w_4660_n6791.t65 9.52217
R16948 w_4660_n6791.n332 w_4660_n6791.t42 9.52217
R16949 w_4660_n6791.n332 w_4660_n6791.t137 9.52217
R16950 w_4660_n6791.n333 w_4660_n6791.t55 9.52217
R16951 w_4660_n6791.n333 w_4660_n6791.t142 9.52217
R16952 w_4660_n6791.n2393 w_4660_n6791.t412 9.52217
R16953 w_4660_n6791.n2393 w_4660_n6791.t411 9.52217
R16954 w_4660_n6791.n2392 w_4660_n6791.t1 9.52217
R16955 w_4660_n6791.n2392 w_4660_n6791.t448 9.52217
R16956 w_4660_n6791.n357 w_4660_n6791.t415 9.52217
R16957 w_4660_n6791.n357 w_4660_n6791.t165 9.52217
R16958 w_4660_n6791.n358 w_4660_n6791.t12 9.52217
R16959 w_4660_n6791.n358 w_4660_n6791.t113 9.52217
R16960 w_4660_n6791.n359 w_4660_n6791.t450 9.52217
R16961 w_4660_n6791.n359 w_4660_n6791.t409 9.52217
R16962 w_4660_n6791.n2354 w_4660_n6791.t162 9.52217
R16963 w_4660_n6791.n2354 w_4660_n6791.t160 9.52217
R16964 w_4660_n6791.n2353 w_4660_n6791.t91 9.52217
R16965 w_4660_n6791.n2353 w_4660_n6791.t89 9.52217
R16966 w_4660_n6791.n382 w_4660_n6791.t449 9.52217
R16967 w_4660_n6791.n382 w_4660_n6791.t402 9.52217
R16968 w_4660_n6791.n383 w_4660_n6791.t152 9.52217
R16969 w_4660_n6791.n383 w_4660_n6791.t462 9.52217
R16970 w_4660_n6791.n384 w_4660_n6791.t445 9.52217
R16971 w_4660_n6791.n384 w_4660_n6791.t121 9.52217
R16972 w_4660_n6791.n2326 w_4660_n6791.t81 9.52217
R16973 w_4660_n6791.n2326 w_4660_n6791.t431 9.52217
R16974 w_4660_n6791.n404 w_4660_n6791.t105 9.52217
R16975 w_4660_n6791.n404 w_4660_n6791.t442 9.52217
R16976 w_4660_n6791.n405 w_4660_n6791.t108 9.52217
R16977 w_4660_n6791.n405 w_4660_n6791.t427 9.52217
R16978 w_4660_n6791.n406 w_4660_n6791.t429 9.52217
R16979 w_4660_n6791.n406 w_4660_n6791.t180 9.52217
R16980 w_4660_n6791.n2299 w_4660_n6791.t398 9.52217
R16981 w_4660_n6791.n2299 w_4660_n6791.t432 9.52217
R16982 w_4660_n6791.n425 w_4660_n6791.t456 9.52217
R16983 w_4660_n6791.n425 w_4660_n6791.t469 9.52217
R16984 w_4660_n6791.n426 w_4660_n6791.t96 9.52217
R16985 w_4660_n6791.n426 w_4660_n6791.t404 9.52217
R16986 w_4660_n6791.n149 w_4660_n6791.t171 9.52217
R16987 w_4660_n6791.n149 w_4660_n6791.t151 9.52217
R16988 w_4660_n6791.n148 w_4660_n6791.t111 9.52217
R16989 w_4660_n6791.n148 w_4660_n6791.t436 9.52217
R16990 w_4660_n6791.n151 w_4660_n6791.t139 9.52217
R16991 w_4660_n6791.n151 w_4660_n6791.t390 9.52217
R16992 w_4660_n6791.n150 w_4660_n6791.t28 9.52217
R16993 w_4660_n6791.n150 w_4660_n6791.t183 9.52217
R16994 w_4660_n6791.n1661 w_4660_n6791.t46 9.52217
R16995 w_4660_n6791.n1661 w_4660_n6791.t177 9.52217
R16996 w_4660_n6791.n1660 w_4660_n6791.t135 9.52217
R16997 w_4660_n6791.n1660 w_4660_n6791.t466 9.52217
R16998 w_4660_n6791.n1659 w_4660_n6791.t438 9.52217
R16999 w_4660_n6791.n1659 w_4660_n6791.t75 9.52217
R17000 w_4660_n6791.n1658 w_4660_n6791.t9 9.52217
R17001 w_4660_n6791.n1658 w_4660_n6791.t428 9.52217
R17002 w_4660_n6791.n1657 w_4660_n6791.t24 9.52217
R17003 w_4660_n6791.n1657 w_4660_n6791.t104 9.52217
R17004 w_4660_n6791.n1656 w_4660_n6791.t176 9.52217
R17005 w_4660_n6791.n1656 w_4660_n6791.t76 9.52217
R17006 w_4660_n6791.n1655 w_4660_n6791.t133 9.52217
R17007 w_4660_n6791.n1655 w_4660_n6791.t54 9.52217
R17008 w_4660_n6791.n1654 w_4660_n6791.t179 9.52217
R17009 w_4660_n6791.n1654 w_4660_n6791.t74 9.52217
R17010 w_4660_n6791.n1653 w_4660_n6791.t453 9.52217
R17011 w_4660_n6791.n1653 w_4660_n6791.t406 9.52217
R17012 w_4660_n6791.n1652 w_4660_n6791.t16 9.52217
R17013 w_4660_n6791.n1652 w_4660_n6791.t441 9.52217
R17014 w_4660_n6791.n1651 w_4660_n6791.t73 9.52217
R17015 w_4660_n6791.n1651 w_4660_n6791.t99 9.52217
R17016 w_4660_n6791.n1650 w_4660_n6791.t407 9.52217
R17017 w_4660_n6791.n1650 w_4660_n6791.t391 9.52217
R17018 w_4660_n6791.n1649 w_4660_n6791.t126 9.52217
R17019 w_4660_n6791.n1649 w_4660_n6791.t150 9.52217
R17020 w_4660_n6791.n1648 w_4660_n6791.t408 9.52217
R17021 w_4660_n6791.n1648 w_4660_n6791.t36 9.52217
R17022 w_4660_n6791.n1647 w_4660_n6791.t169 9.52217
R17023 w_4660_n6791.n1647 w_4660_n6791.t114 9.52217
R17024 w_4660_n6791.n1646 w_4660_n6791.t443 9.52217
R17025 w_4660_n6791.n1646 w_4660_n6791.t90 9.52217
R17026 w_4660_n6791.n1645 w_4660_n6791.t85 9.52217
R17027 w_4660_n6791.n1645 w_4660_n6791.t157 9.52217
R17028 w_4660_n6791.n1644 w_4660_n6791.t49 9.52217
R17029 w_4660_n6791.n1644 w_4660_n6791.t451 9.52217
R17030 w_4660_n6791.n1643 w_4660_n6791.t403 9.52217
R17031 w_4660_n6791.n1643 w_4660_n6791.t164 9.52217
R17032 w_4660_n6791.n1642 w_4660_n6791.t44 9.52217
R17033 w_4660_n6791.n1642 w_4660_n6791.t174 9.52217
R17034 w_4660_n6791.n1608 w_4660_n6791.t100 9.52217
R17035 w_4660_n6791.n1608 w_4660_n6791.t464 9.52217
R17036 w_4660_n6791.n1607 w_4660_n6791.t140 9.52217
R17037 w_4660_n6791.n1607 w_4660_n6791.t161 9.52217
R17038 w_4660_n6791.n1610 w_4660_n6791.t68 9.52217
R17039 w_4660_n6791.n1610 w_4660_n6791.t478 9.52217
R17040 w_4660_n6791.n1609 w_4660_n6791.t430 9.52217
R17041 w_4660_n6791.n1609 w_4660_n6791.t156 9.52217
R17042 w_4660_n6791.n1612 w_4660_n6791.t117 9.52217
R17043 w_4660_n6791.n1612 w_4660_n6791.t38 9.52217
R17044 w_4660_n6791.n1611 w_4660_n6791.t87 9.52217
R17045 w_4660_n6791.n1611 w_4660_n6791.t393 9.52217
R17046 w_4660_n6791.n1614 w_4660_n6791.t400 9.52217
R17047 w_4660_n6791.n1614 w_4660_n6791.t147 9.52217
R17048 w_4660_n6791.n1613 w_4660_n6791.t475 9.52217
R17049 w_4660_n6791.n1613 w_4660_n6791.t128 9.52217
R17050 w_4660_n6791.n1616 w_4660_n6791.t48 9.52217
R17051 w_4660_n6791.n1616 w_4660_n6791.t392 9.52217
R17052 w_4660_n6791.n1615 w_4660_n6791.t120 9.52217
R17053 w_4660_n6791.n1615 w_4660_n6791.t31 9.52217
R17054 w_4660_n6791.n1618 w_4660_n6791.t4 9.52217
R17055 w_4660_n6791.n1618 w_4660_n6791.t71 9.52217
R17056 w_4660_n6791.n1617 w_4660_n6791.t416 9.52217
R17057 w_4660_n6791.n1617 w_4660_n6791.t127 9.52217
R17058 w_4660_n6791.n1620 w_4660_n6791.t8 9.52217
R17059 w_4660_n6791.n1620 w_4660_n6791.t34 9.52217
R17060 w_4660_n6791.n1619 w_4660_n6791.t418 9.52217
R17061 w_4660_n6791.n1619 w_4660_n6791.t66 9.52217
R17062 w_4660_n6791.n1622 w_4660_n6791.t426 9.52217
R17063 w_4660_n6791.n1622 w_4660_n6791.t95 9.52217
R17064 w_4660_n6791.n1621 w_4660_n6791.t477 9.52217
R17065 w_4660_n6791.n1621 w_4660_n6791.t479 9.52217
R17066 w_4660_n6791.n1624 w_4660_n6791.t173 9.52217
R17067 w_4660_n6791.n1624 w_4660_n6791.t101 9.52217
R17068 w_4660_n6791.n1623 w_4660_n6791.t119 9.52217
R17069 w_4660_n6791.n1623 w_4660_n6791.t61 9.52217
R17070 w_4660_n6791.n1626 w_4660_n6791.t422 9.52217
R17071 w_4660_n6791.n1626 w_4660_n6791.t154 9.52217
R17072 w_4660_n6791.n1625 w_4660_n6791.t397 9.52217
R17073 w_4660_n6791.n1625 w_4660_n6791.t155 9.52217
R17074 w_4660_n6791.n1628 w_4660_n6791.t26 9.52217
R17075 w_4660_n6791.n1628 w_4660_n6791.t167 9.52217
R17076 w_4660_n6791.n1627 w_4660_n6791.t465 9.52217
R17077 w_4660_n6791.n1627 w_4660_n6791.t413 9.52217
R17078 w_4660_n6791.n1630 w_4660_n6791.t18 9.52217
R17079 w_4660_n6791.n1630 w_4660_n6791.t396 9.52217
R17080 w_4660_n6791.n1629 w_4660_n6791.t417 9.52217
R17081 w_4660_n6791.n1629 w_4660_n6791.t405 9.52217
R17082 w_4660_n6791.n688 w_4660_n6791.t270 9.52217
R17083 w_4660_n6791.n688 w_4660_n6791.t252 9.52217
R17084 w_4660_n6791.n687 w_4660_n6791.t110 9.52217
R17085 w_4660_n6791.n687 w_4660_n6791.t149 9.52217
R17086 w_4660_n6791.n690 w_4660_n6791.t344 9.52217
R17087 w_4660_n6791.n690 w_4660_n6791.t197 9.52217
R17088 w_4660_n6791.n689 w_4660_n6791.t471 9.52217
R17089 w_4660_n6791.n689 w_4660_n6791.t186 9.52217
R17090 w_4660_n6791.n692 w_4660_n6791.t335 9.52217
R17091 w_4660_n6791.n692 w_4660_n6791.t339 9.52217
R17092 w_4660_n6791.n691 w_4660_n6791.t181 9.52217
R17093 w_4660_n6791.n691 w_4660_n6791.t138 9.52217
R17094 w_4660_n6791.n694 w_4660_n6791.t260 9.52217
R17095 w_4660_n6791.n694 w_4660_n6791.t329 9.52217
R17096 w_4660_n6791.n693 w_4660_n6791.t420 9.52217
R17097 w_4660_n6791.n693 w_4660_n6791.t40 9.52217
R17098 w_4660_n6791.n696 w_4660_n6791.t216 9.52217
R17099 w_4660_n6791.n696 w_4660_n6791.t201 9.52217
R17100 w_4660_n6791.n695 w_4660_n6791.t458 9.52217
R17101 w_4660_n6791.n695 w_4660_n6791.t389 9.52217
R17102 w_4660_n6791.n698 w_4660_n6791.t207 9.52217
R17103 w_4660_n6791.n698 w_4660_n6791.t210 9.52217
R17104 w_4660_n6791.n697 w_4660_n6791.t476 9.52217
R17105 w_4660_n6791.n697 w_4660_n6791.t53 9.52217
R17106 w_4660_n6791.n700 w_4660_n6791.t289 9.52217
R17107 w_4660_n6791.n700 w_4660_n6791.t205 9.52217
R17108 w_4660_n6791.n699 w_4660_n6791.t29 9.52217
R17109 w_4660_n6791.n699 w_4660_n6791.t454 9.52217
R17110 w_4660_n6791.n702 w_4660_n6791.t281 9.52217
R17111 w_4660_n6791.n702 w_4660_n6791.t285 9.52217
R17112 w_4660_n6791.n701 w_4660_n6791.t175 9.52217
R17113 w_4660_n6791.n701 w_4660_n6791.t172 9.52217
R17114 w_4660_n6791.n704 w_4660_n6791.t269 9.52217
R17115 w_4660_n6791.n704 w_4660_n6791.t277 9.52217
R17116 w_4660_n6791.n703 w_4660_n6791.t153 9.52217
R17117 w_4660_n6791.n703 w_4660_n6791.t185 9.52217
R17118 w_4660_n6791.n706 w_4660_n6791.t371 9.52217
R17119 w_4660_n6791.n706 w_4660_n6791.t231 9.52217
R17120 w_4660_n6791.n705 w_4660_n6791.t446 9.52217
R17121 w_4660_n6791.n705 w_4660_n6791.t51 9.52217
R17122 w_4660_n6791.n708 w_4660_n6791.t357 9.52217
R17123 w_4660_n6791.n708 w_4660_n6791.t362 9.52217
R17124 w_4660_n6791.n707 w_4660_n6791.t158 9.52217
R17125 w_4660_n6791.n707 w_4660_n6791.t170 9.52217
R17126 w_4660_n6791.n710 w_4660_n6791.t302 9.52217
R17127 w_4660_n6791.n710 w_4660_n6791.t350 9.52217
R17128 w_4660_n6791.n709 w_4660_n6791.t394 9.52217
R17129 w_4660_n6791.n709 w_4660_n6791.t178 9.52217
R17130 w_4660_n6791.n712 w_4660_n6791.t215 9.52217
R17131 w_4660_n6791.n712 w_4660_n6791.t219 9.52217
R17132 w_4660_n6791.n711 w_4660_n6791.t84 9.52217
R17133 w_4660_n6791.n711 w_4660_n6791.t80 9.52217
R17134 w_4660_n6791.n714 w_4660_n6791.t227 9.52217
R17135 w_4660_n6791.n714 w_4660_n6791.t238 9.52217
R17136 w_4660_n6791.n713 w_4660_n6791.t115 9.52217
R17137 w_4660_n6791.n713 w_4660_n6791.t421 9.52217
R17138 w_4660_n6791.n716 w_4660_n6791.t382 9.52217
R17139 w_4660_n6791.n716 w_4660_n6791.t387 9.52217
R17140 w_4660_n6791.n715 w_4660_n6791.t444 9.52217
R17141 w_4660_n6791.n715 w_4660_n6791.t59 9.52217
R17142 w_4660_n6791.n718 w_4660_n6791.t306 9.52217
R17143 w_4660_n6791.n718 w_4660_n6791.t309 9.52217
R17144 w_4660_n6791.n717 w_4660_n6791.t63 9.52217
R17145 w_4660_n6791.n717 w_4660_n6791.t103 9.52217
R17146 w_4660_n6791.n720 w_4660_n6791.t243 9.52217
R17147 w_4660_n6791.n720 w_4660_n6791.t299 9.52217
R17148 w_4660_n6791.n719 w_4660_n6791.t106 9.52217
R17149 w_4660_n6791.n719 w_4660_n6791.t399 9.52217
R17150 w_4660_n6791.n722 w_4660_n6791.t190 9.52217
R17151 w_4660_n6791.n722 w_4660_n6791.t230 9.52217
R17152 w_4660_n6791.n721 w_4660_n6791.t3 9.52217
R17153 w_4660_n6791.n721 w_4660_n6791.t439 9.52217
R17154 w_4660_n6791.n724 w_4660_n6791.t384 9.52217
R17155 w_4660_n6791.n724 w_4660_n6791.t188 9.52217
R17156 w_4660_n6791.n723 w_4660_n6791.t32 9.52217
R17157 w_4660_n6791.n723 w_4660_n6791.t423 9.52217
R17158 w_4660_n6791.n726 w_4660_n6791.t320 9.52217
R17159 w_4660_n6791.n726 w_4660_n6791.t324 9.52217
R17160 w_4660_n6791.n725 w_4660_n6791.t182 9.52217
R17161 w_4660_n6791.n725 w_4660_n6791.t419 9.52217
R17162 w_4660_n6791.n728 w_4660_n6791.t246 9.52217
R17163 w_4660_n6791.n728 w_4660_n6791.t318 9.52217
R17164 w_4660_n6791.n727 w_4660_n6791.t132 9.52217
R17165 w_4660_n6791.n727 w_4660_n6791.t401 9.52217
R17166 w_4660_n6791.n730 w_4660_n6791.t375 9.52217
R17167 w_4660_n6791.n730 w_4660_n6791.t237 9.52217
R17168 w_4660_n6791.n729 w_4660_n6791.t437 9.52217
R17169 w_4660_n6791.n729 w_4660_n6791.t145 9.52217
R17170 w_4660_n6791.n732 w_4660_n6791.t360 9.52217
R17171 w_4660_n6791.n732 w_4660_n6791.t368 9.52217
R17172 w_4660_n6791.n731 w_4660_n6791.t27 9.52217
R17173 w_4660_n6791.n731 w_4660_n6791.t424 9.52217
R17174 w_4660_n6791.n734 w_4660_n6791.t287 9.52217
R17175 w_4660_n6791.n734 w_4660_n6791.t293 9.52217
R17176 w_4660_n6791.n733 w_4660_n6791.t116 9.52217
R17177 w_4660_n6791.n733 w_4660_n6791.t395 9.52217
R17178 w_4660_n6791.n1189 w_4660_n6791.t308 9.52217
R17179 w_4660_n6791.n1189 w_4660_n6791.t311 9.52217
R17180 w_4660_n6791.n1188 w_4660_n6791.t268 9.52217
R17181 w_4660_n6791.n1188 w_4660_n6791.t251 9.52217
R17182 w_4660_n6791.n1187 w_4660_n6791.t338 9.52217
R17183 w_4660_n6791.n1187 w_4660_n6791.t211 9.52217
R17184 w_4660_n6791.n1186 w_4660_n6791.t343 9.52217
R17185 w_4660_n6791.n1186 w_4660_n6791.t195 9.52217
R17186 w_4660_n6791.n1185 w_4660_n6791.t271 9.52217
R17187 w_4660_n6791.n1185 w_4660_n6791.t202 9.52217
R17188 w_4660_n6791.n1184 w_4660_n6791.t333 9.52217
R17189 w_4660_n6791.n1184 w_4660_n6791.t337 9.52217
R17190 w_4660_n6791.n1183 w_4660_n6791.t253 9.52217
R17191 w_4660_n6791.n1183 w_4660_n6791.t336 9.52217
R17192 w_4660_n6791.n1182 w_4660_n6791.t259 9.52217
R17193 w_4660_n6791.n1182 w_4660_n6791.t327 9.52217
R17194 w_4660_n6791.n1181 w_4660_n6791.t374 9.52217
R17195 w_4660_n6791.n1181 w_4660_n6791.t376 9.52217
R17196 w_4660_n6791.n1180 w_4660_n6791.t213 9.52217
R17197 w_4660_n6791.n1180 w_4660_n6791.t200 9.52217
R17198 w_4660_n6791.n1179 w_4660_n6791.t305 9.52217
R17199 w_4660_n6791.n1179 w_4660_n6791.t225 9.52217
R17200 w_4660_n6791.n1178 w_4660_n6791.t206 9.52217
R17201 w_4660_n6791.n1178 w_4660_n6791.t209 9.52217
R17202 w_4660_n6791.n1177 w_4660_n6791.t334 9.52217
R17203 w_4660_n6791.n1177 w_4660_n6791.t372 9.52217
R17204 w_4660_n6791.n1176 w_4660_n6791.t288 9.52217
R17205 w_4660_n6791.n1176 w_4660_n6791.t204 9.52217
R17206 w_4660_n6791.n1175 w_4660_n6791.t265 9.52217
R17207 w_4660_n6791.n1175 w_4660_n6791.t199 9.52217
R17208 w_4660_n6791.n1174 w_4660_n6791.t279 9.52217
R17209 w_4660_n6791.n1174 w_4660_n6791.t284 9.52217
R17210 w_4660_n6791.n1173 w_4660_n6791.t198 9.52217
R17211 w_4660_n6791.n1173 w_4660_n6791.t331 9.52217
R17212 w_4660_n6791.n1172 w_4660_n6791.t267 9.52217
R17213 w_4660_n6791.n1172 w_4660_n6791.t275 9.52217
R17214 w_4660_n6791.n1171 w_4660_n6791.t366 9.52217
R17215 w_4660_n6791.n1171 w_4660_n6791.t249 9.52217
R17216 w_4660_n6791.n1170 w_4660_n6791.t369 9.52217
R17217 w_4660_n6791.n1170 w_4660_n6791.t229 9.52217
R17218 w_4660_n6791.n1169 w_4660_n6791.t298 9.52217
R17219 w_4660_n6791.n1169 w_4660_n6791.t222 9.52217
R17220 w_4660_n6791.n1168 w_4660_n6791.t356 9.52217
R17221 w_4660_n6791.n1168 w_4660_n6791.t361 9.52217
R17222 w_4660_n6791.n1167 w_4660_n6791.t282 9.52217
R17223 w_4660_n6791.n1167 w_4660_n6791.t363 9.52217
R17224 w_4660_n6791.n1166 w_4660_n6791.t301 9.52217
R17225 w_4660_n6791.n1166 w_4660_n6791.t348 9.52217
R17226 w_4660_n6791.n1165 w_4660_n6791.t262 9.52217
R17227 w_4660_n6791.n1165 w_4660_n6791.t194 9.52217
R17228 w_4660_n6791.n1164 w_4660_n6791.t212 9.52217
R17229 w_4660_n6791.n1164 w_4660_n6791.t217 9.52217
R17230 w_4660_n6791.n1163 w_4660_n6791.t325 9.52217
R17231 w_4660_n6791.n1163 w_4660_n6791.t261 9.52217
R17232 w_4660_n6791.n1162 w_4660_n6791.t226 9.52217
R17233 w_4660_n6791.n1162 w_4660_n6791.t235 9.52217
R17234 w_4660_n6791.n1161 w_4660_n6791.t314 9.52217
R17235 w_4660_n6791.n1161 w_4660_n6791.t245 9.52217
R17236 w_4660_n6791.n1160 w_4660_n6791.t381 9.52217
R17237 w_4660_n6791.n1160 w_4660_n6791.t385 9.52217
R17238 w_4660_n6791.n1159 w_4660_n6791.t295 9.52217
R17239 w_4660_n6791.n1159 w_4660_n6791.t218 9.52217
R17240 w_4660_n6791.n1158 w_4660_n6791.t304 9.52217
R17241 w_4660_n6791.n1158 w_4660_n6791.t307 9.52217
R17242 w_4660_n6791.n1157 w_4660_n6791.t278 9.52217
R17243 w_4660_n6791.n1157 w_4660_n6791.t358 9.52217
R17244 w_4660_n6791.n1156 w_4660_n6791.t242 9.52217
R17245 w_4660_n6791.n1156 w_4660_n6791.t297 9.52217
R17246 w_4660_n6791.n1155 w_4660_n6791.t193 9.52217
R17247 w_4660_n6791.n1155 w_4660_n6791.t342 9.52217
R17248 w_4660_n6791.n1154 w_4660_n6791.t189 9.52217
R17249 w_4660_n6791.n1154 w_4660_n6791.t228 9.52217
R17250 w_4660_n6791.n1153 w_4660_n6791.t321 9.52217
R17251 w_4660_n6791.n1153 w_4660_n6791.t255 9.52217
R17252 w_4660_n6791.n1152 w_4660_n6791.t383 9.52217
R17253 w_4660_n6791.n1152 w_4660_n6791.t187 9.52217
R17254 w_4660_n6791.n1151 w_4660_n6791.t310 9.52217
R17255 w_4660_n6791.n1151 w_4660_n6791.t234 9.52217
R17256 w_4660_n6791.n1150 w_4660_n6791.t319 9.52217
R17257 w_4660_n6791.n1150 w_4660_n6791.t323 9.52217
R17258 w_4660_n6791.n1149 w_4660_n6791.t290 9.52217
R17259 w_4660_n6791.n1149 w_4660_n6791.t377 9.52217
R17260 w_4660_n6791.n1148 w_4660_n6791.t244 9.52217
R17261 w_4660_n6791.n1148 w_4660_n6791.t317 9.52217
R17262 w_4660_n6791.n1147 w_4660_n6791.t241 9.52217
R17263 w_4660_n6791.n1147 w_4660_n6791.t351 9.52217
R17264 w_4660_n6791.n1146 w_4660_n6791.t373 9.52217
R17265 w_4660_n6791.n1146 w_4660_n6791.t233 9.52217
R17266 w_4660_n6791.n1145 w_4660_n6791.t379 9.52217
R17267 w_4660_n6791.n1145 w_4660_n6791.t313 9.52217
R17268 w_4660_n6791.n1144 w_4660_n6791.t359 9.52217
R17269 w_4660_n6791.n1144 w_4660_n6791.t365 9.52217
R17270 w_4660_n6791.n1143 w_4660_n6791.t352 9.52217
R17271 w_4660_n6791.n1143 w_4660_n6791.t294 9.52217
R17272 w_4660_n6791.n1142 w_4660_n6791.t286 9.52217
R17273 w_4660_n6791.n1142 w_4660_n6791.t292 9.52217
R17274 w_4660_n6791.n2704 w_4660_n6791.t266 9.52217
R17275 w_4660_n6791.t388 w_4660_n6791.n2704 9.52217
R17276 w_4660_n6791.n72 w_4660_n6791.n66 9.3005
R17277 w_4660_n6791.n1474 w_4660_n6791.n1473 9.3005
R17278 w_4660_n6791.n460 w_4660_n6791.n459 9.3005
R17279 w_4660_n6791.n1467 w_4660_n6791.n464 9.3005
R17280 w_4660_n6791.n1460 w_4660_n6791.n463 9.3005
R17281 w_4660_n6791.n1462 w_4660_n6791.n1461 9.3005
R17282 w_4660_n6791.n1459 w_4660_n6791.n466 9.3005
R17283 w_4660_n6791.n1458 w_4660_n6791.n1457 9.3005
R17284 w_4660_n6791.n469 w_4660_n6791.n468 9.3005
R17285 w_4660_n6791.n1453 w_4660_n6791.n1452 9.3005
R17286 w_4660_n6791.n1451 w_4660_n6791.n473 9.3005
R17287 w_4660_n6791.n1450 w_4660_n6791.n1449 9.3005
R17288 w_4660_n6791.n477 w_4660_n6791.n476 9.3005
R17289 w_4660_n6791.n1444 w_4660_n6791.n1443 9.3005
R17290 w_4660_n6791.n1442 w_4660_n6791.n481 9.3005
R17291 w_4660_n6791.n1441 w_4660_n6791.n1440 9.3005
R17292 w_4660_n6791.n485 w_4660_n6791.n484 9.3005
R17293 w_4660_n6791.n1436 w_4660_n6791.n1435 9.3005
R17294 w_4660_n6791.n1434 w_4660_n6791.n489 9.3005
R17295 w_4660_n6791.n1433 w_4660_n6791.n1432 9.3005
R17296 w_4660_n6791.n493 w_4660_n6791.n492 9.3005
R17297 w_4660_n6791.n1428 w_4660_n6791.n1427 9.3005
R17298 w_4660_n6791.n1426 w_4660_n6791.n497 9.3005
R17299 w_4660_n6791.n1425 w_4660_n6791.n1424 9.3005
R17300 w_4660_n6791.n501 w_4660_n6791.n500 9.3005
R17301 w_4660_n6791.n1419 w_4660_n6791.n1418 9.3005
R17302 w_4660_n6791.n70 w_4660_n6791.n66 9.3005
R17303 w_4660_n6791.n74 w_4660_n6791.n71 9.3005
R17304 w_4660_n6791.n141 w_4660_n6791.n138 9.3005
R17305 w_4660_n6791.n2626 w_4660_n6791.n2625 9.3005
R17306 w_4660_n6791.n2627 w_4660_n6791.n137 9.3005
R17307 w_4660_n6791.n2629 w_4660_n6791.n2628 9.3005
R17308 w_4660_n6791.n133 w_4660_n6791.n130 9.3005
R17309 w_4660_n6791.n2634 w_4660_n6791.n2633 9.3005
R17310 w_4660_n6791.n2635 w_4660_n6791.n129 9.3005
R17311 w_4660_n6791.n2637 w_4660_n6791.n2636 9.3005
R17312 w_4660_n6791.n125 w_4660_n6791.n122 9.3005
R17313 w_4660_n6791.n2642 w_4660_n6791.n2641 9.3005
R17314 w_4660_n6791.n2643 w_4660_n6791.n120 9.3005
R17315 w_4660_n6791.n2645 w_4660_n6791.n2644 9.3005
R17316 w_4660_n6791.n121 w_4660_n6791.n118 9.3005
R17317 w_4660_n6791.n1498 w_4660_n6791.n1497 9.3005
R17318 w_4660_n6791.n1499 w_4660_n6791.n1492 9.3005
R17319 w_4660_n6791.n1501 w_4660_n6791.n1500 9.3005
R17320 w_4660_n6791.n1488 w_4660_n6791.n1485 9.3005
R17321 w_4660_n6791.n1506 w_4660_n6791.n1505 9.3005
R17322 w_4660_n6791.n1507 w_4660_n6791.n1484 9.3005
R17323 w_4660_n6791.n1509 w_4660_n6791.n1508 9.3005
R17324 w_4660_n6791.n1480 w_4660_n6791.n1477 9.3005
R17325 w_4660_n6791.n1514 w_4660_n6791.n1513 9.3005
R17326 w_4660_n6791.n1515 w_4660_n6791.n457 9.3005
R17327 w_4660_n6791.n1517 w_4660_n6791.n1516 9.3005
R17328 w_4660_n6791.n1476 w_4660_n6791.n455 9.3005
R17329 w_4660_n6791.n255 w_4660_n6791.n141 9.3005
R17330 w_4660_n6791.n2625 w_4660_n6791.n140 9.3005
R17331 w_4660_n6791.n139 w_4660_n6791.n137 9.3005
R17332 w_4660_n6791.n2629 w_4660_n6791.n136 9.3005
R17333 w_4660_n6791.n135 w_4660_n6791.n133 9.3005
R17334 w_4660_n6791.n2633 w_4660_n6791.n132 9.3005
R17335 w_4660_n6791.n131 w_4660_n6791.n129 9.3005
R17336 w_4660_n6791.n2637 w_4660_n6791.n128 9.3005
R17337 w_4660_n6791.n127 w_4660_n6791.n125 9.3005
R17338 w_4660_n6791.n2641 w_4660_n6791.n124 9.3005
R17339 w_4660_n6791.n123 w_4660_n6791.n120 9.3005
R17340 w_4660_n6791.n2645 w_4660_n6791.n119 9.3005
R17341 w_4660_n6791.n1494 w_4660_n6791.n118 9.3005
R17342 w_4660_n6791.n1497 w_4660_n6791.n1495 9.3005
R17343 w_4660_n6791.n1493 w_4660_n6791.n1492 9.3005
R17344 w_4660_n6791.n1501 w_4660_n6791.n1491 9.3005
R17345 w_4660_n6791.n1490 w_4660_n6791.n1488 9.3005
R17346 w_4660_n6791.n1505 w_4660_n6791.n1487 9.3005
R17347 w_4660_n6791.n1486 w_4660_n6791.n1484 9.3005
R17348 w_4660_n6791.n1509 w_4660_n6791.n1483 9.3005
R17349 w_4660_n6791.n1482 w_4660_n6791.n1480 9.3005
R17350 w_4660_n6791.n1513 w_4660_n6791.n1479 9.3005
R17351 w_4660_n6791.n1478 w_4660_n6791.n457 9.3005
R17352 w_4660_n6791.n1517 w_4660_n6791.n456 9.3005
R17353 w_4660_n6791.n1470 w_4660_n6791.n455 9.3005
R17354 w_4660_n6791.n1473 w_4660_n6791.n1472 9.3005
R17355 w_4660_n6791.n1469 w_4660_n6791.n460 9.3005
R17356 w_4660_n6791.n1468 w_4660_n6791.n1467 9.3005
R17357 w_4660_n6791.n463 w_4660_n6791.n462 9.3005
R17358 w_4660_n6791.n1462 w_4660_n6791.n467 9.3005
R17359 w_4660_n6791.n470 w_4660_n6791.n466 9.3005
R17360 w_4660_n6791.n1457 w_4660_n6791.n471 9.3005
R17361 w_4660_n6791.n474 w_4660_n6791.n469 9.3005
R17362 w_4660_n6791.n1453 w_4660_n6791.n475 9.3005
R17363 w_4660_n6791.n478 w_4660_n6791.n473 9.3005
R17364 w_4660_n6791.n1449 w_4660_n6791.n479 9.3005
R17365 w_4660_n6791.n482 w_4660_n6791.n477 9.3005
R17366 w_4660_n6791.n1444 w_4660_n6791.n483 9.3005
R17367 w_4660_n6791.n486 w_4660_n6791.n481 9.3005
R17368 w_4660_n6791.n1440 w_4660_n6791.n487 9.3005
R17369 w_4660_n6791.n490 w_4660_n6791.n485 9.3005
R17370 w_4660_n6791.n1436 w_4660_n6791.n491 9.3005
R17371 w_4660_n6791.n494 w_4660_n6791.n489 9.3005
R17372 w_4660_n6791.n1432 w_4660_n6791.n495 9.3005
R17373 w_4660_n6791.n498 w_4660_n6791.n493 9.3005
R17374 w_4660_n6791.n1428 w_4660_n6791.n499 9.3005
R17375 w_4660_n6791.n502 w_4660_n6791.n497 9.3005
R17376 w_4660_n6791.n1424 w_4660_n6791.n503 9.3005
R17377 w_4660_n6791.n940 w_4660_n6791.n501 9.3005
R17378 w_4660_n6791.n1419 w_4660_n6791.n941 9.3005
R17379 w_4660_n6791.n76 w_4660_n6791.n66 9.3005
R17380 w_4660_n6791.n75 w_4660_n6791.n74 9.3005
R17381 w_4660_n6791.n1415 w_4660_n6791.n945 9.3005
R17382 w_4660_n6791.n980 w_4660_n6791.n943 9.3005
R17383 w_4660_n6791.n982 w_4660_n6791.n981 9.3005
R17384 w_4660_n6791.n979 w_4660_n6791.n947 9.3005
R17385 w_4660_n6791.n978 w_4660_n6791.n977 9.3005
R17386 w_4660_n6791.n950 w_4660_n6791.n949 9.3005
R17387 w_4660_n6791.n973 w_4660_n6791.n972 9.3005
R17388 w_4660_n6791.n971 w_4660_n6791.n954 9.3005
R17389 w_4660_n6791.n970 w_4660_n6791.n969 9.3005
R17390 w_4660_n6791.n958 w_4660_n6791.n957 9.3005
R17391 w_4660_n6791.n965 w_4660_n6791.n964 9.3005
R17392 w_4660_n6791.n108 w_4660_n6791.n105 9.3005
R17393 w_4660_n6791.n2654 w_4660_n6791.n2653 9.3005
R17394 w_4660_n6791.n2655 w_4660_n6791.n104 9.3005
R17395 w_4660_n6791.n2657 w_4660_n6791.n2656 9.3005
R17396 w_4660_n6791.n100 w_4660_n6791.n97 9.3005
R17397 w_4660_n6791.n2662 w_4660_n6791.n2661 9.3005
R17398 w_4660_n6791.n2663 w_4660_n6791.n96 9.3005
R17399 w_4660_n6791.n2665 w_4660_n6791.n2664 9.3005
R17400 w_4660_n6791.n91 w_4660_n6791.n88 9.3005
R17401 w_4660_n6791.n2670 w_4660_n6791.n2669 9.3005
R17402 w_4660_n6791.n2671 w_4660_n6791.n87 9.3005
R17403 w_4660_n6791.n2673 w_4660_n6791.n2672 9.3005
R17404 w_4660_n6791.n2674 w_4660_n6791.n77 9.3005
R17405 w_4660_n6791.n1416 w_4660_n6791.n1415 9.3005
R17406 w_4660_n6791.n943 w_4660_n6791.n942 9.3005
R17407 w_4660_n6791.n982 w_4660_n6791.n948 9.3005
R17408 w_4660_n6791.n951 w_4660_n6791.n947 9.3005
R17409 w_4660_n6791.n977 w_4660_n6791.n952 9.3005
R17410 w_4660_n6791.n955 w_4660_n6791.n950 9.3005
R17411 w_4660_n6791.n973 w_4660_n6791.n956 9.3005
R17412 w_4660_n6791.n959 w_4660_n6791.n954 9.3005
R17413 w_4660_n6791.n969 w_4660_n6791.n960 9.3005
R17414 w_4660_n6791.n962 w_4660_n6791.n958 9.3005
R17415 w_4660_n6791.n965 w_4660_n6791.n963 9.3005
R17416 w_4660_n6791.n961 w_4660_n6791.n108 9.3005
R17417 w_4660_n6791.n2653 w_4660_n6791.n107 9.3005
R17418 w_4660_n6791.n106 w_4660_n6791.n104 9.3005
R17419 w_4660_n6791.n2657 w_4660_n6791.n103 9.3005
R17420 w_4660_n6791.n102 w_4660_n6791.n100 9.3005
R17421 w_4660_n6791.n2661 w_4660_n6791.n99 9.3005
R17422 w_4660_n6791.n98 w_4660_n6791.n96 9.3005
R17423 w_4660_n6791.n2665 w_4660_n6791.n95 9.3005
R17424 w_4660_n6791.n94 w_4660_n6791.n91 9.3005
R17425 w_4660_n6791.n2669 w_4660_n6791.n90 9.3005
R17426 w_4660_n6791.n89 w_4660_n6791.n87 9.3005
R17427 w_4660_n6791.n2673 w_4660_n6791.n86 9.3005
R17428 w_4660_n6791.n2674 w_4660_n6791.n85 9.3005
R17429 w_4660_n6791.n2679 w_4660_n6791.n2678 9.3005
R17430 w_4660_n6791.n2680 w_4660_n6791.n68 9.3005
R17431 w_4660_n6791.n1 w_4660_n6791.n2681 9.3005
R17432 w_4660_n6791.n2678 w_4660_n6791.n80 9.3005
R17433 w_4660_n6791.n79 w_4660_n6791.n68 9.3005
R17434 w_4660_n6791.n1 w_4660_n6791.n67 9.3005
R17435 w_4660_n6791.n2 w_4660_n6791.n1 1.87786
R17436 w_4660_n6791.n2 w_4660_n6791.n65 5.54729
R17437 w_4660_n6791.n2264 w_4660_n6791.n450 9.3005
R17438 w_4660_n6791.n1770 w_4660_n6791.n449 9.3005
R17439 w_4660_n6791.n2260 w_4660_n6791.n2259 9.3005
R17440 w_4660_n6791.n2258 w_4660_n6791.n2257 9.3005
R17441 w_4660_n6791.n2256 w_4660_n6791.n1771 9.3005
R17442 w_4660_n6791.n1777 w_4660_n6791.n5 9.3005
R17443 w_4660_n6791.n6 w_4660_n6791.n2252 9.3005
R17444 w_4660_n6791.n2251 w_4660_n6791.n2250 9.3005
R17445 w_4660_n6791.n2249 w_4660_n6791.n1778 9.3005
R17446 w_4660_n6791.n1787 w_4660_n6791.n1781 9.3005
R17447 w_4660_n6791.n2245 w_4660_n6791.n2244 9.3005
R17448 w_4660_n6791.n2243 w_4660_n6791.n1786 9.3005
R17449 w_4660_n6791.n2242 w_4660_n6791.n2241 9.3005
R17450 w_4660_n6791.n2238 w_4660_n6791.n1788 9.3005
R17451 w_4660_n6791.n2237 w_4660_n6791.n2236 9.3005
R17452 w_4660_n6791.n2235 w_4660_n6791.n1795 9.3005
R17453 w_4660_n6791.n2234 w_4660_n6791.n2233 9.3005
R17454 w_4660_n6791.n1800 w_4660_n6791.n1796 9.3005
R17455 w_4660_n6791.n2229 w_4660_n6791.n2228 9.3005
R17456 w_4660_n6791.n2227 w_4660_n6791.n1805 9.3005
R17457 w_4660_n6791.n2226 w_4660_n6791.n2225 9.3005
R17458 w_4660_n6791.n1810 w_4660_n6791.n1806 9.3005
R17459 w_4660_n6791.n2221 w_4660_n6791.n2220 9.3005
R17460 w_4660_n6791.n2219 w_4660_n6791.n2218 9.3005
R17461 w_4660_n6791.n2217 w_4660_n6791.n1815 9.3005
R17462 w_4660_n6791.n1824 w_4660_n6791.n1818 9.3005
R17463 w_4660_n6791.n2213 w_4660_n6791.n2212 9.3005
R17464 w_4660_n6791.n2211 w_4660_n6791.n1823 9.3005
R17465 w_4660_n6791.n2210 w_4660_n6791.n2209 9.3005
R17466 w_4660_n6791.n8 w_4660_n6791.n7 9.3005
R17467 w_4660_n6791.n2206 w_4660_n6791.n2205 9.3005
R17468 w_4660_n6791.n2204 w_4660_n6791.n1830 9.3005
R17469 w_4660_n6791.n2203 w_4660_n6791.n2202 9.3005
R17470 w_4660_n6791.n2199 w_4660_n6791.n1831 9.3005
R17471 w_4660_n6791.n2198 w_4660_n6791.n2197 9.3005
R17472 w_4660_n6791.n2196 w_4660_n6791.n1839 9.3005
R17473 w_4660_n6791.n2195 w_4660_n6791.n2194 9.3005
R17474 w_4660_n6791.n1844 w_4660_n6791.n1840 9.3005
R17475 w_4660_n6791.n2190 w_4660_n6791.n2189 9.3005
R17476 w_4660_n6791.n2188 w_4660_n6791.n2187 9.3005
R17477 w_4660_n6791.n2186 w_4660_n6791.n1850 9.3005
R17478 w_4660_n6791.n1858 w_4660_n6791.n1853 9.3005
R17479 w_4660_n6791.n2181 w_4660_n6791.n2180 9.3005
R17480 w_4660_n6791.n2179 w_4660_n6791.n2178 9.3005
R17481 w_4660_n6791.n2177 w_4660_n6791.n1859 9.3005
R17482 w_4660_n6791.n1868 w_4660_n6791.n1862 9.3005
R17483 w_4660_n6791.n2173 w_4660_n6791.n2172 9.3005
R17484 w_4660_n6791.n2171 w_4660_n6791.n1867 9.3005
R17485 w_4660_n6791.n2170 w_4660_n6791.n2169 9.3005
R17486 w_4660_n6791.n2166 w_4660_n6791.n1869 9.3005
R17487 w_4660_n6791.n2165 w_4660_n6791.n2164 9.3005
R17488 w_4660_n6791.n2163 w_4660_n6791.n1876 9.3005
R17489 w_4660_n6791.n2162 w_4660_n6791.n2161 9.3005
R17490 w_4660_n6791.n1880 w_4660_n6791.n1877 9.3005
R17491 w_4660_n6791.n2157 w_4660_n6791.n2156 9.3005
R17492 w_4660_n6791.n2155 w_4660_n6791.n1885 9.3005
R17493 w_4660_n6791.n2154 w_4660_n6791.n2153 9.3005
R17494 w_4660_n6791.n1890 w_4660_n6791.n1886 9.3005
R17495 w_4660_n6791.n2149 w_4660_n6791.n2148 9.3005
R17496 w_4660_n6791.n2147 w_4660_n6791.n2146 9.3005
R17497 w_4660_n6791.n2145 w_4660_n6791.n1895 9.3005
R17498 w_4660_n6791.n1904 w_4660_n6791.n1898 9.3005
R17499 w_4660_n6791.n2141 w_4660_n6791.n2140 9.3005
R17500 w_4660_n6791.n2139 w_4660_n6791.n1903 9.3005
R17501 w_4660_n6791.n2138 w_4660_n6791.n2137 9.3005
R17502 w_4660_n6791.n10 w_4660_n6791.n9 9.3005
R17503 w_4660_n6791.n2133 w_4660_n6791.n2132 9.3005
R17504 w_4660_n6791.n2131 w_4660_n6791.n1910 9.3005
R17505 w_4660_n6791.n2130 w_4660_n6791.n2129 9.3005
R17506 w_4660_n6791.n2126 w_4660_n6791.n1911 9.3005
R17507 w_4660_n6791.n2125 w_4660_n6791.n2124 9.3005
R17508 w_4660_n6791.n2123 w_4660_n6791.n1918 9.3005
R17509 w_4660_n6791.n2122 w_4660_n6791.n2121 9.3005
R17510 w_4660_n6791.n2117 w_4660_n6791.n1920 9.3005
R17511 w_4660_n6791.n1919 w_4660_n6791.n47 9.3005
R17512 w_4660_n6791.n2695 w_4660_n6791.n50 9.3005
R17513 w_4660_n6791.n56 w_4660_n6791.n49 9.3005
R17514 w_4660_n6791.n2691 w_4660_n6791.n2690 9.3005
R17515 w_4660_n6791.n2689 w_4660_n6791.n55 9.3005
R17516 w_4660_n6791.n2688 w_4660_n6791.n2687 9.3005
R17517 w_4660_n6791.n60 w_4660_n6791.n57 9.3005
R17518 w_4660_n6791.n2683 w_4660_n6791.n2682 9.3005
R17519 w_4660_n6791.n2264 w_4660_n6791.n448 9.3005
R17520 w_4660_n6791.n1767 w_4660_n6791.n449 9.3005
R17521 w_4660_n6791.n2260 w_4660_n6791.n1768 9.3005
R17522 w_4660_n6791.n2257 w_4660_n6791.n1772 9.3005
R17523 w_4660_n6791.n2256 w_4660_n6791.n1773 9.3005
R17524 w_4660_n6791.n1775 w_4660_n6791.n5 9.3005
R17525 w_4660_n6791.n6 w_4660_n6791.n1776 9.3005
R17526 w_4660_n6791.n2250 w_4660_n6791.n1779 9.3005
R17527 w_4660_n6791.n2249 w_4660_n6791.n1780 9.3005
R17528 w_4660_n6791.n1784 w_4660_n6791.n1781 9.3005
R17529 w_4660_n6791.n2245 w_4660_n6791.n1785 9.3005
R17530 w_4660_n6791.n1789 w_4660_n6791.n1786 9.3005
R17531 w_4660_n6791.n2241 w_4660_n6791.n1790 9.3005
R17532 w_4660_n6791.n2238 w_4660_n6791.n1793 9.3005
R17533 w_4660_n6791.n2237 w_4660_n6791.n1794 9.3005
R17534 w_4660_n6791.n1798 w_4660_n6791.n1795 9.3005
R17535 w_4660_n6791.n2233 w_4660_n6791.n1799 9.3005
R17536 w_4660_n6791.n1803 w_4660_n6791.n1800 9.3005
R17537 w_4660_n6791.n2229 w_4660_n6791.n1804 9.3005
R17538 w_4660_n6791.n1808 w_4660_n6791.n1805 9.3005
R17539 w_4660_n6791.n2225 w_4660_n6791.n1809 9.3005
R17540 w_4660_n6791.n1812 w_4660_n6791.n1810 9.3005
R17541 w_4660_n6791.n2221 w_4660_n6791.n1813 9.3005
R17542 w_4660_n6791.n2218 w_4660_n6791.n1816 9.3005
R17543 w_4660_n6791.n2217 w_4660_n6791.n1817 9.3005
R17544 w_4660_n6791.n1821 w_4660_n6791.n1818 9.3005
R17545 w_4660_n6791.n2213 w_4660_n6791.n1822 9.3005
R17546 w_4660_n6791.n1825 w_4660_n6791.n1823 9.3005
R17547 w_4660_n6791.n2209 w_4660_n6791.n1826 9.3005
R17548 w_4660_n6791.n8 w_4660_n6791.n1828 9.3005
R17549 w_4660_n6791.n2206 w_4660_n6791.n1829 9.3005
R17550 w_4660_n6791.n1832 w_4660_n6791.n1830 9.3005
R17551 w_4660_n6791.n2202 w_4660_n6791.n1833 9.3005
R17552 w_4660_n6791.n2199 w_4660_n6791.n1837 9.3005
R17553 w_4660_n6791.n2198 w_4660_n6791.n1838 9.3005
R17554 w_4660_n6791.n1842 w_4660_n6791.n1839 9.3005
R17555 w_4660_n6791.n2194 w_4660_n6791.n1843 9.3005
R17556 w_4660_n6791.n1847 w_4660_n6791.n1844 9.3005
R17557 w_4660_n6791.n2190 w_4660_n6791.n1848 9.3005
R17558 w_4660_n6791.n2187 w_4660_n6791.n1851 9.3005
R17559 w_4660_n6791.n2186 w_4660_n6791.n1852 9.3005
R17560 w_4660_n6791.n1855 w_4660_n6791.n1853 9.3005
R17561 w_4660_n6791.n2181 w_4660_n6791.n1856 9.3005
R17562 w_4660_n6791.n2178 w_4660_n6791.n1860 9.3005
R17563 w_4660_n6791.n2177 w_4660_n6791.n1861 9.3005
R17564 w_4660_n6791.n1865 w_4660_n6791.n1862 9.3005
R17565 w_4660_n6791.n2173 w_4660_n6791.n1866 9.3005
R17566 w_4660_n6791.n1870 w_4660_n6791.n1867 9.3005
R17567 w_4660_n6791.n2169 w_4660_n6791.n1871 9.3005
R17568 w_4660_n6791.n2166 w_4660_n6791.n1874 9.3005
R17569 w_4660_n6791.n2165 w_4660_n6791.n1875 9.3005
R17570 w_4660_n6791.n1878 w_4660_n6791.n1876 9.3005
R17571 w_4660_n6791.n2161 w_4660_n6791.n1879 9.3005
R17572 w_4660_n6791.n1883 w_4660_n6791.n1880 9.3005
R17573 w_4660_n6791.n2157 w_4660_n6791.n1884 9.3005
R17574 w_4660_n6791.n1888 w_4660_n6791.n1885 9.3005
R17575 w_4660_n6791.n2153 w_4660_n6791.n1889 9.3005
R17576 w_4660_n6791.n1892 w_4660_n6791.n1890 9.3005
R17577 w_4660_n6791.n2149 w_4660_n6791.n1893 9.3005
R17578 w_4660_n6791.n2146 w_4660_n6791.n1896 9.3005
R17579 w_4660_n6791.n2145 w_4660_n6791.n1897 9.3005
R17580 w_4660_n6791.n1901 w_4660_n6791.n1898 9.3005
R17581 w_4660_n6791.n2141 w_4660_n6791.n1902 9.3005
R17582 w_4660_n6791.n1905 w_4660_n6791.n1903 9.3005
R17583 w_4660_n6791.n2137 w_4660_n6791.n1906 9.3005
R17584 w_4660_n6791.n1908 w_4660_n6791.n10 9.3005
R17585 w_4660_n6791.n2133 w_4660_n6791.n1909 9.3005
R17586 w_4660_n6791.n1912 w_4660_n6791.n1910 9.3005
R17587 w_4660_n6791.n2129 w_4660_n6791.n1913 9.3005
R17588 w_4660_n6791.n2126 w_4660_n6791.n1916 9.3005
R17589 w_4660_n6791.n2125 w_4660_n6791.n1917 9.3005
R17590 w_4660_n6791.n2113 w_4660_n6791.n1918 9.3005
R17591 w_4660_n6791.n2121 w_4660_n6791.n2114 9.3005
R17592 w_4660_n6791.n2117 w_4660_n6791.n2116 9.3005
R17593 w_4660_n6791.n2115 w_4660_n6791.n47 9.3005
R17594 w_4660_n6791.n2695 w_4660_n6791.n48 9.3005
R17595 w_4660_n6791.n53 w_4660_n6791.n49 9.3005
R17596 w_4660_n6791.n2691 w_4660_n6791.n54 9.3005
R17597 w_4660_n6791.n58 w_4660_n6791.n55 9.3005
R17598 w_4660_n6791.n2687 w_4660_n6791.n59 9.3005
R17599 w_4660_n6791.n62 w_4660_n6791.n60 9.3005
R17600 w_4660_n6791.n2683 w_4660_n6791.n63 9.3005
R17601 w_4660_n6791.n83 w_4660_n6791.n68 9.3005
R17602 w_4660_n6791.n82 w_4660_n6791.n78 9.3005
R17603 w_4660_n6791.n2678 w_4660_n6791.n2677 9.3005
R17604 w_4660_n6791.n2675 w_4660_n6791.n2674 9.3005
R17605 w_4660_n6791.n1415 w_4660_n6791.n1414 9.3005
R17606 w_4660_n6791.n984 w_4660_n6791.n943 9.3005
R17607 w_4660_n6791.n983 w_4660_n6791.n982 9.3005
R17608 w_4660_n6791.n947 w_4660_n6791.n946 9.3005
R17609 w_4660_n6791.n977 w_4660_n6791.n976 9.3005
R17610 w_4660_n6791.n975 w_4660_n6791.n950 9.3005
R17611 w_4660_n6791.n974 w_4660_n6791.n973 9.3005
R17612 w_4660_n6791.n954 w_4660_n6791.n953 9.3005
R17613 w_4660_n6791.n969 w_4660_n6791.n968 9.3005
R17614 w_4660_n6791.n967 w_4660_n6791.n958 9.3005
R17615 w_4660_n6791.n966 w_4660_n6791.n965 9.3005
R17616 w_4660_n6791.n109 w_4660_n6791.n108 9.3005
R17617 w_4660_n6791.n2653 w_4660_n6791.n2652 9.3005
R17618 w_4660_n6791.n104 w_4660_n6791.n101 9.3005
R17619 w_4660_n6791.n2658 w_4660_n6791.n2657 9.3005
R17620 w_4660_n6791.n2659 w_4660_n6791.n100 9.3005
R17621 w_4660_n6791.n2661 w_4660_n6791.n2660 9.3005
R17622 w_4660_n6791.n96 w_4660_n6791.n93 9.3005
R17623 w_4660_n6791.n2666 w_4660_n6791.n2665 9.3005
R17624 w_4660_n6791.n2667 w_4660_n6791.n91 9.3005
R17625 w_4660_n6791.n2669 w_4660_n6791.n2668 9.3005
R17626 w_4660_n6791.n92 w_4660_n6791.n87 9.3005
R17627 w_4660_n6791.n2673 w_4660_n6791.n84 9.3005
R17628 w_4660_n6791.n1765 w_4660_n6791.n447 9.3005
R17629 w_4660_n6791.n2264 w_4660_n6791.n2263 9.3005
R17630 w_4660_n6791.n2262 w_4660_n6791.n449 9.3005
R17631 w_4660_n6791.n2261 w_4660_n6791.n2260 9.3005
R17632 w_4660_n6791.n2257 w_4660_n6791.n1766 9.3005
R17633 w_4660_n6791.n2256 w_4660_n6791.n2255 9.3005
R17634 w_4660_n6791.n2254 w_4660_n6791.n5 9.3005
R17635 w_4660_n6791.n2253 w_4660_n6791.n6 9.3005
R17636 w_4660_n6791.n2250 w_4660_n6791.n1774 9.3005
R17637 w_4660_n6791.n2249 w_4660_n6791.n2248 9.3005
R17638 w_4660_n6791.n2247 w_4660_n6791.n1781 9.3005
R17639 w_4660_n6791.n2246 w_4660_n6791.n2245 9.3005
R17640 w_4660_n6791.n1786 w_4660_n6791.n1782 9.3005
R17641 w_4660_n6791.n2241 w_4660_n6791.n2240 9.3005
R17642 w_4660_n6791.n2239 w_4660_n6791.n2238 9.3005
R17643 w_4660_n6791.n2237 w_4660_n6791.n1792 9.3005
R17644 w_4660_n6791.n1801 w_4660_n6791.n1795 9.3005
R17645 w_4660_n6791.n2233 w_4660_n6791.n2232 9.3005
R17646 w_4660_n6791.n2231 w_4660_n6791.n1800 9.3005
R17647 w_4660_n6791.n2230 w_4660_n6791.n2229 9.3005
R17648 w_4660_n6791.n1805 w_4660_n6791.n1802 9.3005
R17649 w_4660_n6791.n2225 w_4660_n6791.n2224 9.3005
R17650 w_4660_n6791.n2223 w_4660_n6791.n1810 9.3005
R17651 w_4660_n6791.n2222 w_4660_n6791.n2221 9.3005
R17652 w_4660_n6791.n2218 w_4660_n6791.n1811 9.3005
R17653 w_4660_n6791.n2217 w_4660_n6791.n2216 9.3005
R17654 w_4660_n6791.n2215 w_4660_n6791.n1818 9.3005
R17655 w_4660_n6791.n2214 w_4660_n6791.n2213 9.3005
R17656 w_4660_n6791.n1823 w_4660_n6791.n1819 9.3005
R17657 w_4660_n6791.n2209 w_4660_n6791.n2208 9.3005
R17658 w_4660_n6791.n2207 w_4660_n6791.n8 9.3005
R17659 w_4660_n6791.n2206 w_4660_n6791.n1827 9.3005
R17660 w_4660_n6791.n1835 w_4660_n6791.n1830 9.3005
R17661 w_4660_n6791.n2202 w_4660_n6791.n2201 9.3005
R17662 w_4660_n6791.n2200 w_4660_n6791.n2199 9.3005
R17663 w_4660_n6791.n2198 w_4660_n6791.n1836 9.3005
R17664 w_4660_n6791.n1845 w_4660_n6791.n1839 9.3005
R17665 w_4660_n6791.n2194 w_4660_n6791.n2193 9.3005
R17666 w_4660_n6791.n2192 w_4660_n6791.n1844 9.3005
R17667 w_4660_n6791.n2191 w_4660_n6791.n2190 9.3005
R17668 w_4660_n6791.n2187 w_4660_n6791.n1846 9.3005
R17669 w_4660_n6791.n2186 w_4660_n6791.n2185 9.3005
R17670 w_4660_n6791.n2183 w_4660_n6791.n1853 9.3005
R17671 w_4660_n6791.n2182 w_4660_n6791.n2181 9.3005
R17672 w_4660_n6791.n2178 w_4660_n6791.n1854 9.3005
R17673 w_4660_n6791.n2177 w_4660_n6791.n2176 9.3005
R17674 w_4660_n6791.n2175 w_4660_n6791.n1862 9.3005
R17675 w_4660_n6791.n2174 w_4660_n6791.n2173 9.3005
R17676 w_4660_n6791.n1867 w_4660_n6791.n1863 9.3005
R17677 w_4660_n6791.n2169 w_4660_n6791.n2168 9.3005
R17678 w_4660_n6791.n2167 w_4660_n6791.n2166 9.3005
R17679 w_4660_n6791.n2165 w_4660_n6791.n1873 9.3005
R17680 w_4660_n6791.n1881 w_4660_n6791.n1876 9.3005
R17681 w_4660_n6791.n2161 w_4660_n6791.n2160 9.3005
R17682 w_4660_n6791.n2159 w_4660_n6791.n1880 9.3005
R17683 w_4660_n6791.n2158 w_4660_n6791.n2157 9.3005
R17684 w_4660_n6791.n1885 w_4660_n6791.n1882 9.3005
R17685 w_4660_n6791.n2153 w_4660_n6791.n2152 9.3005
R17686 w_4660_n6791.n2151 w_4660_n6791.n1890 9.3005
R17687 w_4660_n6791.n2150 w_4660_n6791.n2149 9.3005
R17688 w_4660_n6791.n2146 w_4660_n6791.n1891 9.3005
R17689 w_4660_n6791.n2145 w_4660_n6791.n2144 9.3005
R17690 w_4660_n6791.n2143 w_4660_n6791.n1898 9.3005
R17691 w_4660_n6791.n2142 w_4660_n6791.n2141 9.3005
R17692 w_4660_n6791.n1903 w_4660_n6791.n1899 9.3005
R17693 w_4660_n6791.n2137 w_4660_n6791.n2136 9.3005
R17694 w_4660_n6791.n2135 w_4660_n6791.n10 9.3005
R17695 w_4660_n6791.n2134 w_4660_n6791.n2133 9.3005
R17696 w_4660_n6791.n1910 w_4660_n6791.n1907 9.3005
R17697 w_4660_n6791.n2129 w_4660_n6791.n2128 9.3005
R17698 w_4660_n6791.n2127 w_4660_n6791.n2126 9.3005
R17699 w_4660_n6791.n2125 w_4660_n6791.n1915 9.3005
R17700 w_4660_n6791.n2118 w_4660_n6791.n1918 9.3005
R17701 w_4660_n6791.n2121 w_4660_n6791.n2120 9.3005
R17702 w_4660_n6791.n2119 w_4660_n6791.n2117 9.3005
R17703 w_4660_n6791.n51 w_4660_n6791.n47 9.3005
R17704 w_4660_n6791.n2695 w_4660_n6791.n2694 9.3005
R17705 w_4660_n6791.n2693 w_4660_n6791.n49 9.3005
R17706 w_4660_n6791.n2692 w_4660_n6791.n2691 9.3005
R17707 w_4660_n6791.n55 w_4660_n6791.n52 9.3005
R17708 w_4660_n6791.n2687 w_4660_n6791.n2686 9.3005
R17709 w_4660_n6791.n2685 w_4660_n6791.n60 9.3005
R17710 w_4660_n6791.n2684 w_4660_n6791.n2683 9.3005
R17711 w_4660_n6791.n81 w_4660_n6791.n61 9.3005
R17712 w_4660_n6791.n1222 w_4660_n6791.n1221 9.3005
R17713 w_4660_n6791.n1223 w_4660_n6791.n1140 9.3005
R17714 w_4660_n6791.n1226 w_4660_n6791.n1225 9.3005
R17715 w_4660_n6791.n1224 w_4660_n6791.n1136 9.3005
R17716 w_4660_n6791.n1230 w_4660_n6791.n1138 9.3005
R17717 w_4660_n6791.n1137 w_4660_n6791.n1134 9.3005
R17718 w_4660_n6791.n1234 w_4660_n6791.n1129 9.3005
R17719 w_4660_n6791.n1238 w_4660_n6791.n1237 9.3005
R17720 w_4660_n6791.n1239 w_4660_n6791.n1128 9.3005
R17721 w_4660_n6791.n1241 w_4660_n6791.n1240 9.3005
R17722 w_4660_n6791.n1244 w_4660_n6791.n1126 9.3005
R17723 w_4660_n6791.n1125 w_4660_n6791.n1122 9.3005
R17724 w_4660_n6791.n1248 w_4660_n6791.n1117 9.3005
R17725 w_4660_n6791.n1252 w_4660_n6791.n1251 9.3005
R17726 w_4660_n6791.n1253 w_4660_n6791.n1114 9.3005
R17727 w_4660_n6791.n1255 w_4660_n6791.n1254 9.3005
R17728 w_4660_n6791.n12 w_4660_n6791.n11 9.3005
R17729 w_4660_n6791.n1260 w_4660_n6791.n1259 9.3005
R17730 w_4660_n6791.n1261 w_4660_n6791.n1110 9.3005
R17731 w_4660_n6791.n1263 w_4660_n6791.n1262 9.3005
R17732 w_4660_n6791.n1266 w_4660_n6791.n1108 9.3005
R17733 w_4660_n6791.n1107 w_4660_n6791.n1104 9.3005
R17734 w_4660_n6791.n1270 w_4660_n6791.n1099 9.3005
R17735 w_4660_n6791.n1274 w_4660_n6791.n1273 9.3005
R17736 w_4660_n6791.n1275 w_4660_n6791.n1096 9.3005
R17737 w_4660_n6791.n1278 w_4660_n6791.n1277 9.3005
R17738 w_4660_n6791.n1276 w_4660_n6791.n1092 9.3005
R17739 w_4660_n6791.n1282 w_4660_n6791.n1094 9.3005
R17740 w_4660_n6791.n1093 w_4660_n6791.n1090 9.3005
R17741 w_4660_n6791.n1286 w_4660_n6791.n1085 9.3005
R17742 w_4660_n6791.n1290 w_4660_n6791.n1289 9.3005
R17743 w_4660_n6791.n1291 w_4660_n6791.n1084 9.3005
R17744 w_4660_n6791.n1293 w_4660_n6791.n1292 9.3005
R17745 w_4660_n6791.n1296 w_4660_n6791.n1082 9.3005
R17746 w_4660_n6791.n1081 w_4660_n6791.n1078 9.3005
R17747 w_4660_n6791.n1300 w_4660_n6791.n1073 9.3005
R17748 w_4660_n6791.n1304 w_4660_n6791.n1303 9.3005
R17749 w_4660_n6791.n1305 w_4660_n6791.n1072 9.3005
R17750 w_4660_n6791.n1307 w_4660_n6791.n1306 9.3005
R17751 w_4660_n6791.n1311 w_4660_n6791.n1070 9.3005
R17752 w_4660_n6791.n1069 w_4660_n6791.n1066 9.3005
R17753 w_4660_n6791.n1317 w_4660_n6791.n1316 9.3005
R17754 w_4660_n6791.n1319 w_4660_n6791.n1318 9.3005
R17755 w_4660_n6791.n1322 w_4660_n6791.n1064 9.3005
R17756 w_4660_n6791.n1063 w_4660_n6791.n1060 9.3005
R17757 w_4660_n6791.n1326 w_4660_n6791.n1055 9.3005
R17758 w_4660_n6791.n1330 w_4660_n6791.n1329 9.3005
R17759 w_4660_n6791.n1331 w_4660_n6791.n1052 9.3005
R17760 w_4660_n6791.n1334 w_4660_n6791.n1333 9.3005
R17761 w_4660_n6791.n1332 w_4660_n6791.n1048 9.3005
R17762 w_4660_n6791.n1338 w_4660_n6791.n1050 9.3005
R17763 w_4660_n6791.n1049 w_4660_n6791.n1046 9.3005
R17764 w_4660_n6791.n14 w_4660_n6791.n13 9.3005
R17765 w_4660_n6791.n1345 w_4660_n6791.n1344 9.3005
R17766 w_4660_n6791.n1346 w_4660_n6791.n1042 9.3005
R17767 w_4660_n6791.n1348 w_4660_n6791.n1347 9.3005
R17768 w_4660_n6791.n1351 w_4660_n6791.n1040 9.3005
R17769 w_4660_n6791.n1039 w_4660_n6791.n1036 9.3005
R17770 w_4660_n6791.n1355 w_4660_n6791.n1031 9.3005
R17771 w_4660_n6791.n1359 w_4660_n6791.n1358 9.3005
R17772 w_4660_n6791.n1360 w_4660_n6791.n1028 9.3005
R17773 w_4660_n6791.n1363 w_4660_n6791.n1362 9.3005
R17774 w_4660_n6791.n1361 w_4660_n6791.n1024 9.3005
R17775 w_4660_n6791.n1367 w_4660_n6791.n1026 9.3005
R17776 w_4660_n6791.n1025 w_4660_n6791.n1022 9.3005
R17777 w_4660_n6791.n1371 w_4660_n6791.n1017 9.3005
R17778 w_4660_n6791.n1375 w_4660_n6791.n1374 9.3005
R17779 w_4660_n6791.n1376 w_4660_n6791.n1016 9.3005
R17780 w_4660_n6791.n1378 w_4660_n6791.n1377 9.3005
R17781 w_4660_n6791.n1381 w_4660_n6791.n1014 9.3005
R17782 w_4660_n6791.n1013 w_4660_n6791.n1010 9.3005
R17783 w_4660_n6791.n1385 w_4660_n6791.n1005 9.3005
R17784 w_4660_n6791.n1389 w_4660_n6791.n1388 9.3005
R17785 w_4660_n6791.n1390 w_4660_n6791.n1003 9.3005
R17786 w_4660_n6791.n1393 w_4660_n6791.n1392 9.3005
R17787 w_4660_n6791.n1391 w_4660_n6791.n16 9.3005
R17788 w_4660_n6791.n1397 w_4660_n6791.n1001 9.3005
R17789 w_4660_n6791.n1000 w_4660_n6791.n999 9.3005
R17790 w_4660_n6791.n1401 w_4660_n6791.n994 9.3005
R17791 w_4660_n6791.n1405 w_4660_n6791.n1404 9.3005
R17792 w_4660_n6791.n1406 w_4660_n6791.n993 9.3005
R17793 w_4660_n6791.n1408 w_4660_n6791.n1407 9.3005
R17794 w_4660_n6791.n1221 w_4660_n6791.n1219 9.3005
R17795 w_4660_n6791.n1218 w_4660_n6791.n1140 9.3005
R17796 w_4660_n6791.n1226 w_4660_n6791.n1141 9.3005
R17797 w_4660_n6791.n1136 w_4660_n6791.n1135 9.3005
R17798 w_4660_n6791.n1231 w_4660_n6791.n1230 9.3005
R17799 w_4660_n6791.n1232 w_4660_n6791.n1134 9.3005
R17800 w_4660_n6791.n1234 w_4660_n6791.n1233 9.3005
R17801 w_4660_n6791.n1237 w_4660_n6791.n1132 9.3005
R17802 w_4660_n6791.n1131 w_4660_n6791.n1128 9.3005
R17803 w_4660_n6791.n1241 w_4660_n6791.n1123 9.3005
R17804 w_4660_n6791.n1245 w_4660_n6791.n1244 9.3005
R17805 w_4660_n6791.n1246 w_4660_n6791.n1122 9.3005
R17806 w_4660_n6791.n1248 w_4660_n6791.n1247 9.3005
R17807 w_4660_n6791.n1251 w_4660_n6791.n1120 9.3005
R17808 w_4660_n6791.n1119 w_4660_n6791.n1114 9.3005
R17809 w_4660_n6791.n1255 w_4660_n6791.n1116 9.3005
R17810 w_4660_n6791.n1115 w_4660_n6791.n12 9.3005
R17811 w_4660_n6791.n1259 w_4660_n6791.n1112 9.3005
R17812 w_4660_n6791.n1111 w_4660_n6791.n1110 9.3005
R17813 w_4660_n6791.n1263 w_4660_n6791.n1105 9.3005
R17814 w_4660_n6791.n1267 w_4660_n6791.n1266 9.3005
R17815 w_4660_n6791.n1268 w_4660_n6791.n1104 9.3005
R17816 w_4660_n6791.n1270 w_4660_n6791.n1269 9.3005
R17817 w_4660_n6791.n1273 w_4660_n6791.n1102 9.3005
R17818 w_4660_n6791.n1101 w_4660_n6791.n1096 9.3005
R17819 w_4660_n6791.n1278 w_4660_n6791.n1097 9.3005
R17820 w_4660_n6791.n1092 w_4660_n6791.n1091 9.3005
R17821 w_4660_n6791.n1283 w_4660_n6791.n1282 9.3005
R17822 w_4660_n6791.n1284 w_4660_n6791.n1090 9.3005
R17823 w_4660_n6791.n1286 w_4660_n6791.n1285 9.3005
R17824 w_4660_n6791.n1289 w_4660_n6791.n1088 9.3005
R17825 w_4660_n6791.n1087 w_4660_n6791.n1084 9.3005
R17826 w_4660_n6791.n1293 w_4660_n6791.n1079 9.3005
R17827 w_4660_n6791.n1297 w_4660_n6791.n1296 9.3005
R17828 w_4660_n6791.n1298 w_4660_n6791.n1078 9.3005
R17829 w_4660_n6791.n1300 w_4660_n6791.n1299 9.3005
R17830 w_4660_n6791.n1303 w_4660_n6791.n1076 9.3005
R17831 w_4660_n6791.n1075 w_4660_n6791.n1072 9.3005
R17832 w_4660_n6791.n1307 w_4660_n6791.n1067 9.3005
R17833 w_4660_n6791.n1312 w_4660_n6791.n1311 9.3005
R17834 w_4660_n6791.n1313 w_4660_n6791.n1066 9.3005
R17835 w_4660_n6791.n1316 w_4660_n6791.n1315 9.3005
R17836 w_4660_n6791.n1319 w_4660_n6791.n1061 9.3005
R17837 w_4660_n6791.n1323 w_4660_n6791.n1322 9.3005
R17838 w_4660_n6791.n1324 w_4660_n6791.n1060 9.3005
R17839 w_4660_n6791.n1326 w_4660_n6791.n1325 9.3005
R17840 w_4660_n6791.n1329 w_4660_n6791.n1058 9.3005
R17841 w_4660_n6791.n1057 w_4660_n6791.n1052 9.3005
R17842 w_4660_n6791.n1334 w_4660_n6791.n1053 9.3005
R17843 w_4660_n6791.n1048 w_4660_n6791.n1047 9.3005
R17844 w_4660_n6791.n1339 w_4660_n6791.n1338 9.3005
R17845 w_4660_n6791.n1340 w_4660_n6791.n1046 9.3005
R17846 w_4660_n6791.n14 w_4660_n6791.n1341 9.3005
R17847 w_4660_n6791.n1344 w_4660_n6791.n1044 9.3005
R17848 w_4660_n6791.n1043 w_4660_n6791.n1042 9.3005
R17849 w_4660_n6791.n1348 w_4660_n6791.n1037 9.3005
R17850 w_4660_n6791.n1352 w_4660_n6791.n1351 9.3005
R17851 w_4660_n6791.n1353 w_4660_n6791.n1036 9.3005
R17852 w_4660_n6791.n1355 w_4660_n6791.n1354 9.3005
R17853 w_4660_n6791.n1358 w_4660_n6791.n1034 9.3005
R17854 w_4660_n6791.n1033 w_4660_n6791.n1028 9.3005
R17855 w_4660_n6791.n1363 w_4660_n6791.n1029 9.3005
R17856 w_4660_n6791.n1024 w_4660_n6791.n1023 9.3005
R17857 w_4660_n6791.n1368 w_4660_n6791.n1367 9.3005
R17858 w_4660_n6791.n1369 w_4660_n6791.n1022 9.3005
R17859 w_4660_n6791.n1371 w_4660_n6791.n1370 9.3005
R17860 w_4660_n6791.n1374 w_4660_n6791.n1020 9.3005
R17861 w_4660_n6791.n1019 w_4660_n6791.n1016 9.3005
R17862 w_4660_n6791.n1378 w_4660_n6791.n1011 9.3005
R17863 w_4660_n6791.n1382 w_4660_n6791.n1381 9.3005
R17864 w_4660_n6791.n1383 w_4660_n6791.n1010 9.3005
R17865 w_4660_n6791.n1385 w_4660_n6791.n1384 9.3005
R17866 w_4660_n6791.n1388 w_4660_n6791.n1008 9.3005
R17867 w_4660_n6791.n1007 w_4660_n6791.n1003 9.3005
R17868 w_4660_n6791.n1393 w_4660_n6791.n1004 9.3005
R17869 w_4660_n6791.n16 w_4660_n6791.n15 9.3005
R17870 w_4660_n6791.n1398 w_4660_n6791.n1397 9.3005
R17871 w_4660_n6791.n1399 w_4660_n6791.n999 9.3005
R17872 w_4660_n6791.n1401 w_4660_n6791.n1400 9.3005
R17873 w_4660_n6791.n1404 w_4660_n6791.n997 9.3005
R17874 w_4660_n6791.n996 w_4660_n6791.n993 9.3005
R17875 w_4660_n6791.n1408 w_4660_n6791.n986 9.3005
R17876 w_4660_n6791.n1216 w_4660_n6791.n451 9.3005
R17877 w_4660_n6791.n1411 w_4660_n6791.n991 9.3005
R17878 w_4660_n6791.n988 w_4660_n6791.n985 9.3005
R17879 w_4660_n6791.n1412 w_4660_n6791.n1411 9.3005
R17880 w_4660_n6791.n1221 w_4660_n6791.n1220 9.3005
R17881 w_4660_n6791.n1140 w_4660_n6791.n1139 9.3005
R17882 w_4660_n6791.n1227 w_4660_n6791.n1226 9.3005
R17883 w_4660_n6791.n1228 w_4660_n6791.n1136 9.3005
R17884 w_4660_n6791.n1230 w_4660_n6791.n1229 9.3005
R17885 w_4660_n6791.n1134 w_4660_n6791.n1133 9.3005
R17886 w_4660_n6791.n1235 w_4660_n6791.n1234 9.3005
R17887 w_4660_n6791.n1237 w_4660_n6791.n1236 9.3005
R17888 w_4660_n6791.n1128 w_4660_n6791.n1127 9.3005
R17889 w_4660_n6791.n1242 w_4660_n6791.n1241 9.3005
R17890 w_4660_n6791.n1244 w_4660_n6791.n1243 9.3005
R17891 w_4660_n6791.n1122 w_4660_n6791.n1121 9.3005
R17892 w_4660_n6791.n1249 w_4660_n6791.n1248 9.3005
R17893 w_4660_n6791.n1251 w_4660_n6791.n1250 9.3005
R17894 w_4660_n6791.n1114 w_4660_n6791.n1113 9.3005
R17895 w_4660_n6791.n1256 w_4660_n6791.n1255 9.3005
R17896 w_4660_n6791.n1257 w_4660_n6791.n12 9.3005
R17897 w_4660_n6791.n1259 w_4660_n6791.n1258 9.3005
R17898 w_4660_n6791.n1110 w_4660_n6791.n1109 9.3005
R17899 w_4660_n6791.n1264 w_4660_n6791.n1263 9.3005
R17900 w_4660_n6791.n1266 w_4660_n6791.n1265 9.3005
R17901 w_4660_n6791.n1104 w_4660_n6791.n1103 9.3005
R17902 w_4660_n6791.n1271 w_4660_n6791.n1270 9.3005
R17903 w_4660_n6791.n1273 w_4660_n6791.n1272 9.3005
R17904 w_4660_n6791.n1096 w_4660_n6791.n1095 9.3005
R17905 w_4660_n6791.n1279 w_4660_n6791.n1278 9.3005
R17906 w_4660_n6791.n1280 w_4660_n6791.n1092 9.3005
R17907 w_4660_n6791.n1282 w_4660_n6791.n1281 9.3005
R17908 w_4660_n6791.n1090 w_4660_n6791.n1089 9.3005
R17909 w_4660_n6791.n1287 w_4660_n6791.n1286 9.3005
R17910 w_4660_n6791.n1289 w_4660_n6791.n1288 9.3005
R17911 w_4660_n6791.n1084 w_4660_n6791.n1083 9.3005
R17912 w_4660_n6791.n1294 w_4660_n6791.n1293 9.3005
R17913 w_4660_n6791.n1296 w_4660_n6791.n1295 9.3005
R17914 w_4660_n6791.n1078 w_4660_n6791.n1077 9.3005
R17915 w_4660_n6791.n1301 w_4660_n6791.n1300 9.3005
R17916 w_4660_n6791.n1303 w_4660_n6791.n1302 9.3005
R17917 w_4660_n6791.n1072 w_4660_n6791.n1071 9.3005
R17918 w_4660_n6791.n1308 w_4660_n6791.n1307 9.3005
R17919 w_4660_n6791.n1311 w_4660_n6791.n1310 9.3005
R17920 w_4660_n6791.n1309 w_4660_n6791.n1066 9.3005
R17921 w_4660_n6791.n1316 w_4660_n6791.n1065 9.3005
R17922 w_4660_n6791.n1320 w_4660_n6791.n1319 9.3005
R17923 w_4660_n6791.n1322 w_4660_n6791.n1321 9.3005
R17924 w_4660_n6791.n1060 w_4660_n6791.n1059 9.3005
R17925 w_4660_n6791.n1327 w_4660_n6791.n1326 9.3005
R17926 w_4660_n6791.n1329 w_4660_n6791.n1328 9.3005
R17927 w_4660_n6791.n1052 w_4660_n6791.n1051 9.3005
R17928 w_4660_n6791.n1335 w_4660_n6791.n1334 9.3005
R17929 w_4660_n6791.n1336 w_4660_n6791.n1048 9.3005
R17930 w_4660_n6791.n1338 w_4660_n6791.n1337 9.3005
R17931 w_4660_n6791.n1046 w_4660_n6791.n1045 9.3005
R17932 w_4660_n6791.n1342 w_4660_n6791.n14 9.3005
R17933 w_4660_n6791.n1344 w_4660_n6791.n1343 9.3005
R17934 w_4660_n6791.n1042 w_4660_n6791.n1041 9.3005
R17935 w_4660_n6791.n1349 w_4660_n6791.n1348 9.3005
R17936 w_4660_n6791.n1351 w_4660_n6791.n1350 9.3005
R17937 w_4660_n6791.n1036 w_4660_n6791.n1035 9.3005
R17938 w_4660_n6791.n1356 w_4660_n6791.n1355 9.3005
R17939 w_4660_n6791.n1358 w_4660_n6791.n1357 9.3005
R17940 w_4660_n6791.n1028 w_4660_n6791.n1027 9.3005
R17941 w_4660_n6791.n1364 w_4660_n6791.n1363 9.3005
R17942 w_4660_n6791.n1365 w_4660_n6791.n1024 9.3005
R17943 w_4660_n6791.n1367 w_4660_n6791.n1366 9.3005
R17944 w_4660_n6791.n1022 w_4660_n6791.n1021 9.3005
R17945 w_4660_n6791.n1372 w_4660_n6791.n1371 9.3005
R17946 w_4660_n6791.n1374 w_4660_n6791.n1373 9.3005
R17947 w_4660_n6791.n1016 w_4660_n6791.n1015 9.3005
R17948 w_4660_n6791.n1379 w_4660_n6791.n1378 9.3005
R17949 w_4660_n6791.n1381 w_4660_n6791.n1380 9.3005
R17950 w_4660_n6791.n1010 w_4660_n6791.n1009 9.3005
R17951 w_4660_n6791.n1386 w_4660_n6791.n1385 9.3005
R17952 w_4660_n6791.n1388 w_4660_n6791.n1387 9.3005
R17953 w_4660_n6791.n1003 w_4660_n6791.n1002 9.3005
R17954 w_4660_n6791.n1394 w_4660_n6791.n1393 9.3005
R17955 w_4660_n6791.n1395 w_4660_n6791.n16 9.3005
R17956 w_4660_n6791.n1397 w_4660_n6791.n1396 9.3005
R17957 w_4660_n6791.n999 w_4660_n6791.n998 9.3005
R17958 w_4660_n6791.n1402 w_4660_n6791.n1401 9.3005
R17959 w_4660_n6791.n1404 w_4660_n6791.n1403 9.3005
R17960 w_4660_n6791.n993 w_4660_n6791.n992 9.3005
R17961 w_4660_n6791.n1409 w_4660_n6791.n1408 9.3005
R17962 w_4660_n6791.n1411 w_4660_n6791.n1410 9.3005
R17963 w_4660_n6791.n1420 w_4660_n6791.n1419 9.3005
R17964 w_4660_n6791.n1422 w_4660_n6791.n501 9.3005
R17965 w_4660_n6791.n1473 w_4660_n6791.n461 9.3005
R17966 w_4660_n6791.n1465 w_4660_n6791.n460 9.3005
R17967 w_4660_n6791.n1467 w_4660_n6791.n1466 9.3005
R17968 w_4660_n6791.n1464 w_4660_n6791.n463 9.3005
R17969 w_4660_n6791.n1463 w_4660_n6791.n1462 9.3005
R17970 w_4660_n6791.n466 w_4660_n6791.n465 9.3005
R17971 w_4660_n6791.n1457 w_4660_n6791.n1456 9.3005
R17972 w_4660_n6791.n1455 w_4660_n6791.n469 9.3005
R17973 w_4660_n6791.n1454 w_4660_n6791.n1453 9.3005
R17974 w_4660_n6791.n473 w_4660_n6791.n472 9.3005
R17975 w_4660_n6791.n1449 w_4660_n6791.n1448 9.3005
R17976 w_4660_n6791.n1446 w_4660_n6791.n477 9.3005
R17977 w_4660_n6791.n1445 w_4660_n6791.n1444 9.3005
R17978 w_4660_n6791.n481 w_4660_n6791.n480 9.3005
R17979 w_4660_n6791.n1440 w_4660_n6791.n1439 9.3005
R17980 w_4660_n6791.n1438 w_4660_n6791.n485 9.3005
R17981 w_4660_n6791.n1437 w_4660_n6791.n1436 9.3005
R17982 w_4660_n6791.n489 w_4660_n6791.n488 9.3005
R17983 w_4660_n6791.n1432 w_4660_n6791.n1431 9.3005
R17984 w_4660_n6791.n1430 w_4660_n6791.n493 9.3005
R17985 w_4660_n6791.n1429 w_4660_n6791.n1428 9.3005
R17986 w_4660_n6791.n497 w_4660_n6791.n496 9.3005
R17987 w_4660_n6791.n1424 w_4660_n6791.n1423 9.3005
R17988 w_4660_n6791.n932 w_4660_n6791.n506 9.3005
R17989 w_4660_n6791.n931 w_4660_n6791.n930 9.3005
R17990 w_4660_n6791.n929 w_4660_n6791.n509 9.3005
R17991 w_4660_n6791.n928 w_4660_n6791.n927 9.3005
R17992 w_4660_n6791.n514 w_4660_n6791.n510 9.3005
R17993 w_4660_n6791.n923 w_4660_n6791.n922 9.3005
R17994 w_4660_n6791.n921 w_4660_n6791.n519 9.3005
R17995 w_4660_n6791.n920 w_4660_n6791.n919 9.3005
R17996 w_4660_n6791.n524 w_4660_n6791.n520 9.3005
R17997 w_4660_n6791.n915 w_4660_n6791.n914 9.3005
R17998 w_4660_n6791.n913 w_4660_n6791.n912 9.3005
R17999 w_4660_n6791.n911 w_4660_n6791.n529 9.3005
R18000 w_4660_n6791.n538 w_4660_n6791.n532 9.3005
R18001 w_4660_n6791.n907 w_4660_n6791.n906 9.3005
R18002 w_4660_n6791.n905 w_4660_n6791.n537 9.3005
R18003 w_4660_n6791.n904 w_4660_n6791.n903 9.3005
R18004 w_4660_n6791.n18 w_4660_n6791.n17 9.3005
R18005 w_4660_n6791.n900 w_4660_n6791.n899 9.3005
R18006 w_4660_n6791.n898 w_4660_n6791.n544 9.3005
R18007 w_4660_n6791.n897 w_4660_n6791.n896 9.3005
R18008 w_4660_n6791.n893 w_4660_n6791.n545 9.3005
R18009 w_4660_n6791.n892 w_4660_n6791.n891 9.3005
R18010 w_4660_n6791.n890 w_4660_n6791.n553 9.3005
R18011 w_4660_n6791.n889 w_4660_n6791.n888 9.3005
R18012 w_4660_n6791.n558 w_4660_n6791.n554 9.3005
R18013 w_4660_n6791.n884 w_4660_n6791.n883 9.3005
R18014 w_4660_n6791.n882 w_4660_n6791.n881 9.3005
R18015 w_4660_n6791.n880 w_4660_n6791.n564 9.3005
R18016 w_4660_n6791.n572 w_4660_n6791.n567 9.3005
R18017 w_4660_n6791.n876 w_4660_n6791.n875 9.3005
R18018 w_4660_n6791.n874 w_4660_n6791.n873 9.3005
R18019 w_4660_n6791.n872 w_4660_n6791.n573 9.3005
R18020 w_4660_n6791.n582 w_4660_n6791.n576 9.3005
R18021 w_4660_n6791.n868 w_4660_n6791.n867 9.3005
R18022 w_4660_n6791.n866 w_4660_n6791.n581 9.3005
R18023 w_4660_n6791.n865 w_4660_n6791.n864 9.3005
R18024 w_4660_n6791.n861 w_4660_n6791.n583 9.3005
R18025 w_4660_n6791.n860 w_4660_n6791.n859 9.3005
R18026 w_4660_n6791.n858 w_4660_n6791.n590 9.3005
R18027 w_4660_n6791.n857 w_4660_n6791.n856 9.3005
R18028 w_4660_n6791.n852 w_4660_n6791.n591 9.3005
R18029 w_4660_n6791.n851 w_4660_n6791.n599 9.3005
R18030 w_4660_n6791.n605 w_4660_n6791.n598 9.3005
R18031 w_4660_n6791.n847 w_4660_n6791.n846 9.3005
R18032 w_4660_n6791.n845 w_4660_n6791.n604 9.3005
R18033 w_4660_n6791.n844 w_4660_n6791.n843 9.3005
R18034 w_4660_n6791.n840 w_4660_n6791.n606 9.3005
R18035 w_4660_n6791.n839 w_4660_n6791.n838 9.3005
R18036 w_4660_n6791.n837 w_4660_n6791.n613 9.3005
R18037 w_4660_n6791.n836 w_4660_n6791.n835 9.3005
R18038 w_4660_n6791.n618 w_4660_n6791.n614 9.3005
R18039 w_4660_n6791.n831 w_4660_n6791.n830 9.3005
R18040 w_4660_n6791.n829 w_4660_n6791.n20 9.3005
R18041 w_4660_n6791.n828 w_4660_n6791.n827 9.3005
R18042 w_4660_n6791.n625 w_4660_n6791.n622 9.3005
R18043 w_4660_n6791.n823 w_4660_n6791.n822 9.3005
R18044 w_4660_n6791.n821 w_4660_n6791.n820 9.3005
R18045 w_4660_n6791.n819 w_4660_n6791.n630 9.3005
R18046 w_4660_n6791.n639 w_4660_n6791.n633 9.3005
R18047 w_4660_n6791.n815 w_4660_n6791.n814 9.3005
R18048 w_4660_n6791.n813 w_4660_n6791.n638 9.3005
R18049 w_4660_n6791.n812 w_4660_n6791.n811 9.3005
R18050 w_4660_n6791.n808 w_4660_n6791.n640 9.3005
R18051 w_4660_n6791.n807 w_4660_n6791.n806 9.3005
R18052 w_4660_n6791.n805 w_4660_n6791.n647 9.3005
R18053 w_4660_n6791.n804 w_4660_n6791.n803 9.3005
R18054 w_4660_n6791.n800 w_4660_n6791.n648 9.3005
R18055 w_4660_n6791.n799 w_4660_n6791.n798 9.3005
R18056 w_4660_n6791.n797 w_4660_n6791.n656 9.3005
R18057 w_4660_n6791.n796 w_4660_n6791.n795 9.3005
R18058 w_4660_n6791.n661 w_4660_n6791.n657 9.3005
R18059 w_4660_n6791.n791 w_4660_n6791.n790 9.3005
R18060 w_4660_n6791.n789 w_4660_n6791.n788 9.3005
R18061 w_4660_n6791.n787 w_4660_n6791.n667 9.3005
R18062 w_4660_n6791.n674 w_4660_n6791.n21 9.3005
R18063 w_4660_n6791.n22 w_4660_n6791.n783 9.3005
R18064 w_4660_n6791.n782 w_4660_n6791.n673 9.3005
R18065 w_4660_n6791.n781 w_4660_n6791.n780 9.3005
R18066 w_4660_n6791.n678 w_4660_n6791.n675 9.3005
R18067 w_4660_n6791.n776 w_4660_n6791.n775 9.3005
R18068 w_4660_n6791.n774 w_4660_n6791.n683 9.3005
R18069 w_4660_n6791.n773 w_4660_n6791.n772 9.3005
R18070 w_4660_n6791.n932 w_4660_n6791.n504 9.3005
R18071 w_4660_n6791.n931 w_4660_n6791.n508 9.3005
R18072 w_4660_n6791.n512 w_4660_n6791.n509 9.3005
R18073 w_4660_n6791.n927 w_4660_n6791.n513 9.3005
R18074 w_4660_n6791.n517 w_4660_n6791.n514 9.3005
R18075 w_4660_n6791.n923 w_4660_n6791.n518 9.3005
R18076 w_4660_n6791.n522 w_4660_n6791.n519 9.3005
R18077 w_4660_n6791.n919 w_4660_n6791.n523 9.3005
R18078 w_4660_n6791.n526 w_4660_n6791.n524 9.3005
R18079 w_4660_n6791.n915 w_4660_n6791.n527 9.3005
R18080 w_4660_n6791.n912 w_4660_n6791.n530 9.3005
R18081 w_4660_n6791.n911 w_4660_n6791.n531 9.3005
R18082 w_4660_n6791.n535 w_4660_n6791.n532 9.3005
R18083 w_4660_n6791.n907 w_4660_n6791.n536 9.3005
R18084 w_4660_n6791.n539 w_4660_n6791.n537 9.3005
R18085 w_4660_n6791.n903 w_4660_n6791.n540 9.3005
R18086 w_4660_n6791.n18 w_4660_n6791.n542 9.3005
R18087 w_4660_n6791.n900 w_4660_n6791.n543 9.3005
R18088 w_4660_n6791.n546 w_4660_n6791.n544 9.3005
R18089 w_4660_n6791.n896 w_4660_n6791.n547 9.3005
R18090 w_4660_n6791.n893 w_4660_n6791.n551 9.3005
R18091 w_4660_n6791.n892 w_4660_n6791.n552 9.3005
R18092 w_4660_n6791.n556 w_4660_n6791.n553 9.3005
R18093 w_4660_n6791.n888 w_4660_n6791.n557 9.3005
R18094 w_4660_n6791.n561 w_4660_n6791.n558 9.3005
R18095 w_4660_n6791.n884 w_4660_n6791.n562 9.3005
R18096 w_4660_n6791.n881 w_4660_n6791.n565 9.3005
R18097 w_4660_n6791.n880 w_4660_n6791.n566 9.3005
R18098 w_4660_n6791.n569 w_4660_n6791.n567 9.3005
R18099 w_4660_n6791.n876 w_4660_n6791.n570 9.3005
R18100 w_4660_n6791.n873 w_4660_n6791.n574 9.3005
R18101 w_4660_n6791.n872 w_4660_n6791.n575 9.3005
R18102 w_4660_n6791.n579 w_4660_n6791.n576 9.3005
R18103 w_4660_n6791.n868 w_4660_n6791.n580 9.3005
R18104 w_4660_n6791.n584 w_4660_n6791.n581 9.3005
R18105 w_4660_n6791.n864 w_4660_n6791.n585 9.3005
R18106 w_4660_n6791.n861 w_4660_n6791.n588 9.3005
R18107 w_4660_n6791.n860 w_4660_n6791.n589 9.3005
R18108 w_4660_n6791.n593 w_4660_n6791.n590 9.3005
R18109 w_4660_n6791.n856 w_4660_n6791.n594 9.3005
R18110 w_4660_n6791.n852 w_4660_n6791.n595 9.3005
R18111 w_4660_n6791.n851 w_4660_n6791.n597 9.3005
R18112 w_4660_n6791.n602 w_4660_n6791.n598 9.3005
R18113 w_4660_n6791.n847 w_4660_n6791.n603 9.3005
R18114 w_4660_n6791.n607 w_4660_n6791.n604 9.3005
R18115 w_4660_n6791.n843 w_4660_n6791.n608 9.3005
R18116 w_4660_n6791.n840 w_4660_n6791.n611 9.3005
R18117 w_4660_n6791.n839 w_4660_n6791.n612 9.3005
R18118 w_4660_n6791.n616 w_4660_n6791.n613 9.3005
R18119 w_4660_n6791.n835 w_4660_n6791.n617 9.3005
R18120 w_4660_n6791.n620 w_4660_n6791.n618 9.3005
R18121 w_4660_n6791.n831 w_4660_n6791.n621 9.3005
R18122 w_4660_n6791.n623 w_4660_n6791.n20 9.3005
R18123 w_4660_n6791.n827 w_4660_n6791.n624 9.3005
R18124 w_4660_n6791.n627 w_4660_n6791.n625 9.3005
R18125 w_4660_n6791.n823 w_4660_n6791.n628 9.3005
R18126 w_4660_n6791.n820 w_4660_n6791.n631 9.3005
R18127 w_4660_n6791.n819 w_4660_n6791.n632 9.3005
R18128 w_4660_n6791.n636 w_4660_n6791.n633 9.3005
R18129 w_4660_n6791.n815 w_4660_n6791.n637 9.3005
R18130 w_4660_n6791.n641 w_4660_n6791.n638 9.3005
R18131 w_4660_n6791.n811 w_4660_n6791.n642 9.3005
R18132 w_4660_n6791.n808 w_4660_n6791.n645 9.3005
R18133 w_4660_n6791.n807 w_4660_n6791.n646 9.3005
R18134 w_4660_n6791.n649 w_4660_n6791.n647 9.3005
R18135 w_4660_n6791.n803 w_4660_n6791.n650 9.3005
R18136 w_4660_n6791.n800 w_4660_n6791.n654 9.3005
R18137 w_4660_n6791.n799 w_4660_n6791.n655 9.3005
R18138 w_4660_n6791.n659 w_4660_n6791.n656 9.3005
R18139 w_4660_n6791.n795 w_4660_n6791.n660 9.3005
R18140 w_4660_n6791.n664 w_4660_n6791.n661 9.3005
R18141 w_4660_n6791.n791 w_4660_n6791.n665 9.3005
R18142 w_4660_n6791.n788 w_4660_n6791.n668 9.3005
R18143 w_4660_n6791.n787 w_4660_n6791.n669 9.3005
R18144 w_4660_n6791.n671 w_4660_n6791.n21 9.3005
R18145 w_4660_n6791.n22 w_4660_n6791.n672 9.3005
R18146 w_4660_n6791.n676 w_4660_n6791.n673 9.3005
R18147 w_4660_n6791.n780 w_4660_n6791.n677 9.3005
R18148 w_4660_n6791.n681 w_4660_n6791.n678 9.3005
R18149 w_4660_n6791.n776 w_4660_n6791.n682 9.3005
R18150 w_4660_n6791.n685 w_4660_n6791.n683 9.3005
R18151 w_4660_n6791.n772 w_4660_n6791.n686 9.3005
R18152 w_4660_n6791.n935 w_4660_n6791.n934 9.3005
R18153 w_4660_n6791.n768 w_4660_n6791.n765 9.3005
R18154 w_4660_n6791.n769 w_4660_n6791.n684 9.3005
R18155 w_4660_n6791.n768 w_4660_n6791.n763 9.3005
R18156 w_4660_n6791.n769 w_4660_n6791.n762 9.3005
R18157 w_4660_n6791.n933 w_4660_n6791.n932 9.3005
R18158 w_4660_n6791.n931 w_4660_n6791.n507 9.3005
R18159 w_4660_n6791.n515 w_4660_n6791.n509 9.3005
R18160 w_4660_n6791.n927 w_4660_n6791.n926 9.3005
R18161 w_4660_n6791.n925 w_4660_n6791.n514 9.3005
R18162 w_4660_n6791.n924 w_4660_n6791.n923 9.3005
R18163 w_4660_n6791.n519 w_4660_n6791.n516 9.3005
R18164 w_4660_n6791.n919 w_4660_n6791.n918 9.3005
R18165 w_4660_n6791.n917 w_4660_n6791.n524 9.3005
R18166 w_4660_n6791.n916 w_4660_n6791.n915 9.3005
R18167 w_4660_n6791.n912 w_4660_n6791.n525 9.3005
R18168 w_4660_n6791.n911 w_4660_n6791.n910 9.3005
R18169 w_4660_n6791.n909 w_4660_n6791.n532 9.3005
R18170 w_4660_n6791.n908 w_4660_n6791.n907 9.3005
R18171 w_4660_n6791.n537 w_4660_n6791.n533 9.3005
R18172 w_4660_n6791.n903 w_4660_n6791.n902 9.3005
R18173 w_4660_n6791.n901 w_4660_n6791.n18 9.3005
R18174 w_4660_n6791.n900 w_4660_n6791.n541 9.3005
R18175 w_4660_n6791.n549 w_4660_n6791.n544 9.3005
R18176 w_4660_n6791.n896 w_4660_n6791.n895 9.3005
R18177 w_4660_n6791.n894 w_4660_n6791.n893 9.3005
R18178 w_4660_n6791.n892 w_4660_n6791.n550 9.3005
R18179 w_4660_n6791.n559 w_4660_n6791.n553 9.3005
R18180 w_4660_n6791.n888 w_4660_n6791.n887 9.3005
R18181 w_4660_n6791.n886 w_4660_n6791.n558 9.3005
R18182 w_4660_n6791.n885 w_4660_n6791.n884 9.3005
R18183 w_4660_n6791.n881 w_4660_n6791.n560 9.3005
R18184 w_4660_n6791.n880 w_4660_n6791.n879 9.3005
R18185 w_4660_n6791.n878 w_4660_n6791.n567 9.3005
R18186 w_4660_n6791.n877 w_4660_n6791.n876 9.3005
R18187 w_4660_n6791.n873 w_4660_n6791.n568 9.3005
R18188 w_4660_n6791.n872 w_4660_n6791.n871 9.3005
R18189 w_4660_n6791.n870 w_4660_n6791.n576 9.3005
R18190 w_4660_n6791.n869 w_4660_n6791.n868 9.3005
R18191 w_4660_n6791.n581 w_4660_n6791.n577 9.3005
R18192 w_4660_n6791.n864 w_4660_n6791.n863 9.3005
R18193 w_4660_n6791.n862 w_4660_n6791.n861 9.3005
R18194 w_4660_n6791.n860 w_4660_n6791.n587 9.3005
R18195 w_4660_n6791.n853 w_4660_n6791.n590 9.3005
R18196 w_4660_n6791.n856 w_4660_n6791.n855 9.3005
R18197 w_4660_n6791.n854 w_4660_n6791.n852 9.3005
R18198 w_4660_n6791.n851 w_4660_n6791.n850 9.3005
R18199 w_4660_n6791.n849 w_4660_n6791.n598 9.3005
R18200 w_4660_n6791.n848 w_4660_n6791.n847 9.3005
R18201 w_4660_n6791.n604 w_4660_n6791.n600 9.3005
R18202 w_4660_n6791.n843 w_4660_n6791.n842 9.3005
R18203 w_4660_n6791.n841 w_4660_n6791.n840 9.3005
R18204 w_4660_n6791.n839 w_4660_n6791.n610 9.3005
R18205 w_4660_n6791.n619 w_4660_n6791.n613 9.3005
R18206 w_4660_n6791.n835 w_4660_n6791.n834 9.3005
R18207 w_4660_n6791.n833 w_4660_n6791.n618 9.3005
R18208 w_4660_n6791.n832 w_4660_n6791.n831 9.3005
R18209 w_4660_n6791.n20 w_4660_n6791.n19 9.3005
R18210 w_4660_n6791.n827 w_4660_n6791.n826 9.3005
R18211 w_4660_n6791.n825 w_4660_n6791.n625 9.3005
R18212 w_4660_n6791.n824 w_4660_n6791.n823 9.3005
R18213 w_4660_n6791.n820 w_4660_n6791.n626 9.3005
R18214 w_4660_n6791.n819 w_4660_n6791.n818 9.3005
R18215 w_4660_n6791.n817 w_4660_n6791.n633 9.3005
R18216 w_4660_n6791.n816 w_4660_n6791.n815 9.3005
R18217 w_4660_n6791.n638 w_4660_n6791.n634 9.3005
R18218 w_4660_n6791.n811 w_4660_n6791.n810 9.3005
R18219 w_4660_n6791.n809 w_4660_n6791.n808 9.3005
R18220 w_4660_n6791.n807 w_4660_n6791.n644 9.3005
R18221 w_4660_n6791.n652 w_4660_n6791.n647 9.3005
R18222 w_4660_n6791.n803 w_4660_n6791.n802 9.3005
R18223 w_4660_n6791.n801 w_4660_n6791.n800 9.3005
R18224 w_4660_n6791.n799 w_4660_n6791.n653 9.3005
R18225 w_4660_n6791.n662 w_4660_n6791.n656 9.3005
R18226 w_4660_n6791.n795 w_4660_n6791.n794 9.3005
R18227 w_4660_n6791.n793 w_4660_n6791.n661 9.3005
R18228 w_4660_n6791.n792 w_4660_n6791.n791 9.3005
R18229 w_4660_n6791.n788 w_4660_n6791.n663 9.3005
R18230 w_4660_n6791.n787 w_4660_n6791.n786 9.3005
R18231 w_4660_n6791.n785 w_4660_n6791.n21 9.3005
R18232 w_4660_n6791.n784 w_4660_n6791.n22 9.3005
R18233 w_4660_n6791.n673 w_4660_n6791.n670 9.3005
R18234 w_4660_n6791.n780 w_4660_n6791.n779 9.3005
R18235 w_4660_n6791.n778 w_4660_n6791.n678 9.3005
R18236 w_4660_n6791.n777 w_4660_n6791.n776 9.3005
R18237 w_4660_n6791.n683 w_4660_n6791.n679 9.3005
R18238 w_4660_n6791.n772 w_4660_n6791.n771 9.3005
R18239 w_4660_n6791.n770 w_4660_n6791.n769 9.3005
R18240 w_4660_n6791.n455 w_4660_n6791.n453 9.3005
R18241 w_4660_n6791.n1518 w_4660_n6791.n1517 9.3005
R18242 w_4660_n6791.n2623 w_4660_n6791.n141 9.3005
R18243 w_4660_n6791.n2625 w_4660_n6791.n2624 9.3005
R18244 w_4660_n6791.n137 w_4660_n6791.n134 9.3005
R18245 w_4660_n6791.n2630 w_4660_n6791.n2629 9.3005
R18246 w_4660_n6791.n2631 w_4660_n6791.n133 9.3005
R18247 w_4660_n6791.n2633 w_4660_n6791.n2632 9.3005
R18248 w_4660_n6791.n129 w_4660_n6791.n126 9.3005
R18249 w_4660_n6791.n2638 w_4660_n6791.n2637 9.3005
R18250 w_4660_n6791.n2639 w_4660_n6791.n125 9.3005
R18251 w_4660_n6791.n2641 w_4660_n6791.n2640 9.3005
R18252 w_4660_n6791.n120 w_4660_n6791.n117 9.3005
R18253 w_4660_n6791.n2646 w_4660_n6791.n2645 9.3005
R18254 w_4660_n6791.n118 w_4660_n6791.n116 9.3005
R18255 w_4660_n6791.n1497 w_4660_n6791.n1496 9.3005
R18256 w_4660_n6791.n1492 w_4660_n6791.n1489 9.3005
R18257 w_4660_n6791.n1502 w_4660_n6791.n1501 9.3005
R18258 w_4660_n6791.n1503 w_4660_n6791.n1488 9.3005
R18259 w_4660_n6791.n1505 w_4660_n6791.n1504 9.3005
R18260 w_4660_n6791.n1484 w_4660_n6791.n1481 9.3005
R18261 w_4660_n6791.n1510 w_4660_n6791.n1509 9.3005
R18262 w_4660_n6791.n1511 w_4660_n6791.n1480 9.3005
R18263 w_4660_n6791.n1513 w_4660_n6791.n1512 9.3005
R18264 w_4660_n6791.n457 w_4660_n6791.n454 9.3005
R18265 w_4660_n6791.n1757 w_4660_n6791.n1756 9.3005
R18266 w_4660_n6791.n1755 w_4660_n6791.n1524 9.3005
R18267 w_4660_n6791.n1532 w_4660_n6791.n1526 9.3005
R18268 w_4660_n6791.n1751 w_4660_n6791.n1750 9.3005
R18269 w_4660_n6791.n1749 w_4660_n6791.n1531 9.3005
R18270 w_4660_n6791.n1748 w_4660_n6791.n1747 9.3005
R18271 w_4660_n6791.n24 w_4660_n6791.n23 9.3005
R18272 w_4660_n6791.n1743 w_4660_n6791.n1742 9.3005
R18273 w_4660_n6791.n1741 w_4660_n6791.n1538 9.3005
R18274 w_4660_n6791.n1740 w_4660_n6791.n1739 9.3005
R18275 w_4660_n6791.n1736 w_4660_n6791.n1539 9.3005
R18276 w_4660_n6791.n1735 w_4660_n6791.n1734 9.3005
R18277 w_4660_n6791.n1733 w_4660_n6791.n1546 9.3005
R18278 w_4660_n6791.n1732 w_4660_n6791.n1731 9.3005
R18279 w_4660_n6791.n1551 w_4660_n6791.n1547 9.3005
R18280 w_4660_n6791.n1727 w_4660_n6791.n1726 9.3005
R18281 w_4660_n6791.n1725 w_4660_n6791.n1724 9.3005
R18282 w_4660_n6791.n1723 w_4660_n6791.n1557 9.3005
R18283 w_4660_n6791.n1565 w_4660_n6791.n1560 9.3005
R18284 w_4660_n6791.n1719 w_4660_n6791.n1718 9.3005
R18285 w_4660_n6791.n1717 w_4660_n6791.n1716 9.3005
R18286 w_4660_n6791.n1715 w_4660_n6791.n1566 9.3005
R18287 w_4660_n6791.n1575 w_4660_n6791.n1569 9.3005
R18288 w_4660_n6791.n1711 w_4660_n6791.n1710 9.3005
R18289 w_4660_n6791.n1709 w_4660_n6791.n1574 9.3005
R18290 w_4660_n6791.n1708 w_4660_n6791.n1707 9.3005
R18291 w_4660_n6791.n1704 w_4660_n6791.n1576 9.3005
R18292 w_4660_n6791.n1703 w_4660_n6791.n1702 9.3005
R18293 w_4660_n6791.n1701 w_4660_n6791.n25 9.3005
R18294 w_4660_n6791.n1700 w_4660_n6791.n26 9.3005
R18295 w_4660_n6791.n1586 w_4660_n6791.n1583 9.3005
R18296 w_4660_n6791.n1696 w_4660_n6791.n1695 9.3005
R18297 w_4660_n6791.n1694 w_4660_n6791.n1591 9.3005
R18298 w_4660_n6791.n1693 w_4660_n6791.n1692 9.3005
R18299 w_4660_n6791.n1596 w_4660_n6791.n1592 9.3005
R18300 w_4660_n6791.n1688 w_4660_n6791.n1687 9.3005
R18301 w_4660_n6791.n1686 w_4660_n6791.n1685 9.3005
R18302 w_4660_n6791.n1684 w_4660_n6791.n1601 9.3005
R18303 w_4660_n6791.n1677 w_4660_n6791.n1604 9.3005
R18304 w_4660_n6791.n1680 w_4660_n6791.n1679 9.3005
R18305 w_4660_n6791.n1678 w_4660_n6791.n1676 9.3005
R18306 w_4660_n6791.n242 w_4660_n6791.n233 9.3005
R18307 w_4660_n6791.n2526 w_4660_n6791.n228 9.3005
R18308 w_4660_n6791.n2530 w_4660_n6791.n2529 9.3005
R18309 w_4660_n6791.n2531 w_4660_n6791.n227 9.3005
R18310 w_4660_n6791.n2533 w_4660_n6791.n2532 9.3005
R18311 w_4660_n6791.n2536 w_4660_n6791.n225 9.3005
R18312 w_4660_n6791.n224 w_4660_n6791.n221 9.3005
R18313 w_4660_n6791.n2540 w_4660_n6791.n216 9.3005
R18314 w_4660_n6791.n2544 w_4660_n6791.n2543 9.3005
R18315 w_4660_n6791.n2545 w_4660_n6791.n212 9.3005
R18316 w_4660_n6791.n2547 w_4660_n6791.n2546 9.3005
R18317 w_4660_n6791.n208 w_4660_n6791.n207 9.3005
R18318 w_4660_n6791.n2552 w_4660_n6791.n2551 9.3005
R18319 w_4660_n6791.n2553 w_4660_n6791.n206 9.3005
R18320 w_4660_n6791.n2555 w_4660_n6791.n2554 9.3005
R18321 w_4660_n6791.n2558 w_4660_n6791.n204 9.3005
R18322 w_4660_n6791.n203 w_4660_n6791.n200 9.3005
R18323 w_4660_n6791.n2562 w_4660_n6791.n195 9.3005
R18324 w_4660_n6791.n2566 w_4660_n6791.n2565 9.3005
R18325 w_4660_n6791.n2567 w_4660_n6791.n191 9.3005
R18326 w_4660_n6791.n2569 w_4660_n6791.n2568 9.3005
R18327 w_4660_n6791.n187 w_4660_n6791.n186 9.3005
R18328 w_4660_n6791.n2574 w_4660_n6791.n2573 9.3005
R18329 w_4660_n6791.n2575 w_4660_n6791.n185 9.3005
R18330 w_4660_n6791.n28 w_4660_n6791.n2576 9.3005
R18331 w_4660_n6791.n2579 w_4660_n6791.n183 9.3005
R18332 w_4660_n6791.n182 w_4660_n6791.n181 9.3005
R18333 w_4660_n6791.n2583 w_4660_n6791.n176 9.3005
R18334 w_4660_n6791.n2587 w_4660_n6791.n2586 9.3005
R18335 w_4660_n6791.n2588 w_4660_n6791.n175 9.3005
R18336 w_4660_n6791.n2590 w_4660_n6791.n2589 9.3005
R18337 w_4660_n6791.n2593 w_4660_n6791.n173 9.3005
R18338 w_4660_n6791.n172 w_4660_n6791.n169 9.3005
R18339 w_4660_n6791.n2597 w_4660_n6791.n164 9.3005
R18340 w_4660_n6791.n2601 w_4660_n6791.n2600 9.3005
R18341 w_4660_n6791.n2602 w_4660_n6791.n161 9.3005
R18342 w_4660_n6791.n2605 w_4660_n6791.n2604 9.3005
R18343 w_4660_n6791.n2603 w_4660_n6791.n153 9.3005
R18344 w_4660_n6791.n2611 w_4660_n6791.n159 9.3005
R18345 w_4660_n6791.n158 w_4660_n6791.n157 9.3005
R18346 w_4660_n6791.n147 w_4660_n6791.n146 9.3005
R18347 w_4660_n6791.n1756 w_4660_n6791.n1522 9.3005
R18348 w_4660_n6791.n1755 w_4660_n6791.n1525 9.3005
R18349 w_4660_n6791.n1529 w_4660_n6791.n1526 9.3005
R18350 w_4660_n6791.n1751 w_4660_n6791.n1530 9.3005
R18351 w_4660_n6791.n1533 w_4660_n6791.n1531 9.3005
R18352 w_4660_n6791.n1747 w_4660_n6791.n1534 9.3005
R18353 w_4660_n6791.n1536 w_4660_n6791.n24 9.3005
R18354 w_4660_n6791.n1743 w_4660_n6791.n1537 9.3005
R18355 w_4660_n6791.n1540 w_4660_n6791.n1538 9.3005
R18356 w_4660_n6791.n1739 w_4660_n6791.n1541 9.3005
R18357 w_4660_n6791.n1736 w_4660_n6791.n1544 9.3005
R18358 w_4660_n6791.n1735 w_4660_n6791.n1545 9.3005
R18359 w_4660_n6791.n1549 w_4660_n6791.n1546 9.3005
R18360 w_4660_n6791.n1731 w_4660_n6791.n1550 9.3005
R18361 w_4660_n6791.n1554 w_4660_n6791.n1551 9.3005
R18362 w_4660_n6791.n1727 w_4660_n6791.n1555 9.3005
R18363 w_4660_n6791.n1724 w_4660_n6791.n1558 9.3005
R18364 w_4660_n6791.n1723 w_4660_n6791.n1559 9.3005
R18365 w_4660_n6791.n1562 w_4660_n6791.n1560 9.3005
R18366 w_4660_n6791.n1719 w_4660_n6791.n1563 9.3005
R18367 w_4660_n6791.n1716 w_4660_n6791.n1567 9.3005
R18368 w_4660_n6791.n1715 w_4660_n6791.n1568 9.3005
R18369 w_4660_n6791.n1572 w_4660_n6791.n1569 9.3005
R18370 w_4660_n6791.n1711 w_4660_n6791.n1573 9.3005
R18371 w_4660_n6791.n1577 w_4660_n6791.n1574 9.3005
R18372 w_4660_n6791.n1707 w_4660_n6791.n1578 9.3005
R18373 w_4660_n6791.n1704 w_4660_n6791.n1581 9.3005
R18374 w_4660_n6791.n1703 w_4660_n6791.n1582 9.3005
R18375 w_4660_n6791.n1584 w_4660_n6791.n25 9.3005
R18376 w_4660_n6791.n26 w_4660_n6791.n1585 9.3005
R18377 w_4660_n6791.n1589 w_4660_n6791.n1586 9.3005
R18378 w_4660_n6791.n1696 w_4660_n6791.n1590 9.3005
R18379 w_4660_n6791.n1594 w_4660_n6791.n1591 9.3005
R18380 w_4660_n6791.n1692 w_4660_n6791.n1595 9.3005
R18381 w_4660_n6791.n1598 w_4660_n6791.n1596 9.3005
R18382 w_4660_n6791.n1688 w_4660_n6791.n1599 9.3005
R18383 w_4660_n6791.n1685 w_4660_n6791.n1602 9.3005
R18384 w_4660_n6791.n1684 w_4660_n6791.n1603 9.3005
R18385 w_4660_n6791.n1674 w_4660_n6791.n1604 9.3005
R18386 w_4660_n6791.n1680 w_4660_n6791.n1675 9.3005
R18387 w_4660_n6791.n1676 w_4660_n6791.n234 9.3005
R18388 w_4660_n6791.n2524 w_4660_n6791.n233 9.3005
R18389 w_4660_n6791.n2526 w_4660_n6791.n2525 9.3005
R18390 w_4660_n6791.n2529 w_4660_n6791.n231 9.3005
R18391 w_4660_n6791.n230 w_4660_n6791.n227 9.3005
R18392 w_4660_n6791.n2533 w_4660_n6791.n222 9.3005
R18393 w_4660_n6791.n2537 w_4660_n6791.n2536 9.3005
R18394 w_4660_n6791.n2538 w_4660_n6791.n221 9.3005
R18395 w_4660_n6791.n2540 w_4660_n6791.n2539 9.3005
R18396 w_4660_n6791.n2543 w_4660_n6791.n219 9.3005
R18397 w_4660_n6791.n218 w_4660_n6791.n212 9.3005
R18398 w_4660_n6791.n2547 w_4660_n6791.n214 9.3005
R18399 w_4660_n6791.n213 w_4660_n6791.n208 9.3005
R18400 w_4660_n6791.n2551 w_4660_n6791.n210 9.3005
R18401 w_4660_n6791.n209 w_4660_n6791.n206 9.3005
R18402 w_4660_n6791.n2555 w_4660_n6791.n201 9.3005
R18403 w_4660_n6791.n2559 w_4660_n6791.n2558 9.3005
R18404 w_4660_n6791.n2560 w_4660_n6791.n200 9.3005
R18405 w_4660_n6791.n2562 w_4660_n6791.n2561 9.3005
R18406 w_4660_n6791.n2565 w_4660_n6791.n198 9.3005
R18407 w_4660_n6791.n197 w_4660_n6791.n191 9.3005
R18408 w_4660_n6791.n2569 w_4660_n6791.n193 9.3005
R18409 w_4660_n6791.n192 w_4660_n6791.n187 9.3005
R18410 w_4660_n6791.n2573 w_4660_n6791.n189 9.3005
R18411 w_4660_n6791.n188 w_4660_n6791.n185 9.3005
R18412 w_4660_n6791.n28 w_4660_n6791.n27 9.3005
R18413 w_4660_n6791.n2580 w_4660_n6791.n2579 9.3005
R18414 w_4660_n6791.n2581 w_4660_n6791.n181 9.3005
R18415 w_4660_n6791.n2583 w_4660_n6791.n2582 9.3005
R18416 w_4660_n6791.n2586 w_4660_n6791.n179 9.3005
R18417 w_4660_n6791.n178 w_4660_n6791.n175 9.3005
R18418 w_4660_n6791.n2590 w_4660_n6791.n170 9.3005
R18419 w_4660_n6791.n2594 w_4660_n6791.n2593 9.3005
R18420 w_4660_n6791.n2595 w_4660_n6791.n169 9.3005
R18421 w_4660_n6791.n2597 w_4660_n6791.n2596 9.3005
R18422 w_4660_n6791.n2600 w_4660_n6791.n167 9.3005
R18423 w_4660_n6791.n166 w_4660_n6791.n161 9.3005
R18424 w_4660_n6791.n2605 w_4660_n6791.n163 9.3005
R18425 w_4660_n6791.n162 w_4660_n6791.n153 9.3005
R18426 w_4660_n6791.n2611 w_4660_n6791.n154 9.3005
R18427 w_4660_n6791.n157 w_4660_n6791.n156 9.3005
R18428 w_4660_n6791.n155 w_4660_n6791.n147 9.3005
R18429 w_4660_n6791.n1756 w_4660_n6791.n1521 9.3005
R18430 w_4660_n6791.n1755 w_4660_n6791.n1754 9.3005
R18431 w_4660_n6791.n1753 w_4660_n6791.n1526 9.3005
R18432 w_4660_n6791.n1752 w_4660_n6791.n1751 9.3005
R18433 w_4660_n6791.n1531 w_4660_n6791.n1527 9.3005
R18434 w_4660_n6791.n1747 w_4660_n6791.n1746 9.3005
R18435 w_4660_n6791.n1745 w_4660_n6791.n24 9.3005
R18436 w_4660_n6791.n1744 w_4660_n6791.n1743 9.3005
R18437 w_4660_n6791.n1538 w_4660_n6791.n1535 9.3005
R18438 w_4660_n6791.n1739 w_4660_n6791.n1738 9.3005
R18439 w_4660_n6791.n1737 w_4660_n6791.n1736 9.3005
R18440 w_4660_n6791.n1735 w_4660_n6791.n1543 9.3005
R18441 w_4660_n6791.n1552 w_4660_n6791.n1546 9.3005
R18442 w_4660_n6791.n1731 w_4660_n6791.n1730 9.3005
R18443 w_4660_n6791.n1729 w_4660_n6791.n1551 9.3005
R18444 w_4660_n6791.n1728 w_4660_n6791.n1727 9.3005
R18445 w_4660_n6791.n1724 w_4660_n6791.n1553 9.3005
R18446 w_4660_n6791.n1723 w_4660_n6791.n1722 9.3005
R18447 w_4660_n6791.n1721 w_4660_n6791.n1560 9.3005
R18448 w_4660_n6791.n1720 w_4660_n6791.n1719 9.3005
R18449 w_4660_n6791.n1716 w_4660_n6791.n1561 9.3005
R18450 w_4660_n6791.n1715 w_4660_n6791.n1714 9.3005
R18451 w_4660_n6791.n1713 w_4660_n6791.n1569 9.3005
R18452 w_4660_n6791.n1712 w_4660_n6791.n1711 9.3005
R18453 w_4660_n6791.n1574 w_4660_n6791.n1570 9.3005
R18454 w_4660_n6791.n1707 w_4660_n6791.n1706 9.3005
R18455 w_4660_n6791.n1705 w_4660_n6791.n1704 9.3005
R18456 w_4660_n6791.n1703 w_4660_n6791.n1580 9.3005
R18457 w_4660_n6791.n1587 w_4660_n6791.n25 9.3005
R18458 w_4660_n6791.n26 w_4660_n6791.n1699 9.3005
R18459 w_4660_n6791.n1698 w_4660_n6791.n1586 9.3005
R18460 w_4660_n6791.n1697 w_4660_n6791.n1696 9.3005
R18461 w_4660_n6791.n1591 w_4660_n6791.n1588 9.3005
R18462 w_4660_n6791.n1692 w_4660_n6791.n1691 9.3005
R18463 w_4660_n6791.n1690 w_4660_n6791.n1596 9.3005
R18464 w_4660_n6791.n1689 w_4660_n6791.n1688 9.3005
R18465 w_4660_n6791.n1685 w_4660_n6791.n1597 9.3005
R18466 w_4660_n6791.n1684 w_4660_n6791.n1683 9.3005
R18467 w_4660_n6791.n1682 w_4660_n6791.n1604 9.3005
R18468 w_4660_n6791.n1681 w_4660_n6791.n1680 9.3005
R18469 w_4660_n6791.n1676 w_4660_n6791.n1606 9.3005
R18470 w_4660_n6791.n233 w_4660_n6791.n232 9.3005
R18471 w_4660_n6791.n2527 w_4660_n6791.n2526 9.3005
R18472 w_4660_n6791.n2529 w_4660_n6791.n2528 9.3005
R18473 w_4660_n6791.n227 w_4660_n6791.n226 9.3005
R18474 w_4660_n6791.n2534 w_4660_n6791.n2533 9.3005
R18475 w_4660_n6791.n2536 w_4660_n6791.n2535 9.3005
R18476 w_4660_n6791.n221 w_4660_n6791.n220 9.3005
R18477 w_4660_n6791.n2541 w_4660_n6791.n2540 9.3005
R18478 w_4660_n6791.n2543 w_4660_n6791.n2542 9.3005
R18479 w_4660_n6791.n212 w_4660_n6791.n211 9.3005
R18480 w_4660_n6791.n2548 w_4660_n6791.n2547 9.3005
R18481 w_4660_n6791.n2549 w_4660_n6791.n208 9.3005
R18482 w_4660_n6791.n2551 w_4660_n6791.n2550 9.3005
R18483 w_4660_n6791.n206 w_4660_n6791.n205 9.3005
R18484 w_4660_n6791.n2556 w_4660_n6791.n2555 9.3005
R18485 w_4660_n6791.n2558 w_4660_n6791.n2557 9.3005
R18486 w_4660_n6791.n200 w_4660_n6791.n199 9.3005
R18487 w_4660_n6791.n2563 w_4660_n6791.n2562 9.3005
R18488 w_4660_n6791.n2565 w_4660_n6791.n2564 9.3005
R18489 w_4660_n6791.n191 w_4660_n6791.n190 9.3005
R18490 w_4660_n6791.n2570 w_4660_n6791.n2569 9.3005
R18491 w_4660_n6791.n2571 w_4660_n6791.n187 9.3005
R18492 w_4660_n6791.n2573 w_4660_n6791.n2572 9.3005
R18493 w_4660_n6791.n185 w_4660_n6791.n184 9.3005
R18494 w_4660_n6791.n2577 w_4660_n6791.n28 9.3005
R18495 w_4660_n6791.n2579 w_4660_n6791.n2578 9.3005
R18496 w_4660_n6791.n181 w_4660_n6791.n180 9.3005
R18497 w_4660_n6791.n2584 w_4660_n6791.n2583 9.3005
R18498 w_4660_n6791.n2586 w_4660_n6791.n2585 9.3005
R18499 w_4660_n6791.n175 w_4660_n6791.n174 9.3005
R18500 w_4660_n6791.n2591 w_4660_n6791.n2590 9.3005
R18501 w_4660_n6791.n2593 w_4660_n6791.n2592 9.3005
R18502 w_4660_n6791.n169 w_4660_n6791.n168 9.3005
R18503 w_4660_n6791.n2598 w_4660_n6791.n2597 9.3005
R18504 w_4660_n6791.n2600 w_4660_n6791.n2599 9.3005
R18505 w_4660_n6791.n161 w_4660_n6791.n160 9.3005
R18506 w_4660_n6791.n2606 w_4660_n6791.n2605 9.3005
R18507 w_4660_n6791.n2607 w_4660_n6791.n153 9.3005
R18508 w_4660_n6791.n2611 w_4660_n6791.n2610 9.3005
R18509 w_4660_n6791.n2609 w_4660_n6791.n157 9.3005
R18510 w_4660_n6791.n2608 w_4660_n6791.n147 9.3005
R18511 w_4660_n6791.n1759 w_4660_n6791.n1758 9.3005
R18512 w_4660_n6791.n2617 w_4660_n6791.n2616 9.3005
R18513 w_4660_n6791.n2619 w_4660_n6791.n143 9.3005
R18514 w_4660_n6791.n2616 w_4660_n6791.n144 9.3005
R18515 w_4660_n6791.n2616 w_4660_n6791.n142 9.3005
R18516 w_4660_n6791.n2475 w_4660_n6791.n298 9.3005
R18517 w_4660_n6791.n2477 w_4660_n6791.n2476 9.3005
R18518 w_4660_n6791.n294 w_4660_n6791.n291 9.3005
R18519 w_4660_n6791.n2482 w_4660_n6791.n2481 9.3005
R18520 w_4660_n6791.n2483 w_4660_n6791.n290 9.3005
R18521 w_4660_n6791.n2485 w_4660_n6791.n2484 9.3005
R18522 w_4660_n6791.n285 w_4660_n6791.n282 9.3005
R18523 w_4660_n6791.n2490 w_4660_n6791.n2489 9.3005
R18524 w_4660_n6791.n2491 w_4660_n6791.n281 9.3005
R18525 w_4660_n6791.n2493 w_4660_n6791.n2492 9.3005
R18526 w_4660_n6791.n277 w_4660_n6791.n274 9.3005
R18527 w_4660_n6791.n2498 w_4660_n6791.n2497 9.3005
R18528 w_4660_n6791.n2499 w_4660_n6791.n273 9.3005
R18529 w_4660_n6791.n2501 w_4660_n6791.n2500 9.3005
R18530 w_4660_n6791.n269 w_4660_n6791.n266 9.3005
R18531 w_4660_n6791.n2506 w_4660_n6791.n2505 9.3005
R18532 w_4660_n6791.n2507 w_4660_n6791.n265 9.3005
R18533 w_4660_n6791.n2509 w_4660_n6791.n2508 9.3005
R18534 w_4660_n6791.n261 w_4660_n6791.n258 9.3005
R18535 w_4660_n6791.n2514 w_4660_n6791.n2513 9.3005
R18536 w_4660_n6791.n2515 w_4660_n6791.n251 9.3005
R18537 w_4660_n6791.n2517 w_4660_n6791.n2516 9.3005
R18538 w_4660_n6791.n257 w_4660_n6791.n249 9.3005
R18539 w_4660_n6791.n2473 w_4660_n6791.n301 9.3005
R18540 w_4660_n6791.n300 w_4660_n6791.n298 9.3005
R18541 w_4660_n6791.n2477 w_4660_n6791.n297 9.3005
R18542 w_4660_n6791.n296 w_4660_n6791.n294 9.3005
R18543 w_4660_n6791.n2481 w_4660_n6791.n293 9.3005
R18544 w_4660_n6791.n292 w_4660_n6791.n290 9.3005
R18545 w_4660_n6791.n2485 w_4660_n6791.n289 9.3005
R18546 w_4660_n6791.n288 w_4660_n6791.n285 9.3005
R18547 w_4660_n6791.n2489 w_4660_n6791.n284 9.3005
R18548 w_4660_n6791.n283 w_4660_n6791.n281 9.3005
R18549 w_4660_n6791.n2493 w_4660_n6791.n280 9.3005
R18550 w_4660_n6791.n279 w_4660_n6791.n277 9.3005
R18551 w_4660_n6791.n2497 w_4660_n6791.n276 9.3005
R18552 w_4660_n6791.n275 w_4660_n6791.n273 9.3005
R18553 w_4660_n6791.n2501 w_4660_n6791.n272 9.3005
R18554 w_4660_n6791.n271 w_4660_n6791.n269 9.3005
R18555 w_4660_n6791.n2505 w_4660_n6791.n268 9.3005
R18556 w_4660_n6791.n267 w_4660_n6791.n265 9.3005
R18557 w_4660_n6791.n2509 w_4660_n6791.n264 9.3005
R18558 w_4660_n6791.n263 w_4660_n6791.n261 9.3005
R18559 w_4660_n6791.n2513 w_4660_n6791.n260 9.3005
R18560 w_4660_n6791.n259 w_4660_n6791.n251 9.3005
R18561 w_4660_n6791.n2517 w_4660_n6791.n250 9.3005
R18562 w_4660_n6791.n252 w_4660_n6791.n249 9.3005
R18563 w_4660_n6791.n2518 w_4660_n6791.n2517 9.3005
R18564 w_4660_n6791.n2471 w_4660_n6791.n299 9.3005
R18565 w_4660_n6791.n2473 w_4660_n6791.n2472 9.3005
R18566 w_4660_n6791.n298 w_4660_n6791.n295 9.3005
R18567 w_4660_n6791.n2478 w_4660_n6791.n2477 9.3005
R18568 w_4660_n6791.n2479 w_4660_n6791.n294 9.3005
R18569 w_4660_n6791.n2481 w_4660_n6791.n2480 9.3005
R18570 w_4660_n6791.n290 w_4660_n6791.n287 9.3005
R18571 w_4660_n6791.n2486 w_4660_n6791.n2485 9.3005
R18572 w_4660_n6791.n2487 w_4660_n6791.n285 9.3005
R18573 w_4660_n6791.n2489 w_4660_n6791.n2488 9.3005
R18574 w_4660_n6791.n286 w_4660_n6791.n281 9.3005
R18575 w_4660_n6791.n2494 w_4660_n6791.n2493 9.3005
R18576 w_4660_n6791.n2495 w_4660_n6791.n277 9.3005
R18577 w_4660_n6791.n2497 w_4660_n6791.n2496 9.3005
R18578 w_4660_n6791.n273 w_4660_n6791.n270 9.3005
R18579 w_4660_n6791.n2502 w_4660_n6791.n2501 9.3005
R18580 w_4660_n6791.n2503 w_4660_n6791.n269 9.3005
R18581 w_4660_n6791.n2505 w_4660_n6791.n2504 9.3005
R18582 w_4660_n6791.n265 w_4660_n6791.n262 9.3005
R18583 w_4660_n6791.n2510 w_4660_n6791.n2509 9.3005
R18584 w_4660_n6791.n2511 w_4660_n6791.n261 9.3005
R18585 w_4660_n6791.n2513 w_4660_n6791.n2512 9.3005
R18586 w_4660_n6791.n251 w_4660_n6791.n248 9.3005
R18587 w_4660_n6791.n249 w_4660_n6791.n145 9.3005
R18588 w_4660_n6791.n2288 w_4660_n6791.n2284 9.3005
R18589 w_4660_n6791.n2291 w_4660_n6791.n2290 9.3005
R18590 w_4660_n6791.n2289 w_4660_n6791.n2278 9.3005
R18591 w_4660_n6791.n2296 w_4660_n6791.n2279 9.3005
R18592 w_4660_n6791.n2282 w_4660_n6791.n2281 9.3005
R18593 w_4660_n6791.n2280 w_4660_n6791.n422 9.3005
R18594 w_4660_n6791.n30 w_4660_n6791.n424 9.3005
R18595 w_4660_n6791.n423 w_4660_n6791.n29 9.3005
R18596 w_4660_n6791.n2305 w_4660_n6791.n420 9.3005
R18597 w_4660_n6791.n2307 w_4660_n6791.n2306 9.3005
R18598 w_4660_n6791.n2309 w_4660_n6791.n2308 9.3005
R18599 w_4660_n6791.n416 w_4660_n6791.n415 9.3005
R18600 w_4660_n6791.n2314 w_4660_n6791.n2313 9.3005
R18601 w_4660_n6791.n2315 w_4660_n6791.n414 9.3005
R18602 w_4660_n6791.n2318 w_4660_n6791.n2317 9.3005
R18603 w_4660_n6791.n2316 w_4660_n6791.n408 9.3005
R18604 w_4660_n6791.n2323 w_4660_n6791.n409 9.3005
R18605 w_4660_n6791.n412 w_4660_n6791.n411 9.3005
R18606 w_4660_n6791.n410 w_4660_n6791.n401 9.3005
R18607 w_4660_n6791.n2330 w_4660_n6791.n403 9.3005
R18608 w_4660_n6791.n402 w_4660_n6791.n399 9.3005
R18609 w_4660_n6791.n2334 w_4660_n6791.n398 9.3005
R18610 w_4660_n6791.n2336 w_4660_n6791.n2335 9.3005
R18611 w_4660_n6791.n2338 w_4660_n6791.n2337 9.3005
R18612 w_4660_n6791.n394 w_4660_n6791.n393 9.3005
R18613 w_4660_n6791.n2343 w_4660_n6791.n2342 9.3005
R18614 w_4660_n6791.n2344 w_4660_n6791.n392 9.3005
R18615 w_4660_n6791.n2347 w_4660_n6791.n2346 9.3005
R18616 w_4660_n6791.n2345 w_4660_n6791.n386 9.3005
R18617 w_4660_n6791.n31 w_4660_n6791.n387 9.3005
R18618 w_4660_n6791.n390 w_4660_n6791.n389 9.3005
R18619 w_4660_n6791.n388 w_4660_n6791.n379 9.3005
R18620 w_4660_n6791.n2359 w_4660_n6791.n381 9.3005
R18621 w_4660_n6791.n380 w_4660_n6791.n377 9.3005
R18622 w_4660_n6791.n2363 w_4660_n6791.n376 9.3005
R18623 w_4660_n6791.n2365 w_4660_n6791.n2364 9.3005
R18624 w_4660_n6791.n2367 w_4660_n6791.n2366 9.3005
R18625 w_4660_n6791.n372 w_4660_n6791.n371 9.3005
R18626 w_4660_n6791.n2372 w_4660_n6791.n2371 9.3005
R18627 w_4660_n6791.n2373 w_4660_n6791.n370 9.3005
R18628 w_4660_n6791.n2375 w_4660_n6791.n2374 9.3005
R18629 w_4660_n6791.n367 w_4660_n6791.n366 9.3005
R18630 w_4660_n6791.n2381 w_4660_n6791.n2380 9.3005
R18631 w_4660_n6791.n2382 w_4660_n6791.n365 9.3005
R18632 w_4660_n6791.n2385 w_4660_n6791.n2384 9.3005
R18633 w_4660_n6791.n2383 w_4660_n6791.n361 9.3005
R18634 w_4660_n6791.n2389 w_4660_n6791.n363 9.3005
R18635 w_4660_n6791.n362 w_4660_n6791.n354 9.3005
R18636 w_4660_n6791.n2398 w_4660_n6791.n356 9.3005
R18637 w_4660_n6791.n355 w_4660_n6791.n352 9.3005
R18638 w_4660_n6791.n2402 w_4660_n6791.n351 9.3005
R18639 w_4660_n6791.n2404 w_4660_n6791.n2403 9.3005
R18640 w_4660_n6791.n2407 w_4660_n6791.n2406 9.3005
R18641 w_4660_n6791.n2405 w_4660_n6791.n348 9.3005
R18642 w_4660_n6791.n2411 w_4660_n6791.n347 9.3005
R18643 w_4660_n6791.n2413 w_4660_n6791.n2412 9.3005
R18644 w_4660_n6791.n2415 w_4660_n6791.n2414 9.3005
R18645 w_4660_n6791.n343 w_4660_n6791.n342 9.3005
R18646 w_4660_n6791.n2420 w_4660_n6791.n2419 9.3005
R18647 w_4660_n6791.n2421 w_4660_n6791.n341 9.3005
R18648 w_4660_n6791.n2424 w_4660_n6791.n2423 9.3005
R18649 w_4660_n6791.n2422 w_4660_n6791.n335 9.3005
R18650 w_4660_n6791.n2429 w_4660_n6791.n336 9.3005
R18651 w_4660_n6791.n339 w_4660_n6791.n338 9.3005
R18652 w_4660_n6791.n337 w_4660_n6791.n328 9.3005
R18653 w_4660_n6791.n33 w_4660_n6791.n330 9.3005
R18654 w_4660_n6791.n329 w_4660_n6791.n32 9.3005
R18655 w_4660_n6791.n2438 w_4660_n6791.n326 9.3005
R18656 w_4660_n6791.n2440 w_4660_n6791.n2439 9.3005
R18657 w_4660_n6791.n2442 w_4660_n6791.n2441 9.3005
R18658 w_4660_n6791.n322 w_4660_n6791.n321 9.3005
R18659 w_4660_n6791.n2447 w_4660_n6791.n2446 9.3005
R18660 w_4660_n6791.n2448 w_4660_n6791.n320 9.3005
R18661 w_4660_n6791.n2451 w_4660_n6791.n2450 9.3005
R18662 w_4660_n6791.n2449 w_4660_n6791.n314 9.3005
R18663 w_4660_n6791.n2456 w_4660_n6791.n315 9.3005
R18664 w_4660_n6791.n318 w_4660_n6791.n317 9.3005
R18665 w_4660_n6791.n316 w_4660_n6791.n307 9.3005
R18666 w_4660_n6791.n2462 w_4660_n6791.n309 9.3005
R18667 w_4660_n6791.n308 w_4660_n6791.n305 9.3005
R18668 w_4660_n6791.n2466 w_4660_n6791.n304 9.3005
R18669 w_4660_n6791.n2468 w_4660_n6791.n2467 9.3005
R18670 w_4660_n6791.n2284 w_4660_n6791.n2283 9.3005
R18671 w_4660_n6791.n2292 w_4660_n6791.n2291 9.3005
R18672 w_4660_n6791.n2293 w_4660_n6791.n2278 9.3005
R18673 w_4660_n6791.n2296 w_4660_n6791.n2295 9.3005
R18674 w_4660_n6791.n2294 w_4660_n6791.n2282 9.3005
R18675 w_4660_n6791.n422 w_4660_n6791.n421 9.3005
R18676 w_4660_n6791.n2302 w_4660_n6791.n30 9.3005
R18677 w_4660_n6791.n2303 w_4660_n6791.n29 9.3005
R18678 w_4660_n6791.n2305 w_4660_n6791.n2304 9.3005
R18679 w_4660_n6791.n2306 w_4660_n6791.n418 9.3005
R18680 w_4660_n6791.n2310 w_4660_n6791.n2309 9.3005
R18681 w_4660_n6791.n2311 w_4660_n6791.n416 9.3005
R18682 w_4660_n6791.n2313 w_4660_n6791.n2312 9.3005
R18683 w_4660_n6791.n414 w_4660_n6791.n413 9.3005
R18684 w_4660_n6791.n2319 w_4660_n6791.n2318 9.3005
R18685 w_4660_n6791.n2320 w_4660_n6791.n408 9.3005
R18686 w_4660_n6791.n2323 w_4660_n6791.n2322 9.3005
R18687 w_4660_n6791.n2321 w_4660_n6791.n412 9.3005
R18688 w_4660_n6791.n401 w_4660_n6791.n400 9.3005
R18689 w_4660_n6791.n2331 w_4660_n6791.n2330 9.3005
R18690 w_4660_n6791.n2332 w_4660_n6791.n399 9.3005
R18691 w_4660_n6791.n2334 w_4660_n6791.n2333 9.3005
R18692 w_4660_n6791.n2335 w_4660_n6791.n396 9.3005
R18693 w_4660_n6791.n2339 w_4660_n6791.n2338 9.3005
R18694 w_4660_n6791.n2340 w_4660_n6791.n394 9.3005
R18695 w_4660_n6791.n2342 w_4660_n6791.n2341 9.3005
R18696 w_4660_n6791.n392 w_4660_n6791.n391 9.3005
R18697 w_4660_n6791.n2348 w_4660_n6791.n2347 9.3005
R18698 w_4660_n6791.n2349 w_4660_n6791.n386 9.3005
R18699 w_4660_n6791.n31 w_4660_n6791.n2351 9.3005
R18700 w_4660_n6791.n2350 w_4660_n6791.n390 9.3005
R18701 w_4660_n6791.n379 w_4660_n6791.n378 9.3005
R18702 w_4660_n6791.n2360 w_4660_n6791.n2359 9.3005
R18703 w_4660_n6791.n2361 w_4660_n6791.n377 9.3005
R18704 w_4660_n6791.n2363 w_4660_n6791.n2362 9.3005
R18705 w_4660_n6791.n2364 w_4660_n6791.n374 9.3005
R18706 w_4660_n6791.n2368 w_4660_n6791.n2367 9.3005
R18707 w_4660_n6791.n2369 w_4660_n6791.n372 9.3005
R18708 w_4660_n6791.n2371 w_4660_n6791.n2370 9.3005
R18709 w_4660_n6791.n370 w_4660_n6791.n369 9.3005
R18710 w_4660_n6791.n2376 w_4660_n6791.n2375 9.3005
R18711 w_4660_n6791.n2378 w_4660_n6791.n367 9.3005
R18712 w_4660_n6791.n2380 w_4660_n6791.n2379 9.3005
R18713 w_4660_n6791.n365 w_4660_n6791.n364 9.3005
R18714 w_4660_n6791.n2386 w_4660_n6791.n2385 9.3005
R18715 w_4660_n6791.n2387 w_4660_n6791.n361 9.3005
R18716 w_4660_n6791.n2389 w_4660_n6791.n2388 9.3005
R18717 w_4660_n6791.n354 w_4660_n6791.n353 9.3005
R18718 w_4660_n6791.n2399 w_4660_n6791.n2398 9.3005
R18719 w_4660_n6791.n2400 w_4660_n6791.n352 9.3005
R18720 w_4660_n6791.n2402 w_4660_n6791.n2401 9.3005
R18721 w_4660_n6791.n2403 w_4660_n6791.n349 9.3005
R18722 w_4660_n6791.n2408 w_4660_n6791.n2407 9.3005
R18723 w_4660_n6791.n2409 w_4660_n6791.n348 9.3005
R18724 w_4660_n6791.n2411 w_4660_n6791.n2410 9.3005
R18725 w_4660_n6791.n2412 w_4660_n6791.n345 9.3005
R18726 w_4660_n6791.n2416 w_4660_n6791.n2415 9.3005
R18727 w_4660_n6791.n2417 w_4660_n6791.n343 9.3005
R18728 w_4660_n6791.n2419 w_4660_n6791.n2418 9.3005
R18729 w_4660_n6791.n341 w_4660_n6791.n340 9.3005
R18730 w_4660_n6791.n2425 w_4660_n6791.n2424 9.3005
R18731 w_4660_n6791.n2426 w_4660_n6791.n335 9.3005
R18732 w_4660_n6791.n2429 w_4660_n6791.n2428 9.3005
R18733 w_4660_n6791.n2427 w_4660_n6791.n339 9.3005
R18734 w_4660_n6791.n328 w_4660_n6791.n327 9.3005
R18735 w_4660_n6791.n2435 w_4660_n6791.n33 9.3005
R18736 w_4660_n6791.n2436 w_4660_n6791.n32 9.3005
R18737 w_4660_n6791.n2438 w_4660_n6791.n2437 9.3005
R18738 w_4660_n6791.n2439 w_4660_n6791.n324 9.3005
R18739 w_4660_n6791.n2443 w_4660_n6791.n2442 9.3005
R18740 w_4660_n6791.n2444 w_4660_n6791.n322 9.3005
R18741 w_4660_n6791.n2446 w_4660_n6791.n2445 9.3005
R18742 w_4660_n6791.n320 w_4660_n6791.n319 9.3005
R18743 w_4660_n6791.n2452 w_4660_n6791.n2451 9.3005
R18744 w_4660_n6791.n2453 w_4660_n6791.n314 9.3005
R18745 w_4660_n6791.n2456 w_4660_n6791.n2455 9.3005
R18746 w_4660_n6791.n2454 w_4660_n6791.n318 9.3005
R18747 w_4660_n6791.n307 w_4660_n6791.n306 9.3005
R18748 w_4660_n6791.n2463 w_4660_n6791.n2462 9.3005
R18749 w_4660_n6791.n2464 w_4660_n6791.n305 9.3005
R18750 w_4660_n6791.n2466 w_4660_n6791.n2465 9.3005
R18751 w_4660_n6791.n2467 w_4660_n6791.n302 9.3005
R18752 w_4660_n6791.n2470 w_4660_n6791.n2469 9.3005
R18753 w_4660_n6791.n1519 w_4660_n6791.n453 9.22941
R18754 w_4660_n6791.n989 w_4660_n6791.n938 8.79188
R18755 w_4660_n6791.n2651 w_4660_n6791.n109 8.41193
R18756 w_4660_n6791.n2622 w_4660_n6791.n2621 7.79915
R18757 w_4660_n6791.n278 w_4660_n6791.n113 7.70883
R18758 w_4660_n6791.n2649 w_4660_n6791.n113 7.70883
R18759 w_4660_n6791.n247 w_4660_n6791.n246 7.70883
R18760 w_4660_n6791.n1762 w_4660_n6791.n246 7.70883
R18761 w_4660_n6791.n2648 w_4660_n6791.n2647 7.70883
R18762 w_4660_n6791.n2649 w_4660_n6791.n2648 7.70883
R18763 w_4660_n6791.n1761 w_4660_n6791.n1760 7.70883
R18764 w_4660_n6791.n1762 w_4660_n6791.n1761 7.70883
R18765 w_4660_n6791.n1447 w_4660_n6791.n112 7.70883
R18766 w_4660_n6791.n2649 w_4660_n6791.n112 7.70883
R18767 w_4660_n6791.n936 w_4660_n6791.n452 7.70883
R18768 w_4660_n6791.n1762 w_4660_n6791.n452 7.70883
R18769 w_4660_n6791.n2651 w_4660_n6791.n2650 7.70883
R18770 w_4660_n6791.n2650 w_4660_n6791.n2649 7.70883
R18771 w_4660_n6791.n1764 w_4660_n6791.n1763 7.70883
R18772 w_4660_n6791.n1763 w_4660_n6791.n1762 7.70883
R18773 w_4660_n6791.n767 w_4660_n6791.n766 7.49675
R18774 w_4660_n6791.n2522 w_4660_n6791.t79 6.70505
R18775 w_4660_n6791.n2522 w_4660_n6791.t43 6.70505
R18776 w_4660_n6791.n2621 w_4660_n6791.n2620 5.23915
R18777 w_4660_n6791.n2519 w_4660_n6791.n2518 4.75479
R18778 w_4660_n6791.n767 w_4660_n6791.n761 4.48498
R18779 w_4660_n6791.n990 w_4660_n6791.n989 4.27423
R18780 w_4660_n6791.n2522 w_4660_n6791.n245 4.20505
R18781 w_4660_n6791.n2522 w_4660_n6791.n241 4.20505
R18782 w_4660_n6791.n2522 w_4660_n6791.n240 4.20505
R18783 w_4660_n6791.n2522 w_4660_n6791.n237 4.20505
R18784 w_4660_n6791.n2522 w_4660_n6791.n236 4.20505
R18785 w_4660_n6791.n2522 w_4660_n6791.n235 4.20505
R18786 w_4660_n6791.n2523 w_4660_n6791.n2522 4.20505
R18787 w_4660_n6791.n2522 w_4660_n6791.n243 4.20505
R18788 w_4660_n6791.n1447 w_4660_n6791.n1446 4.02336
R18789 w_4660_n6791.n2272 w_4660_n6791.n2271 3.4105
R18790 w_4660_n6791.n40 w_4660_n6791.n445 3.4105
R18791 w_4660_n6791.n2273 w_4660_n6791.n433 3.4105
R18792 w_4660_n6791.n2273 w_4660_n6791.n435 3.4105
R18793 w_4660_n6791.n2273 w_4660_n6791.n432 3.4105
R18794 w_4660_n6791.n2273 w_4660_n6791.n436 3.4105
R18795 w_4660_n6791.n2273 w_4660_n6791.n431 3.4105
R18796 w_4660_n6791.n2273 w_4660_n6791.n437 3.4105
R18797 w_4660_n6791.n2273 w_4660_n6791.n430 3.4105
R18798 w_4660_n6791.n2273 w_4660_n6791.n2272 3.4105
R18799 w_4660_n6791.n1422 w_4660_n6791.n1421 3.29193
R18800 w_4660_n6791.n2619 w_4660_n6791.n2618 3.01226
R18801 w_4660_n6791.n2494 w_4660_n6791.n278 2.5605
R18802 w_4660_n6791.n989 w_4660_n6791.n988 2.51438
R18803 w_4660_n6791.n768 w_4660_n6791.n767 2.40901
R18804 w_4660_n6791.n2377 w_4660_n6791.n244 2.10277
R18805 w_4660_n6791.n2522 w_4660_n6791.n244 2.10277
R18806 w_4660_n6791.n2521 w_4660_n6791.n2520 2.10277
R18807 w_4660_n6791.n2522 w_4660_n6791.n2521 2.10277
R18808 w_4660_n6791.n1605 w_4660_n6791.n115 2.10277
R18809 w_4660_n6791.n2522 w_4660_n6791.n115 2.10277
R18810 w_4660_n6791.n1520 w_4660_n6791.n114 2.10277
R18811 w_4660_n6791.n2522 w_4660_n6791.n114 2.10277
R18812 w_4660_n6791.n596 w_4660_n6791.n239 2.10277
R18813 w_4660_n6791.n2522 w_4660_n6791.n239 2.10277
R18814 w_4660_n6791.n937 w_4660_n6791.n238 2.10277
R18815 w_4660_n6791.n2522 w_4660_n6791.n238 2.10277
R18816 w_4660_n6791.n1314 w_4660_n6791.n111 2.10277
R18817 w_4660_n6791.n2522 w_4660_n6791.n111 2.10277
R18818 w_4660_n6791.n2184 w_4660_n6791.n110 2.10277
R18819 w_4660_n6791.n2522 w_4660_n6791.n110 2.10277
R18820 w_4660_n6791.n2621 w_4660_n6791.n143 2.03192
R18821 w_4660_n6791.n40 w_4660_n6791.n444 1.70267
R18822 w_4660_n6791.n2271 w_4660_n6791.n441 1.70263
R18823 w_4660_n6791.n2271 w_4660_n6791.n440 1.70263
R18824 w_4660_n6791.n2271 w_4660_n6791.n439 1.70263
R18825 w_4660_n6791.n2271 w_4660_n6791.n438 1.70263
R18826 w_4660_n6791.n40 w_4660_n6791.n443 1.70263
R18827 w_4660_n6791.n40 w_4660_n6791.n442 1.70263
R18828 w_4660_n6791.n40 w_4660_n6791.n39 1.70263
R18829 w_4660_n6791.n2273 w_4660_n6791.n434 1.70263
R18830 w_4660_n6791.n2270 w_4660_n6791.n2269 1.7018
R18831 w_4660_n6791.n2287 w_4660_n6791.n2286 1.42902
R18832 w_4660_n6791.n2701 w_4660_n6791.n41 1.13717
R18833 w_4660_n6791.n2700 w_4660_n6791.n2699 1.13717
R18834 w_4660_n6791.n2698 w_4660_n6791.n44 1.13717
R18835 w_4660_n6791.n2108 w_4660_n6791.n46 1.13717
R18836 w_4660_n6791.n2110 w_4660_n6791.n2109 1.13717
R18837 w_4660_n6791.n2107 w_4660_n6791.n1922 1.13717
R18838 w_4660_n6791.n2106 w_4660_n6791.n2105 1.13717
R18839 w_4660_n6791.n2104 w_4660_n6791.n1923 1.13717
R18840 w_4660_n6791.n2102 w_4660_n6791.n2101 1.13717
R18841 w_4660_n6791.n2100 w_4660_n6791.n1925 1.13717
R18842 w_4660_n6791.n2099 w_4660_n6791.n2098 1.13717
R18843 w_4660_n6791.n2096 w_4660_n6791.n1926 1.13717
R18844 w_4660_n6791.n2095 w_4660_n6791.n2094 1.13717
R18845 w_4660_n6791.n2093 w_4660_n6791.n1928 1.13717
R18846 w_4660_n6791.n2092 w_4660_n6791.n2091 1.13717
R18847 w_4660_n6791.n2088 w_4660_n6791.n1929 1.13717
R18848 w_4660_n6791.n2087 w_4660_n6791.n2086 1.13717
R18849 w_4660_n6791.n2085 w_4660_n6791.n2084 1.13717
R18850 w_4660_n6791.n2083 w_4660_n6791.n1932 1.13717
R18851 w_4660_n6791.n2082 w_4660_n6791.n2081 1.13717
R18852 w_4660_n6791.n2078 w_4660_n6791.n3 1.13717
R18853 w_4660_n6791.n2080 w_4660_n6791.n2079 1.13717
R18854 w_4660_n6791.n37 w_4660_n6791.n4 1.13717
R18855 w_4660_n6791.n2076 w_4660_n6791.n2075 1.13717
R18856 w_4660_n6791.n2074 w_4660_n6791.n1936 1.13717
R18857 w_4660_n6791.n2072 w_4660_n6791.n2071 1.13717
R18858 w_4660_n6791.n2068 w_4660_n6791.n1938 1.13717
R18859 w_4660_n6791.n2067 w_4660_n6791.n2066 1.13717
R18860 w_4660_n6791.n2064 w_4660_n6791.n2063 1.13717
R18861 w_4660_n6791.n2062 w_4660_n6791.n1942 1.13717
R18862 w_4660_n6791.n2061 w_4660_n6791.n2060 1.13717
R18863 w_4660_n6791.n2058 w_4660_n6791.n2057 1.13717
R18864 w_4660_n6791.n2056 w_4660_n6791.n1946 1.13717
R18865 w_4660_n6791.n2055 w_4660_n6791.n2054 1.13717
R18866 w_4660_n6791.n2052 w_4660_n6791.n2051 1.13717
R18867 w_4660_n6791.n2050 w_4660_n6791.n1950 1.13717
R18868 w_4660_n6791.n2049 w_4660_n6791.n2048 1.13717
R18869 w_4660_n6791.n2046 w_4660_n6791.n2045 1.13717
R18870 w_4660_n6791.n2044 w_4660_n6791.n1954 1.13717
R18871 w_4660_n6791.n2043 w_4660_n6791.n2042 1.13717
R18872 w_4660_n6791.n2040 w_4660_n6791.n2039 1.13717
R18873 w_4660_n6791.n2038 w_4660_n6791.n1958 1.13717
R18874 w_4660_n6791.n2037 w_4660_n6791.n2036 1.13717
R18875 w_4660_n6791.n2034 w_4660_n6791.n2033 1.13717
R18876 w_4660_n6791.n2032 w_4660_n6791.n1961 1.13717
R18877 w_4660_n6791.n2031 w_4660_n6791.n2030 1.13717
R18878 w_4660_n6791.n2028 w_4660_n6791.n1962 1.13717
R18879 w_4660_n6791.n2027 w_4660_n6791.n2026 1.13717
R18880 w_4660_n6791.n2023 w_4660_n6791.n1964 1.13717
R18881 w_4660_n6791.n2022 w_4660_n6791.n2021 1.13717
R18882 w_4660_n6791.n2018 w_4660_n6791.n2017 1.13717
R18883 w_4660_n6791.n2016 w_4660_n6791.n1967 1.13717
R18884 w_4660_n6791.n2011 w_4660_n6791.n2010 1.13717
R18885 w_4660_n6791.n2015 w_4660_n6791.n2014 1.13717
R18886 w_4660_n6791.n2009 w_4660_n6791.n1971 1.13717
R18887 w_4660_n6791.n2008 w_4660_n6791.n2007 1.13717
R18888 w_4660_n6791.n2006 w_4660_n6791.n2005 1.13717
R18889 w_4660_n6791.n2004 w_4660_n6791.n2003 1.13717
R18890 w_4660_n6791.n2002 w_4660_n6791.n1976 1.13717
R18891 w_4660_n6791.n2001 w_4660_n6791.n2000 1.13717
R18892 w_4660_n6791.n1997 w_4660_n6791.n1996 1.13717
R18893 w_4660_n6791.n1995 w_4660_n6791.n0 1.13717
R18894 w_4660_n6791.n1994 w_4660_n6791.n1993 1.13717
R18895 w_4660_n6791.n1991 w_4660_n6791.n1990 1.13717
R18896 w_4660_n6791.n1989 w_4660_n6791.n38 1.13717
R18897 w_4660_n6791.n1988 w_4660_n6791.n1987 1.13717
R18898 w_4660_n6791.n1985 w_4660_n6791.n1984 1.13717
R18899 w_4660_n6791.n1983 w_4660_n6791.n35 1.13717
R18900 w_4660_n6791.n446 w_4660_n6791.n34 1.13717
R18901 w_4660_n6791.n2268 w_4660_n6791.n2267 1.13717
R18902 w_4660_n6791.n1217 w_4660_n6791.n429 1.1255
R18903 w_4660_n6791.n1215 w_4660_n6791.n1214 1.1255
R18904 w_4660_n6791.n1213 w_4660_n6791.n1130 1.1255
R18905 w_4660_n6791.n1212 w_4660_n6791.n1124 1.1255
R18906 w_4660_n6791.n1211 w_4660_n6791.n1118 1.1255
R18907 w_4660_n6791.n1210 w_4660_n6791.n12 1.1255
R18908 w_4660_n6791.n1209 w_4660_n6791.n1106 1.1255
R18909 w_4660_n6791.n1208 w_4660_n6791.n1100 1.1255
R18910 w_4660_n6791.n1207 w_4660_n6791.n1098 1.1255
R18911 w_4660_n6791.n1206 w_4660_n6791.n1086 1.1255
R18912 w_4660_n6791.n1205 w_4660_n6791.n1080 1.1255
R18913 w_4660_n6791.n1204 w_4660_n6791.n1074 1.1255
R18914 w_4660_n6791.n1203 w_4660_n6791.n1068 1.1255
R18915 w_4660_n6791.n1202 w_4660_n6791.n1062 1.1255
R18916 w_4660_n6791.n1201 w_4660_n6791.n1056 1.1255
R18917 w_4660_n6791.n1200 w_4660_n6791.n1054 1.1255
R18918 w_4660_n6791.n1199 w_4660_n6791.n14 1.1255
R18919 w_4660_n6791.n1198 w_4660_n6791.n1038 1.1255
R18920 w_4660_n6791.n1197 w_4660_n6791.n1032 1.1255
R18921 w_4660_n6791.n1196 w_4660_n6791.n1030 1.1255
R18922 w_4660_n6791.n1195 w_4660_n6791.n1018 1.1255
R18923 w_4660_n6791.n1194 w_4660_n6791.n1012 1.1255
R18924 w_4660_n6791.n1193 w_4660_n6791.n1006 1.1255
R18925 w_4660_n6791.n1192 w_4660_n6791.n16 1.1255
R18926 w_4660_n6791.n1191 w_4660_n6791.n995 1.1255
R18927 w_4660_n6791.n1190 w_4660_n6791.n987 1.1255
R18928 w_4660_n6791.n505 w_4660_n6791.n428 1.1255
R18929 w_4660_n6791.n735 w_4660_n6791.n511 1.1255
R18930 w_4660_n6791.n736 w_4660_n6791.n521 1.1255
R18931 w_4660_n6791.n737 w_4660_n6791.n528 1.1255
R18932 w_4660_n6791.n738 w_4660_n6791.n534 1.1255
R18933 w_4660_n6791.n739 w_4660_n6791.n18 1.1255
R18934 w_4660_n6791.n740 w_4660_n6791.n548 1.1255
R18935 w_4660_n6791.n741 w_4660_n6791.n555 1.1255
R18936 w_4660_n6791.n742 w_4660_n6791.n563 1.1255
R18937 w_4660_n6791.n743 w_4660_n6791.n571 1.1255
R18938 w_4660_n6791.n744 w_4660_n6791.n578 1.1255
R18939 w_4660_n6791.n745 w_4660_n6791.n586 1.1255
R18940 w_4660_n6791.n746 w_4660_n6791.n592 1.1255
R18941 w_4660_n6791.n747 w_4660_n6791.n601 1.1255
R18942 w_4660_n6791.n748 w_4660_n6791.n609 1.1255
R18943 w_4660_n6791.n749 w_4660_n6791.n615 1.1255
R18944 w_4660_n6791.n750 w_4660_n6791.n20 1.1255
R18945 w_4660_n6791.n751 w_4660_n6791.n629 1.1255
R18946 w_4660_n6791.n752 w_4660_n6791.n635 1.1255
R18947 w_4660_n6791.n753 w_4660_n6791.n643 1.1255
R18948 w_4660_n6791.n754 w_4660_n6791.n651 1.1255
R18949 w_4660_n6791.n755 w_4660_n6791.n658 1.1255
R18950 w_4660_n6791.n756 w_4660_n6791.n666 1.1255
R18951 w_4660_n6791.n757 w_4660_n6791.n22 1.1255
R18952 w_4660_n6791.n758 w_4660_n6791.n680 1.1255
R18953 w_4660_n6791.n760 w_4660_n6791.n759 1.1255
R18954 w_4660_n6791.n1523 w_4660_n6791.n427 1.1255
R18955 w_4660_n6791.n1631 w_4660_n6791.n1528 1.1255
R18956 w_4660_n6791.n1632 w_4660_n6791.n24 1.1255
R18957 w_4660_n6791.n1633 w_4660_n6791.n1542 1.1255
R18958 w_4660_n6791.n1634 w_4660_n6791.n1548 1.1255
R18959 w_4660_n6791.n1635 w_4660_n6791.n1556 1.1255
R18960 w_4660_n6791.n1636 w_4660_n6791.n1564 1.1255
R18961 w_4660_n6791.n1637 w_4660_n6791.n1571 1.1255
R18962 w_4660_n6791.n1638 w_4660_n6791.n1579 1.1255
R18963 w_4660_n6791.n1639 w_4660_n6791.n26 1.1255
R18964 w_4660_n6791.n1640 w_4660_n6791.n1593 1.1255
R18965 w_4660_n6791.n1641 w_4660_n6791.n1600 1.1255
R18966 w_4660_n6791.n1673 w_4660_n6791.n1672 1.1255
R18967 w_4660_n6791.n1671 w_4660_n6791.n229 1.1255
R18968 w_4660_n6791.n1670 w_4660_n6791.n223 1.1255
R18969 w_4660_n6791.n1669 w_4660_n6791.n217 1.1255
R18970 w_4660_n6791.n1668 w_4660_n6791.n215 1.1255
R18971 w_4660_n6791.n1667 w_4660_n6791.n202 1.1255
R18972 w_4660_n6791.n1666 w_4660_n6791.n196 1.1255
R18973 w_4660_n6791.n1665 w_4660_n6791.n194 1.1255
R18974 w_4660_n6791.n1664 w_4660_n6791.n28 1.1255
R18975 w_4660_n6791.n1663 w_4660_n6791.n177 1.1255
R18976 w_4660_n6791.n1662 w_4660_n6791.n171 1.1255
R18977 w_4660_n6791.n165 w_4660_n6791.n152 1.1255
R18978 w_4660_n6791.n2613 w_4660_n6791.n2612 1.1255
R18979 w_4660_n6791.n2615 w_4660_n6791.n2614 1.1255
R18980 w_4660_n6791.n2285 w_4660_n6791.n2277 1.1255
R18981 w_4660_n6791.n2298 w_4660_n6791.n2297 1.1255
R18982 w_4660_n6791.n30 w_4660_n6791.n2301 1.1255
R18983 w_4660_n6791.n2300 w_4660_n6791.n419 1.1255
R18984 w_4660_n6791.n417 w_4660_n6791.n407 1.1255
R18985 w_4660_n6791.n2325 w_4660_n6791.n2324 1.1255
R18986 w_4660_n6791.n2329 w_4660_n6791.n2328 1.1255
R18987 w_4660_n6791.n2327 w_4660_n6791.n397 1.1255
R18988 w_4660_n6791.n395 w_4660_n6791.n385 1.1255
R18989 w_4660_n6791.n2352 w_4660_n6791.n31 1.1255
R18990 w_4660_n6791.n2358 w_4660_n6791.n2357 1.1255
R18991 w_4660_n6791.n2356 w_4660_n6791.n375 1.1255
R18992 w_4660_n6791.n2355 w_4660_n6791.n373 1.1255
R18993 w_4660_n6791.n368 w_4660_n6791.n360 1.1255
R18994 w_4660_n6791.n2391 w_4660_n6791.n2390 1.1255
R18995 w_4660_n6791.n2397 w_4660_n6791.n2396 1.1255
R18996 w_4660_n6791.n2395 w_4660_n6791.n350 1.1255
R18997 w_4660_n6791.n2394 w_4660_n6791.n346 1.1255
R18998 w_4660_n6791.n344 w_4660_n6791.n334 1.1255
R18999 w_4660_n6791.n2431 w_4660_n6791.n2430 1.1255
R19000 w_4660_n6791.n33 w_4660_n6791.n2434 1.1255
R19001 w_4660_n6791.n2433 w_4660_n6791.n325 1.1255
R19002 w_4660_n6791.n323 w_4660_n6791.n313 1.1255
R19003 w_4660_n6791.n2458 w_4660_n6791.n2457 1.1255
R19004 w_4660_n6791.n2461 w_4660_n6791.n2460 1.1255
R19005 w_4660_n6791.n2459 w_4660_n6791.n303 1.1255
R19006 w_4660_n6791.n2266 w_4660_n6791.n2265 1.1255
R19007 w_4660_n6791.n1982 w_4660_n6791.n1769 1.1255
R19008 w_4660_n6791.n1980 w_4660_n6791.n6 1.1255
R19009 w_4660_n6791.n1978 w_4660_n6791.n1783 1.1255
R19010 w_4660_n6791.n1975 w_4660_n6791.n1791 1.1255
R19011 w_4660_n6791.n1971 w_4660_n6791.n1797 1.1255
R19012 w_4660_n6791.n2013 w_4660_n6791.n1807 1.1255
R19013 w_4660_n6791.n2020 w_4660_n6791.n1814 1.1255
R19014 w_4660_n6791.n2029 w_4660_n6791.n1820 1.1255
R19015 w_4660_n6791.n2035 w_4660_n6791.n8 1.1255
R19016 w_4660_n6791.n2041 w_4660_n6791.n1834 1.1255
R19017 w_4660_n6791.n2047 w_4660_n6791.n1841 1.1255
R19018 w_4660_n6791.n2053 w_4660_n6791.n1849 1.1255
R19019 w_4660_n6791.n2059 w_4660_n6791.n1857 1.1255
R19020 w_4660_n6791.n2065 w_4660_n6791.n1864 1.1255
R19021 w_4660_n6791.n2073 w_4660_n6791.n1872 1.1255
R19022 w_4660_n6791.n37 w_4660_n6791.n36 1.1255
R19023 w_4660_n6791.n1934 w_4660_n6791.n1887 1.1255
R19024 w_4660_n6791.n1931 w_4660_n6791.n1894 1.1255
R19025 w_4660_n6791.n2090 w_4660_n6791.n1900 1.1255
R19026 w_4660_n6791.n2097 w_4660_n6791.n10 1.1255
R19027 w_4660_n6791.n2103 w_4660_n6791.n1914 1.1255
R19028 w_4660_n6791.n2112 w_4660_n6791.n2111 1.1255
R19029 w_4660_n6791.n2697 w_4660_n6791.n2696 1.1255
R19030 w_4660_n6791.n2703 w_4660_n6791.n42 1.1255
R19031 w_4660_n6791.n64 w_4660_n6791.n43 1.1255
R19032 w_4660_n6791.n1413 w_4660_n6791.n985 1.09764
R19033 w_4660_n6791.n1417 w_4660_n6791.n939 0.444266
R19034 w_4660_n6791.n254 w_4660_n6791.n253 0.444266
R19035 w_4660_n6791.n944 w_4660_n6791.n939 0.402766
R19036 w_4660_n6791.n256 w_4660_n6791.n254 0.402766
R19037 w_4660_n6791.n2277 w_4660_n6791.n2276 0.377474
R19038 w_4660_n6791.n2276 w_4660_n6791.n2275 0.332861
R19039 w_4660_n6791.n2275 w_4660_n6791.n2274 0.332698
R19040 w_4660_n6791.n2274 w_4660_n6791.n2273 0.301732
R19041 w_4660_n6791.n2702 w_4660_n6791.n2701 0.291623
R19042 w_4660_n6791.n1475 w_4660_n6791.n458 0.12796
R19043 w_4660_n6791.n1631 w_4660_n6791.n427 0.1185
R19044 w_4660_n6791.n1632 w_4660_n6791.n1631 0.1185
R19045 w_4660_n6791.n1633 w_4660_n6791.n1632 0.1185
R19046 w_4660_n6791.n1634 w_4660_n6791.n1633 0.1185
R19047 w_4660_n6791.n1635 w_4660_n6791.n1634 0.1185
R19048 w_4660_n6791.n1636 w_4660_n6791.n1635 0.1185
R19049 w_4660_n6791.n1637 w_4660_n6791.n1636 0.1185
R19050 w_4660_n6791.n1638 w_4660_n6791.n1637 0.1185
R19051 w_4660_n6791.n1639 w_4660_n6791.n1638 0.1185
R19052 w_4660_n6791.n1640 w_4660_n6791.n1639 0.1185
R19053 w_4660_n6791.n1641 w_4660_n6791.n1640 0.1185
R19054 w_4660_n6791.n1672 w_4660_n6791.n1641 0.1185
R19055 w_4660_n6791.n1672 w_4660_n6791.n1671 0.1185
R19056 w_4660_n6791.n1671 w_4660_n6791.n1670 0.1185
R19057 w_4660_n6791.n1670 w_4660_n6791.n1669 0.1185
R19058 w_4660_n6791.n1669 w_4660_n6791.n1668 0.1185
R19059 w_4660_n6791.n1668 w_4660_n6791.n1667 0.1185
R19060 w_4660_n6791.n1667 w_4660_n6791.n1666 0.1185
R19061 w_4660_n6791.n1666 w_4660_n6791.n1665 0.1185
R19062 w_4660_n6791.n1665 w_4660_n6791.n1664 0.1185
R19063 w_4660_n6791.n1664 w_4660_n6791.n1663 0.1185
R19064 w_4660_n6791.n1663 w_4660_n6791.n1662 0.1185
R19065 w_4660_n6791.n1662 w_4660_n6791.n152 0.1185
R19066 w_4660_n6791.n2613 w_4660_n6791.n152 0.1185
R19067 w_4660_n6791.n2614 w_4660_n6791.n2613 0.1185
R19068 w_4660_n6791.n735 w_4660_n6791.n428 0.11803
R19069 w_4660_n6791.n736 w_4660_n6791.n735 0.11803
R19070 w_4660_n6791.n737 w_4660_n6791.n736 0.11803
R19071 w_4660_n6791.n738 w_4660_n6791.n737 0.11803
R19072 w_4660_n6791.n739 w_4660_n6791.n738 0.11803
R19073 w_4660_n6791.n740 w_4660_n6791.n739 0.11803
R19074 w_4660_n6791.n741 w_4660_n6791.n740 0.11803
R19075 w_4660_n6791.n742 w_4660_n6791.n741 0.11803
R19076 w_4660_n6791.n743 w_4660_n6791.n742 0.11803
R19077 w_4660_n6791.n744 w_4660_n6791.n743 0.11803
R19078 w_4660_n6791.n745 w_4660_n6791.n744 0.11803
R19079 w_4660_n6791.n746 w_4660_n6791.n745 0.11803
R19080 w_4660_n6791.n747 w_4660_n6791.n746 0.11803
R19081 w_4660_n6791.n748 w_4660_n6791.n747 0.11803
R19082 w_4660_n6791.n749 w_4660_n6791.n748 0.11803
R19083 w_4660_n6791.n750 w_4660_n6791.n749 0.11803
R19084 w_4660_n6791.n751 w_4660_n6791.n750 0.11803
R19085 w_4660_n6791.n752 w_4660_n6791.n751 0.11803
R19086 w_4660_n6791.n753 w_4660_n6791.n752 0.11803
R19087 w_4660_n6791.n754 w_4660_n6791.n753 0.11803
R19088 w_4660_n6791.n755 w_4660_n6791.n754 0.11803
R19089 w_4660_n6791.n756 w_4660_n6791.n755 0.11803
R19090 w_4660_n6791.n757 w_4660_n6791.n756 0.11803
R19091 w_4660_n6791.n758 w_4660_n6791.n757 0.11803
R19092 w_4660_n6791.n759 w_4660_n6791.n758 0.11803
R19093 w_4660_n6791.n1214 w_4660_n6791.n429 0.11803
R19094 w_4660_n6791.n1214 w_4660_n6791.n1213 0.11803
R19095 w_4660_n6791.n1213 w_4660_n6791.n1212 0.11803
R19096 w_4660_n6791.n1212 w_4660_n6791.n1211 0.11803
R19097 w_4660_n6791.n1211 w_4660_n6791.n1210 0.11803
R19098 w_4660_n6791.n1210 w_4660_n6791.n1209 0.11803
R19099 w_4660_n6791.n1209 w_4660_n6791.n1208 0.11803
R19100 w_4660_n6791.n1208 w_4660_n6791.n1207 0.11803
R19101 w_4660_n6791.n1207 w_4660_n6791.n1206 0.11803
R19102 w_4660_n6791.n1206 w_4660_n6791.n1205 0.11803
R19103 w_4660_n6791.n1205 w_4660_n6791.n1204 0.11803
R19104 w_4660_n6791.n1204 w_4660_n6791.n1203 0.11803
R19105 w_4660_n6791.n1203 w_4660_n6791.n1202 0.11803
R19106 w_4660_n6791.n1202 w_4660_n6791.n1201 0.11803
R19107 w_4660_n6791.n1201 w_4660_n6791.n1200 0.11803
R19108 w_4660_n6791.n1200 w_4660_n6791.n1199 0.11803
R19109 w_4660_n6791.n1199 w_4660_n6791.n1198 0.11803
R19110 w_4660_n6791.n1198 w_4660_n6791.n1197 0.11803
R19111 w_4660_n6791.n1197 w_4660_n6791.n1196 0.11803
R19112 w_4660_n6791.n1196 w_4660_n6791.n1195 0.11803
R19113 w_4660_n6791.n1195 w_4660_n6791.n1194 0.11803
R19114 w_4660_n6791.n1194 w_4660_n6791.n1193 0.11803
R19115 w_4660_n6791.n1193 w_4660_n6791.n1192 0.11803
R19116 w_4660_n6791.n1192 w_4660_n6791.n1191 0.11803
R19117 w_4660_n6791.n1191 w_4660_n6791.n1190 0.11803
R19118 w_4660_n6791.n2298 w_4660_n6791.n2277 0.11803
R19119 w_4660_n6791.n2301 w_4660_n6791.n2298 0.11803
R19120 w_4660_n6791.n2301 w_4660_n6791.n2300 0.11803
R19121 w_4660_n6791.n2300 w_4660_n6791.n407 0.11803
R19122 w_4660_n6791.n2325 w_4660_n6791.n407 0.11803
R19123 w_4660_n6791.n2328 w_4660_n6791.n2325 0.11803
R19124 w_4660_n6791.n2328 w_4660_n6791.n2327 0.11803
R19125 w_4660_n6791.n2327 w_4660_n6791.n385 0.11803
R19126 w_4660_n6791.n2352 w_4660_n6791.n385 0.11803
R19127 w_4660_n6791.n2357 w_4660_n6791.n2352 0.11803
R19128 w_4660_n6791.n2357 w_4660_n6791.n2356 0.11803
R19129 w_4660_n6791.n2356 w_4660_n6791.n2355 0.11803
R19130 w_4660_n6791.n2355 w_4660_n6791.n360 0.11803
R19131 w_4660_n6791.n2391 w_4660_n6791.n360 0.11803
R19132 w_4660_n6791.n2396 w_4660_n6791.n2391 0.11803
R19133 w_4660_n6791.n2396 w_4660_n6791.n2395 0.11803
R19134 w_4660_n6791.n2395 w_4660_n6791.n2394 0.11803
R19135 w_4660_n6791.n2394 w_4660_n6791.n334 0.11803
R19136 w_4660_n6791.n2431 w_4660_n6791.n334 0.11803
R19137 w_4660_n6791.n2434 w_4660_n6791.n2431 0.11803
R19138 w_4660_n6791.n2434 w_4660_n6791.n2433 0.11803
R19139 w_4660_n6791.n2433 w_4660_n6791.n313 0.11803
R19140 w_4660_n6791.n2458 w_4660_n6791.n313 0.11803
R19141 w_4660_n6791.n2460 w_4660_n6791.n2458 0.11803
R19142 w_4660_n6791.n2460 w_4660_n6791.n2459 0.11803
R19143 w_4660_n6791.n1471 w_4660_n6791.n458 0.0864598
R19144 w_4660_n6791.n2469 w_4660_n6791.n299 0.081038
R19145 w_4660_n6791.n2276 w_4660_n6791.n427 0.0575
R19146 w_4660_n6791.n2275 w_4660_n6791.n428 0.0572729
R19147 w_4660_n6791.n2274 w_4660_n6791.n429 0.0572729
R19148 w_4660_n6791.n2703 w_4660_n6791.n2702 0.0568974
R19149 w_4660_n6791.n2702 w_4660_n6791.n43 0.0472088
R19150 w_4660_n6791.n2098 w_4660_n6791.n1925 0.0457128
R19151 w_4660_n6791.n988 w_4660_n6791.n939 0.042
R19152 w_4660_n6791.n768 w_4660_n6791.n458 0.042
R19153 w_4660_n6791.n254 w_4660_n6791.n143 0.042
R19154 w_4660_n6791.n2697 w_4660_n6791.n46 0.0412801
R19155 w_4660_n6791.n1411 w_4660_n6791.n988 0.041
R19156 w_4660_n6791.n769 w_4660_n6791.n768 0.041
R19157 w_4660_n6791.n2075 w_4660_n6791.n2074 0.0390638
R19158 w_4660_n6791.n74 w_4660_n6791.n66 0.038
R19159 w_4660_n6791.n1419 w_4660_n6791.n501 0.038
R19160 w_4660_n6791.n1424 w_4660_n6791.n501 0.038
R19161 w_4660_n6791.n1424 w_4660_n6791.n497 0.038
R19162 w_4660_n6791.n1428 w_4660_n6791.n497 0.038
R19163 w_4660_n6791.n1428 w_4660_n6791.n493 0.038
R19164 w_4660_n6791.n1432 w_4660_n6791.n493 0.038
R19165 w_4660_n6791.n1432 w_4660_n6791.n489 0.038
R19166 w_4660_n6791.n1436 w_4660_n6791.n489 0.038
R19167 w_4660_n6791.n1436 w_4660_n6791.n485 0.038
R19168 w_4660_n6791.n1440 w_4660_n6791.n485 0.038
R19169 w_4660_n6791.n1440 w_4660_n6791.n481 0.038
R19170 w_4660_n6791.n1444 w_4660_n6791.n481 0.038
R19171 w_4660_n6791.n1444 w_4660_n6791.n477 0.038
R19172 w_4660_n6791.n1449 w_4660_n6791.n477 0.038
R19173 w_4660_n6791.n1449 w_4660_n6791.n473 0.038
R19174 w_4660_n6791.n1453 w_4660_n6791.n473 0.038
R19175 w_4660_n6791.n1453 w_4660_n6791.n469 0.038
R19176 w_4660_n6791.n1457 w_4660_n6791.n469 0.038
R19177 w_4660_n6791.n1457 w_4660_n6791.n466 0.038
R19178 w_4660_n6791.n1462 w_4660_n6791.n466 0.038
R19179 w_4660_n6791.n1462 w_4660_n6791.n463 0.038
R19180 w_4660_n6791.n1467 w_4660_n6791.n463 0.038
R19181 w_4660_n6791.n1467 w_4660_n6791.n460 0.038
R19182 w_4660_n6791.n1473 w_4660_n6791.n460 0.038
R19183 w_4660_n6791.n1517 w_4660_n6791.n455 0.038
R19184 w_4660_n6791.n1517 w_4660_n6791.n457 0.038
R19185 w_4660_n6791.n1513 w_4660_n6791.n457 0.038
R19186 w_4660_n6791.n1513 w_4660_n6791.n1480 0.038
R19187 w_4660_n6791.n1509 w_4660_n6791.n1480 0.038
R19188 w_4660_n6791.n1509 w_4660_n6791.n1484 0.038
R19189 w_4660_n6791.n1505 w_4660_n6791.n1484 0.038
R19190 w_4660_n6791.n1505 w_4660_n6791.n1488 0.038
R19191 w_4660_n6791.n1501 w_4660_n6791.n1488 0.038
R19192 w_4660_n6791.n1501 w_4660_n6791.n1492 0.038
R19193 w_4660_n6791.n1497 w_4660_n6791.n1492 0.038
R19194 w_4660_n6791.n1497 w_4660_n6791.n118 0.038
R19195 w_4660_n6791.n2645 w_4660_n6791.n118 0.038
R19196 w_4660_n6791.n2645 w_4660_n6791.n120 0.038
R19197 w_4660_n6791.n2641 w_4660_n6791.n120 0.038
R19198 w_4660_n6791.n2641 w_4660_n6791.n125 0.038
R19199 w_4660_n6791.n2637 w_4660_n6791.n125 0.038
R19200 w_4660_n6791.n2637 w_4660_n6791.n129 0.038
R19201 w_4660_n6791.n2633 w_4660_n6791.n129 0.038
R19202 w_4660_n6791.n2633 w_4660_n6791.n133 0.038
R19203 w_4660_n6791.n2629 w_4660_n6791.n133 0.038
R19204 w_4660_n6791.n2629 w_4660_n6791.n137 0.038
R19205 w_4660_n6791.n2625 w_4660_n6791.n137 0.038
R19206 w_4660_n6791.n2625 w_4660_n6791.n141 0.038
R19207 w_4660_n6791.n2674 w_4660_n6791.n2673 0.038
R19208 w_4660_n6791.n2673 w_4660_n6791.n87 0.038
R19209 w_4660_n6791.n2669 w_4660_n6791.n87 0.038
R19210 w_4660_n6791.n2669 w_4660_n6791.n91 0.038
R19211 w_4660_n6791.n2665 w_4660_n6791.n91 0.038
R19212 w_4660_n6791.n2665 w_4660_n6791.n96 0.038
R19213 w_4660_n6791.n2661 w_4660_n6791.n96 0.038
R19214 w_4660_n6791.n2661 w_4660_n6791.n100 0.038
R19215 w_4660_n6791.n2657 w_4660_n6791.n100 0.038
R19216 w_4660_n6791.n2657 w_4660_n6791.n104 0.038
R19217 w_4660_n6791.n2653 w_4660_n6791.n104 0.038
R19218 w_4660_n6791.n2653 w_4660_n6791.n108 0.038
R19219 w_4660_n6791.n965 w_4660_n6791.n108 0.038
R19220 w_4660_n6791.n965 w_4660_n6791.n958 0.038
R19221 w_4660_n6791.n969 w_4660_n6791.n958 0.038
R19222 w_4660_n6791.n969 w_4660_n6791.n954 0.038
R19223 w_4660_n6791.n973 w_4660_n6791.n954 0.038
R19224 w_4660_n6791.n973 w_4660_n6791.n950 0.038
R19225 w_4660_n6791.n977 w_4660_n6791.n950 0.038
R19226 w_4660_n6791.n977 w_4660_n6791.n947 0.038
R19227 w_4660_n6791.n982 w_4660_n6791.n947 0.038
R19228 w_4660_n6791.n982 w_4660_n6791.n943 0.038
R19229 w_4660_n6791.n1415 w_4660_n6791.n943 0.038
R19230 w_4660_n6791.n2517 w_4660_n6791.n249 0.038
R19231 w_4660_n6791.n2517 w_4660_n6791.n251 0.038
R19232 w_4660_n6791.n2513 w_4660_n6791.n251 0.038
R19233 w_4660_n6791.n2513 w_4660_n6791.n261 0.038
R19234 w_4660_n6791.n2509 w_4660_n6791.n261 0.038
R19235 w_4660_n6791.n2509 w_4660_n6791.n265 0.038
R19236 w_4660_n6791.n2505 w_4660_n6791.n265 0.038
R19237 w_4660_n6791.n2505 w_4660_n6791.n269 0.038
R19238 w_4660_n6791.n2501 w_4660_n6791.n269 0.038
R19239 w_4660_n6791.n2501 w_4660_n6791.n273 0.038
R19240 w_4660_n6791.n2497 w_4660_n6791.n273 0.038
R19241 w_4660_n6791.n2497 w_4660_n6791.n277 0.038
R19242 w_4660_n6791.n2493 w_4660_n6791.n277 0.038
R19243 w_4660_n6791.n2493 w_4660_n6791.n281 0.038
R19244 w_4660_n6791.n2489 w_4660_n6791.n281 0.038
R19245 w_4660_n6791.n2489 w_4660_n6791.n285 0.038
R19246 w_4660_n6791.n2485 w_4660_n6791.n285 0.038
R19247 w_4660_n6791.n2485 w_4660_n6791.n290 0.038
R19248 w_4660_n6791.n2481 w_4660_n6791.n290 0.038
R19249 w_4660_n6791.n2481 w_4660_n6791.n294 0.038
R19250 w_4660_n6791.n2477 w_4660_n6791.n294 0.038
R19251 w_4660_n6791.n2477 w_4660_n6791.n298 0.038
R19252 w_4660_n6791.n2473 w_4660_n6791.n298 0.038
R19253 w_4660_n6791.n2616 w_4660_n6791.n143 0.037
R19254 w_4660_n6791.n2264 w_4660_n6791.n449 0.0365
R19255 w_4660_n6791.n2260 w_4660_n6791.n449 0.0365
R19256 w_4660_n6791.n2257 w_4660_n6791.n2256 0.0365
R19257 w_4660_n6791.n2256 w_4660_n6791.n5 0.0365
R19258 w_4660_n6791.n6 w_4660_n6791.n5 0.0365
R19259 w_4660_n6791.n2250 w_4660_n6791.n2249 0.0365
R19260 w_4660_n6791.n2249 w_4660_n6791.n1781 0.0365
R19261 w_4660_n6791.n2245 w_4660_n6791.n1786 0.0365
R19262 w_4660_n6791.n2241 w_4660_n6791.n1786 0.0365
R19263 w_4660_n6791.n2238 w_4660_n6791.n2237 0.0365
R19264 w_4660_n6791.n2237 w_4660_n6791.n1795 0.0365
R19265 w_4660_n6791.n2233 w_4660_n6791.n1800 0.0365
R19266 w_4660_n6791.n2229 w_4660_n6791.n1800 0.0365
R19267 w_4660_n6791.n2229 w_4660_n6791.n1805 0.0365
R19268 w_4660_n6791.n2225 w_4660_n6791.n1810 0.0365
R19269 w_4660_n6791.n2221 w_4660_n6791.n1810 0.0365
R19270 w_4660_n6791.n2218 w_4660_n6791.n2217 0.0365
R19271 w_4660_n6791.n2217 w_4660_n6791.n1818 0.0365
R19272 w_4660_n6791.n2213 w_4660_n6791.n1823 0.0365
R19273 w_4660_n6791.n2209 w_4660_n6791.n1823 0.0365
R19274 w_4660_n6791.n8 w_4660_n6791.n2206 0.0365
R19275 w_4660_n6791.n2206 w_4660_n6791.n1830 0.0365
R19276 w_4660_n6791.n2202 w_4660_n6791.n1830 0.0365
R19277 w_4660_n6791.n2199 w_4660_n6791.n2198 0.0365
R19278 w_4660_n6791.n2198 w_4660_n6791.n1839 0.0365
R19279 w_4660_n6791.n2194 w_4660_n6791.n1844 0.0365
R19280 w_4660_n6791.n2190 w_4660_n6791.n1844 0.0365
R19281 w_4660_n6791.n2187 w_4660_n6791.n2186 0.0365
R19282 w_4660_n6791.n2186 w_4660_n6791.n1853 0.0365
R19283 w_4660_n6791.n2181 w_4660_n6791.n1853 0.0365
R19284 w_4660_n6791.n2178 w_4660_n6791.n2177 0.0365
R19285 w_4660_n6791.n2177 w_4660_n6791.n1862 0.0365
R19286 w_4660_n6791.n2173 w_4660_n6791.n1867 0.0365
R19287 w_4660_n6791.n2169 w_4660_n6791.n1867 0.0365
R19288 w_4660_n6791.n2166 w_4660_n6791.n2165 0.0365
R19289 w_4660_n6791.n2165 w_4660_n6791.n1876 0.0365
R19290 w_4660_n6791.n2161 w_4660_n6791.n1880 0.0365
R19291 w_4660_n6791.n2157 w_4660_n6791.n1880 0.0365
R19292 w_4660_n6791.n2157 w_4660_n6791.n1885 0.0365
R19293 w_4660_n6791.n2153 w_4660_n6791.n1890 0.0365
R19294 w_4660_n6791.n2149 w_4660_n6791.n1890 0.0365
R19295 w_4660_n6791.n2146 w_4660_n6791.n2145 0.0365
R19296 w_4660_n6791.n2145 w_4660_n6791.n1898 0.0365
R19297 w_4660_n6791.n2141 w_4660_n6791.n1903 0.0365
R19298 w_4660_n6791.n2137 w_4660_n6791.n1903 0.0365
R19299 w_4660_n6791.n2137 w_4660_n6791.n10 0.0365
R19300 w_4660_n6791.n2133 w_4660_n6791.n1910 0.0365
R19301 w_4660_n6791.n2129 w_4660_n6791.n1910 0.0365
R19302 w_4660_n6791.n2126 w_4660_n6791.n2125 0.0365
R19303 w_4660_n6791.n2125 w_4660_n6791.n1918 0.0365
R19304 w_4660_n6791.n2121 w_4660_n6791.n2117 0.0365
R19305 w_4660_n6791.n2117 w_4660_n6791.n47 0.0365
R19306 w_4660_n6791.n2695 w_4660_n6791.n49 0.0365
R19307 w_4660_n6791.n2691 w_4660_n6791.n49 0.0365
R19308 w_4660_n6791.n2691 w_4660_n6791.n55 0.0365
R19309 w_4660_n6791.n2687 w_4660_n6791.n60 0.0365
R19310 w_4660_n6791.n2683 w_4660_n6791.n60 0.0365
R19311 w_4660_n6791.n1221 w_4660_n6791.n1140 0.0365
R19312 w_4660_n6791.n1226 w_4660_n6791.n1140 0.0365
R19313 w_4660_n6791.n1230 w_4660_n6791.n1136 0.0365
R19314 w_4660_n6791.n1230 w_4660_n6791.n1134 0.0365
R19315 w_4660_n6791.n1234 w_4660_n6791.n1134 0.0365
R19316 w_4660_n6791.n1237 w_4660_n6791.n1128 0.0365
R19317 w_4660_n6791.n1241 w_4660_n6791.n1128 0.0365
R19318 w_4660_n6791.n1244 w_4660_n6791.n1122 0.0365
R19319 w_4660_n6791.n1248 w_4660_n6791.n1122 0.0365
R19320 w_4660_n6791.n1251 w_4660_n6791.n1114 0.0365
R19321 w_4660_n6791.n1255 w_4660_n6791.n1114 0.0365
R19322 w_4660_n6791.n1259 w_4660_n6791.n12 0.0365
R19323 w_4660_n6791.n1259 w_4660_n6791.n1110 0.0365
R19324 w_4660_n6791.n1263 w_4660_n6791.n1110 0.0365
R19325 w_4660_n6791.n1266 w_4660_n6791.n1104 0.0365
R19326 w_4660_n6791.n1270 w_4660_n6791.n1104 0.0365
R19327 w_4660_n6791.n1273 w_4660_n6791.n1096 0.0365
R19328 w_4660_n6791.n1278 w_4660_n6791.n1096 0.0365
R19329 w_4660_n6791.n1282 w_4660_n6791.n1092 0.0365
R19330 w_4660_n6791.n1282 w_4660_n6791.n1090 0.0365
R19331 w_4660_n6791.n1286 w_4660_n6791.n1090 0.0365
R19332 w_4660_n6791.n1289 w_4660_n6791.n1084 0.0365
R19333 w_4660_n6791.n1293 w_4660_n6791.n1084 0.0365
R19334 w_4660_n6791.n1296 w_4660_n6791.n1078 0.0365
R19335 w_4660_n6791.n1300 w_4660_n6791.n1078 0.0365
R19336 w_4660_n6791.n1303 w_4660_n6791.n1072 0.0365
R19337 w_4660_n6791.n1307 w_4660_n6791.n1072 0.0365
R19338 w_4660_n6791.n1311 w_4660_n6791.n1066 0.0365
R19339 w_4660_n6791.n1316 w_4660_n6791.n1066 0.0365
R19340 w_4660_n6791.n1319 w_4660_n6791.n1316 0.0365
R19341 w_4660_n6791.n1322 w_4660_n6791.n1060 0.0365
R19342 w_4660_n6791.n1326 w_4660_n6791.n1060 0.0365
R19343 w_4660_n6791.n1329 w_4660_n6791.n1052 0.0365
R19344 w_4660_n6791.n1334 w_4660_n6791.n1052 0.0365
R19345 w_4660_n6791.n1338 w_4660_n6791.n1048 0.0365
R19346 w_4660_n6791.n1338 w_4660_n6791.n1046 0.0365
R19347 w_4660_n6791.n14 w_4660_n6791.n1046 0.0365
R19348 w_4660_n6791.n1344 w_4660_n6791.n1042 0.0365
R19349 w_4660_n6791.n1348 w_4660_n6791.n1042 0.0365
R19350 w_4660_n6791.n1351 w_4660_n6791.n1036 0.0365
R19351 w_4660_n6791.n1355 w_4660_n6791.n1036 0.0365
R19352 w_4660_n6791.n1358 w_4660_n6791.n1028 0.0365
R19353 w_4660_n6791.n1363 w_4660_n6791.n1028 0.0365
R19354 w_4660_n6791.n1367 w_4660_n6791.n1024 0.0365
R19355 w_4660_n6791.n1367 w_4660_n6791.n1022 0.0365
R19356 w_4660_n6791.n1371 w_4660_n6791.n1022 0.0365
R19357 w_4660_n6791.n1374 w_4660_n6791.n1016 0.0365
R19358 w_4660_n6791.n1378 w_4660_n6791.n1016 0.0365
R19359 w_4660_n6791.n1381 w_4660_n6791.n1010 0.0365
R19360 w_4660_n6791.n1385 w_4660_n6791.n1010 0.0365
R19361 w_4660_n6791.n1388 w_4660_n6791.n1003 0.0365
R19362 w_4660_n6791.n1393 w_4660_n6791.n1003 0.0365
R19363 w_4660_n6791.n1397 w_4660_n6791.n16 0.0365
R19364 w_4660_n6791.n1397 w_4660_n6791.n999 0.0365
R19365 w_4660_n6791.n1401 w_4660_n6791.n999 0.0365
R19366 w_4660_n6791.n1404 w_4660_n6791.n993 0.0365
R19367 w_4660_n6791.n1408 w_4660_n6791.n993 0.0365
R19368 w_4660_n6791.n932 w_4660_n6791.n931 0.0365
R19369 w_4660_n6791.n931 w_4660_n6791.n509 0.0365
R19370 w_4660_n6791.n927 w_4660_n6791.n514 0.0365
R19371 w_4660_n6791.n923 w_4660_n6791.n514 0.0365
R19372 w_4660_n6791.n923 w_4660_n6791.n519 0.0365
R19373 w_4660_n6791.n919 w_4660_n6791.n524 0.0365
R19374 w_4660_n6791.n915 w_4660_n6791.n524 0.0365
R19375 w_4660_n6791.n912 w_4660_n6791.n911 0.0365
R19376 w_4660_n6791.n911 w_4660_n6791.n532 0.0365
R19377 w_4660_n6791.n907 w_4660_n6791.n537 0.0365
R19378 w_4660_n6791.n903 w_4660_n6791.n537 0.0365
R19379 w_4660_n6791.n18 w_4660_n6791.n900 0.0365
R19380 w_4660_n6791.n900 w_4660_n6791.n544 0.0365
R19381 w_4660_n6791.n896 w_4660_n6791.n544 0.0365
R19382 w_4660_n6791.n893 w_4660_n6791.n892 0.0365
R19383 w_4660_n6791.n892 w_4660_n6791.n553 0.0365
R19384 w_4660_n6791.n888 w_4660_n6791.n558 0.0365
R19385 w_4660_n6791.n884 w_4660_n6791.n558 0.0365
R19386 w_4660_n6791.n881 w_4660_n6791.n880 0.0365
R19387 w_4660_n6791.n880 w_4660_n6791.n567 0.0365
R19388 w_4660_n6791.n876 w_4660_n6791.n567 0.0365
R19389 w_4660_n6791.n873 w_4660_n6791.n872 0.0365
R19390 w_4660_n6791.n872 w_4660_n6791.n576 0.0365
R19391 w_4660_n6791.n868 w_4660_n6791.n581 0.0365
R19392 w_4660_n6791.n864 w_4660_n6791.n581 0.0365
R19393 w_4660_n6791.n861 w_4660_n6791.n860 0.0365
R19394 w_4660_n6791.n860 w_4660_n6791.n590 0.0365
R19395 w_4660_n6791.n856 w_4660_n6791.n852 0.0365
R19396 w_4660_n6791.n852 w_4660_n6791.n851 0.0365
R19397 w_4660_n6791.n851 w_4660_n6791.n598 0.0365
R19398 w_4660_n6791.n847 w_4660_n6791.n604 0.0365
R19399 w_4660_n6791.n843 w_4660_n6791.n604 0.0365
R19400 w_4660_n6791.n840 w_4660_n6791.n839 0.0365
R19401 w_4660_n6791.n839 w_4660_n6791.n613 0.0365
R19402 w_4660_n6791.n835 w_4660_n6791.n618 0.0365
R19403 w_4660_n6791.n831 w_4660_n6791.n618 0.0365
R19404 w_4660_n6791.n831 w_4660_n6791.n20 0.0365
R19405 w_4660_n6791.n827 w_4660_n6791.n625 0.0365
R19406 w_4660_n6791.n823 w_4660_n6791.n625 0.0365
R19407 w_4660_n6791.n820 w_4660_n6791.n819 0.0365
R19408 w_4660_n6791.n819 w_4660_n6791.n633 0.0365
R19409 w_4660_n6791.n815 w_4660_n6791.n638 0.0365
R19410 w_4660_n6791.n811 w_4660_n6791.n638 0.0365
R19411 w_4660_n6791.n808 w_4660_n6791.n807 0.0365
R19412 w_4660_n6791.n807 w_4660_n6791.n647 0.0365
R19413 w_4660_n6791.n803 w_4660_n6791.n647 0.0365
R19414 w_4660_n6791.n800 w_4660_n6791.n799 0.0365
R19415 w_4660_n6791.n799 w_4660_n6791.n656 0.0365
R19416 w_4660_n6791.n795 w_4660_n6791.n661 0.0365
R19417 w_4660_n6791.n791 w_4660_n6791.n661 0.0365
R19418 w_4660_n6791.n788 w_4660_n6791.n787 0.0365
R19419 w_4660_n6791.n787 w_4660_n6791.n21 0.0365
R19420 w_4660_n6791.n22 w_4660_n6791.n673 0.0365
R19421 w_4660_n6791.n780 w_4660_n6791.n673 0.0365
R19422 w_4660_n6791.n780 w_4660_n6791.n678 0.0365
R19423 w_4660_n6791.n776 w_4660_n6791.n683 0.0365
R19424 w_4660_n6791.n772 w_4660_n6791.n683 0.0365
R19425 w_4660_n6791.n1756 w_4660_n6791.n1755 0.0365
R19426 w_4660_n6791.n1755 w_4660_n6791.n1526 0.0365
R19427 w_4660_n6791.n1751 w_4660_n6791.n1531 0.0365
R19428 w_4660_n6791.n1747 w_4660_n6791.n1531 0.0365
R19429 w_4660_n6791.n1747 w_4660_n6791.n24 0.0365
R19430 w_4660_n6791.n1743 w_4660_n6791.n1538 0.0365
R19431 w_4660_n6791.n1739 w_4660_n6791.n1538 0.0365
R19432 w_4660_n6791.n1736 w_4660_n6791.n1735 0.0365
R19433 w_4660_n6791.n1735 w_4660_n6791.n1546 0.0365
R19434 w_4660_n6791.n1731 w_4660_n6791.n1551 0.0365
R19435 w_4660_n6791.n1727 w_4660_n6791.n1551 0.0365
R19436 w_4660_n6791.n1724 w_4660_n6791.n1723 0.0365
R19437 w_4660_n6791.n1723 w_4660_n6791.n1560 0.0365
R19438 w_4660_n6791.n1719 w_4660_n6791.n1560 0.0365
R19439 w_4660_n6791.n1716 w_4660_n6791.n1715 0.0365
R19440 w_4660_n6791.n1715 w_4660_n6791.n1569 0.0365
R19441 w_4660_n6791.n1711 w_4660_n6791.n1574 0.0365
R19442 w_4660_n6791.n1707 w_4660_n6791.n1574 0.0365
R19443 w_4660_n6791.n1704 w_4660_n6791.n1703 0.0365
R19444 w_4660_n6791.n1703 w_4660_n6791.n25 0.0365
R19445 w_4660_n6791.n26 w_4660_n6791.n1586 0.0365
R19446 w_4660_n6791.n1696 w_4660_n6791.n1586 0.0365
R19447 w_4660_n6791.n1696 w_4660_n6791.n1591 0.0365
R19448 w_4660_n6791.n1692 w_4660_n6791.n1596 0.0365
R19449 w_4660_n6791.n1688 w_4660_n6791.n1596 0.0365
R19450 w_4660_n6791.n1685 w_4660_n6791.n1684 0.0365
R19451 w_4660_n6791.n1684 w_4660_n6791.n1604 0.0365
R19452 w_4660_n6791.n1680 w_4660_n6791.n1676 0.0365
R19453 w_4660_n6791.n1676 w_4660_n6791.n233 0.0365
R19454 w_4660_n6791.n2526 w_4660_n6791.n233 0.0365
R19455 w_4660_n6791.n2529 w_4660_n6791.n227 0.0365
R19456 w_4660_n6791.n2533 w_4660_n6791.n227 0.0365
R19457 w_4660_n6791.n2536 w_4660_n6791.n221 0.0365
R19458 w_4660_n6791.n2540 w_4660_n6791.n221 0.0365
R19459 w_4660_n6791.n2543 w_4660_n6791.n212 0.0365
R19460 w_4660_n6791.n2547 w_4660_n6791.n212 0.0365
R19461 w_4660_n6791.n2551 w_4660_n6791.n208 0.0365
R19462 w_4660_n6791.n2551 w_4660_n6791.n206 0.0365
R19463 w_4660_n6791.n2555 w_4660_n6791.n206 0.0365
R19464 w_4660_n6791.n2558 w_4660_n6791.n200 0.0365
R19465 w_4660_n6791.n2562 w_4660_n6791.n200 0.0365
R19466 w_4660_n6791.n2565 w_4660_n6791.n191 0.0365
R19467 w_4660_n6791.n2569 w_4660_n6791.n191 0.0365
R19468 w_4660_n6791.n2573 w_4660_n6791.n187 0.0365
R19469 w_4660_n6791.n2573 w_4660_n6791.n185 0.0365
R19470 w_4660_n6791.n28 w_4660_n6791.n185 0.0365
R19471 w_4660_n6791.n2579 w_4660_n6791.n181 0.0365
R19472 w_4660_n6791.n2583 w_4660_n6791.n181 0.0365
R19473 w_4660_n6791.n2586 w_4660_n6791.n175 0.0365
R19474 w_4660_n6791.n2590 w_4660_n6791.n175 0.0365
R19475 w_4660_n6791.n2593 w_4660_n6791.n169 0.0365
R19476 w_4660_n6791.n2597 w_4660_n6791.n169 0.0365
R19477 w_4660_n6791.n2600 w_4660_n6791.n161 0.0365
R19478 w_4660_n6791.n2605 w_4660_n6791.n161 0.0365
R19479 w_4660_n6791.n2605 w_4660_n6791.n153 0.0365
R19480 w_4660_n6791.n2611 w_4660_n6791.n157 0.0365
R19481 w_4660_n6791.n157 w_4660_n6791.n147 0.0365
R19482 w_4660_n6791.n2291 w_4660_n6791.n2284 0.0365
R19483 w_4660_n6791.n2291 w_4660_n6791.n2278 0.0365
R19484 w_4660_n6791.n2296 w_4660_n6791.n2282 0.0365
R19485 w_4660_n6791.n2282 w_4660_n6791.n422 0.0365
R19486 w_4660_n6791.n30 w_4660_n6791.n422 0.0365
R19487 w_4660_n6791.n2305 w_4660_n6791.n29 0.0365
R19488 w_4660_n6791.n2306 w_4660_n6791.n2305 0.0365
R19489 w_4660_n6791.n2309 w_4660_n6791.n416 0.0365
R19490 w_4660_n6791.n2313 w_4660_n6791.n416 0.0365
R19491 w_4660_n6791.n2318 w_4660_n6791.n414 0.0365
R19492 w_4660_n6791.n2318 w_4660_n6791.n408 0.0365
R19493 w_4660_n6791.n2323 w_4660_n6791.n412 0.0365
R19494 w_4660_n6791.n412 w_4660_n6791.n401 0.0365
R19495 w_4660_n6791.n2330 w_4660_n6791.n401 0.0365
R19496 w_4660_n6791.n2334 w_4660_n6791.n399 0.0365
R19497 w_4660_n6791.n2335 w_4660_n6791.n2334 0.0365
R19498 w_4660_n6791.n2338 w_4660_n6791.n394 0.0365
R19499 w_4660_n6791.n2342 w_4660_n6791.n394 0.0365
R19500 w_4660_n6791.n2347 w_4660_n6791.n392 0.0365
R19501 w_4660_n6791.n2347 w_4660_n6791.n386 0.0365
R19502 w_4660_n6791.n31 w_4660_n6791.n390 0.0365
R19503 w_4660_n6791.n390 w_4660_n6791.n379 0.0365
R19504 w_4660_n6791.n2359 w_4660_n6791.n379 0.0365
R19505 w_4660_n6791.n2363 w_4660_n6791.n377 0.0365
R19506 w_4660_n6791.n2364 w_4660_n6791.n2363 0.0365
R19507 w_4660_n6791.n2367 w_4660_n6791.n372 0.0365
R19508 w_4660_n6791.n2371 w_4660_n6791.n372 0.0365
R19509 w_4660_n6791.n2375 w_4660_n6791.n370 0.0365
R19510 w_4660_n6791.n2375 w_4660_n6791.n367 0.0365
R19511 w_4660_n6791.n2380 w_4660_n6791.n367 0.0365
R19512 w_4660_n6791.n2385 w_4660_n6791.n365 0.0365
R19513 w_4660_n6791.n2385 w_4660_n6791.n361 0.0365
R19514 w_4660_n6791.n2389 w_4660_n6791.n354 0.0365
R19515 w_4660_n6791.n2398 w_4660_n6791.n354 0.0365
R19516 w_4660_n6791.n2402 w_4660_n6791.n352 0.0365
R19517 w_4660_n6791.n2403 w_4660_n6791.n2402 0.0365
R19518 w_4660_n6791.n2407 w_4660_n6791.n348 0.0365
R19519 w_4660_n6791.n2411 w_4660_n6791.n348 0.0365
R19520 w_4660_n6791.n2412 w_4660_n6791.n2411 0.0365
R19521 w_4660_n6791.n2415 w_4660_n6791.n343 0.0365
R19522 w_4660_n6791.n2419 w_4660_n6791.n343 0.0365
R19523 w_4660_n6791.n2424 w_4660_n6791.n341 0.0365
R19524 w_4660_n6791.n2424 w_4660_n6791.n335 0.0365
R19525 w_4660_n6791.n2429 w_4660_n6791.n339 0.0365
R19526 w_4660_n6791.n339 w_4660_n6791.n328 0.0365
R19527 w_4660_n6791.n33 w_4660_n6791.n328 0.0365
R19528 w_4660_n6791.n2438 w_4660_n6791.n32 0.0365
R19529 w_4660_n6791.n2439 w_4660_n6791.n2438 0.0365
R19530 w_4660_n6791.n2442 w_4660_n6791.n322 0.0365
R19531 w_4660_n6791.n2446 w_4660_n6791.n322 0.0365
R19532 w_4660_n6791.n2451 w_4660_n6791.n320 0.0365
R19533 w_4660_n6791.n2451 w_4660_n6791.n314 0.0365
R19534 w_4660_n6791.n2456 w_4660_n6791.n318 0.0365
R19535 w_4660_n6791.n318 w_4660_n6791.n307 0.0365
R19536 w_4660_n6791.n2462 w_4660_n6791.n307 0.0365
R19537 w_4660_n6791.n2466 w_4660_n6791.n305 0.0365
R19538 w_4660_n6791.n2467 w_4660_n6791.n2466 0.0365
R19539 w_4660_n6791.n33 w_4660_n6791.n32 0.0365
R19540 w_4660_n6791.n31 w_4660_n6791.n386 0.0365
R19541 w_4660_n6791.n30 w_4660_n6791.n29 0.0365
R19542 w_4660_n6791.n2579 w_4660_n6791.n28 0.0365
R19543 w_4660_n6791.n26 w_4660_n6791.n25 0.0365
R19544 w_4660_n6791.n1743 w_4660_n6791.n24 0.0365
R19545 w_4660_n6791.n22 w_4660_n6791.n21 0.0365
R19546 w_4660_n6791.n827 w_4660_n6791.n20 0.0365
R19547 w_4660_n6791.n903 w_4660_n6791.n18 0.0365
R19548 w_4660_n6791.n1393 w_4660_n6791.n16 0.0365
R19549 w_4660_n6791.n1344 w_4660_n6791.n14 0.0365
R19550 w_4660_n6791.n1255 w_4660_n6791.n12 0.0365
R19551 w_4660_n6791.n2133 w_4660_n6791.n10 0.0365
R19552 w_4660_n6791.n2209 w_4660_n6791.n8 0.0365
R19553 w_4660_n6791.n2250 w_4660_n6791.n6 0.0365
R19554 w_4660_n6791.n2075 w_4660_n6791.n37 0.0364043
R19555 w_4660_n6791.n2267 w_4660_n6791.n40 0.0364043
R19556 w_4660_n6791.n1983 w_4660_n6791.n446 0.0364043
R19557 w_4660_n6791.n1984 w_4660_n6791.n1983 0.0364043
R19558 w_4660_n6791.n1989 w_4660_n6791.n1988 0.0364043
R19559 w_4660_n6791.n1990 w_4660_n6791.n1989 0.0364043
R19560 w_4660_n6791.n1995 w_4660_n6791.n1994 0.0364043
R19561 w_4660_n6791.n1996 w_4660_n6791.n1995 0.0364043
R19562 w_4660_n6791.n2003 w_4660_n6791.n2002 0.0364043
R19563 w_4660_n6791.n2007 w_4660_n6791.n2006 0.0364043
R19564 w_4660_n6791.n2007 w_4660_n6791.n1971 0.0364043
R19565 w_4660_n6791.n2011 w_4660_n6791.n1971 0.0364043
R19566 w_4660_n6791.n2014 w_4660_n6791.n2011 0.0364043
R19567 w_4660_n6791.n2018 w_4660_n6791.n1967 0.0364043
R19568 w_4660_n6791.n2021 w_4660_n6791.n2018 0.0364043
R19569 w_4660_n6791.n2027 w_4660_n6791.n1964 0.0364043
R19570 w_4660_n6791.n2028 w_4660_n6791.n2027 0.0364043
R19571 w_4660_n6791.n2034 w_4660_n6791.n1961 0.0364043
R19572 w_4660_n6791.n2036 w_4660_n6791.n1958 0.0364043
R19573 w_4660_n6791.n2040 w_4660_n6791.n1958 0.0364043
R19574 w_4660_n6791.n2042 w_4660_n6791.n1954 0.0364043
R19575 w_4660_n6791.n2048 w_4660_n6791.n1950 0.0364043
R19576 w_4660_n6791.n2052 w_4660_n6791.n1950 0.0364043
R19577 w_4660_n6791.n2054 w_4660_n6791.n1946 0.0364043
R19578 w_4660_n6791.n2058 w_4660_n6791.n1946 0.0364043
R19579 w_4660_n6791.n2060 w_4660_n6791.n1942 0.0364043
R19580 w_4660_n6791.n2064 w_4660_n6791.n1942 0.0364043
R19581 w_4660_n6791.n2066 w_4660_n6791.n1938 0.0364043
R19582 w_4660_n6791.n2072 w_4660_n6791.n1938 0.0364043
R19583 w_4660_n6791.n2078 w_4660_n6791.n37 0.0364043
R19584 w_4660_n6791.n2079 w_4660_n6791.n2078 0.0364043
R19585 w_4660_n6791.n2083 w_4660_n6791.n2082 0.0364043
R19586 w_4660_n6791.n2084 w_4660_n6791.n2083 0.0364043
R19587 w_4660_n6791.n2088 w_4660_n6791.n2087 0.0364043
R19588 w_4660_n6791.n2091 w_4660_n6791.n2088 0.0364043
R19589 w_4660_n6791.n2095 w_4660_n6791.n1928 0.0364043
R19590 w_4660_n6791.n2096 w_4660_n6791.n2095 0.0364043
R19591 w_4660_n6791.n2102 w_4660_n6791.n1925 0.0364043
R19592 w_4660_n6791.n2105 w_4660_n6791.n2104 0.0364043
R19593 w_4660_n6791.n2105 w_4660_n6791.n1922 0.0364043
R19594 w_4660_n6791.n2110 w_4660_n6791.n46 0.0364043
R19595 w_4660_n6791.n2699 w_4660_n6791.n2698 0.0364043
R19596 w_4660_n6791.n2699 w_4660_n6791.n41 0.0364043
R19597 w_4660_n6791.n2002 w_4660_n6791.n2001 0.035961
R19598 w_4660_n6791.n2030 w_4660_n6791.n1961 0.035961
R19599 w_4660_n6791.n2046 w_4660_n6791.n1954 0.035961
R19600 w_4660_n6791.n1473 w_4660_n6791.n458 0.034875
R19601 w_4660_n6791.n2178 w_4660_n6791.n1857 0.0335
R19602 w_4660_n6791.n36 w_4660_n6791.n1876 0.0335
R19603 w_4660_n6791.n1289 w_4660_n6791.n1086 0.0335
R19604 w_4660_n6791.n1307 w_4660_n6791.n1068 0.0335
R19605 w_4660_n6791.n873 w_4660_n6791.n571 0.0335
R19606 w_4660_n6791.n592 w_4660_n6791.n590 0.0335
R19607 w_4660_n6791.n2529 w_4660_n6791.n229 0.0335
R19608 w_4660_n6791.n2547 w_4660_n6791.n215 0.0335
R19609 w_4660_n6791.n368 w_4660_n6791.n365 0.0335
R19610 w_4660_n6791.n2403 w_4660_n6791.n350 0.0335
R19611 w_4660_n6791.n1 w_4660_n6791.n68 0.0333947
R19612 w_4660_n6791.n1 w_4660_n6791.n66 0.0333125
R19613 w_4660_n6791.n2006 w_4660_n6791.n1975 0.0333014
R19614 w_4660_n6791.n2014 w_4660_n6791.n2013 0.0333014
R19615 w_4660_n6791.n2079 w_4660_n6791.n1934 0.0328582
R19616 w_4660_n6791.n1797 w_4660_n6791.n1795 0.0315
R19617 w_4660_n6791.n2225 w_4660_n6791.n1807 0.0315
R19618 w_4660_n6791.n2696 w_4660_n6791.n47 0.0315
R19619 w_4660_n6791.n2687 w_4660_n6791.n42 0.0315
R19620 w_4660_n6791.n1226 w_4660_n6791.n1215 0.0315
R19621 w_4660_n6791.n1237 w_4660_n6791.n1130 0.0315
R19622 w_4660_n6791.n1363 w_4660_n6791.n1030 0.0315
R19623 w_4660_n6791.n1374 w_4660_n6791.n1018 0.0315
R19624 w_4660_n6791.n511 w_4660_n6791.n509 0.0315
R19625 w_4660_n6791.n919 w_4660_n6791.n521 0.0315
R19626 w_4660_n6791.n811 w_4660_n6791.n643 0.0315
R19627 w_4660_n6791.n800 w_4660_n6791.n651 0.0315
R19628 w_4660_n6791.n1727 w_4660_n6791.n1556 0.0315
R19629 w_4660_n6791.n1716 w_4660_n6791.n1564 0.0315
R19630 w_4660_n6791.n2597 w_4660_n6791.n165 0.0315
R19631 w_4660_n6791.n2612 w_4660_n6791.n2611 0.0315
R19632 w_4660_n6791.n2324 w_4660_n6791.n408 0.0315
R19633 w_4660_n6791.n2329 w_4660_n6791.n399 0.0315
R19634 w_4660_n6791.n2457 w_4660_n6791.n314 0.0315
R19635 w_4660_n6791.n2461 w_4660_n6791.n305 0.0315
R19636 w_4660_n6791.n2074 w_4660_n6791.n2073 0.0310851
R19637 w_4660_n6791.n73 w_4660_n6791.n69 0.0308452
R19638 w_4660_n6791.n2474 w_4660_n6791.n299 0.0308452
R19639 w_4660_n6791.n2001 w_4660_n6791.n1978 0.0306418
R19640 w_4660_n6791.n2084 w_4660_n6791.n1931 0.0297553
R19641 w_4660_n6791.n2190 w_4660_n6791.n1849 0.0295
R19642 w_4660_n6791.n2153 w_4660_n6791.n1887 0.0295
R19643 w_4660_n6791.n1278 w_4660_n6791.n1098 0.0295
R19644 w_4660_n6791.n1322 w_4660_n6791.n1062 0.0295
R19645 w_4660_n6791.n884 w_4660_n6791.n563 0.0295
R19646 w_4660_n6791.n847 w_4660_n6791.n601 0.0295
R19647 w_4660_n6791.n1673 w_4660_n6791.n1604 0.0295
R19648 w_4660_n6791.n2558 w_4660_n6791.n202 0.0295
R19649 w_4660_n6791.n2371 w_4660_n6791.n373 0.0295
R19650 w_4660_n6791.n2415 w_4660_n6791.n346 0.0295
R19651 w_4660_n6791.n2021 w_4660_n6791.n2020 0.0293121
R19652 w_4660_n6791.n2703 w_4660_n6791.n41 0.0288688
R19653 w_4660_n6791.n2111 w_4660_n6791.n2110 0.0284255
R19654 w_4660_n6791.n2066 w_4660_n6791.n2065 0.0279823
R19655 w_4660_n6791.n1994 w_4660_n6791.n1980 0.027539
R19656 w_4660_n6791.n2260 w_4660_n6791.n1769 0.0275
R19657 w_4660_n6791.n2199 w_4660_n6791.n1834 0.0275
R19658 w_4660_n6791.n1900 w_4660_n6791.n1898 0.0275
R19659 w_4660_n6791.n1266 w_4660_n6791.n1106 0.0275
R19660 w_4660_n6791.n1334 w_4660_n6791.n1054 0.0275
R19661 w_4660_n6791.n1404 w_4660_n6791.n995 0.0275
R19662 w_4660_n6791.n893 w_4660_n6791.n548 0.0275
R19663 w_4660_n6791.n615 w_4660_n6791.n613 0.0275
R19664 w_4660_n6791.n776 w_4660_n6791.n680 0.0275
R19665 w_4660_n6791.n1528 w_4660_n6791.n1526 0.0275
R19666 w_4660_n6791.n1692 w_4660_n6791.n1593 0.0275
R19667 w_4660_n6791.n2569 w_4660_n6791.n194 0.0275
R19668 w_4660_n6791.n2297 w_4660_n6791.n2278 0.0275
R19669 w_4660_n6791.n2358 w_4660_n6791.n377 0.0275
R19670 w_4660_n6791.n2430 w_4660_n6791.n335 0.0275
R19671 w_4660_n6791.n2091 w_4660_n6791.n2090 0.0270957
R19672 w_4660_n6791.n2678 w_4660_n6791.n78 0.0263772
R19673 w_4660_n6791.n2029 w_4660_n6791.n2028 0.0262092
R19674 w_4660_n6791.n2245 w_4660_n6791.n1783 0.0255
R19675 w_4660_n6791.n1820 w_4660_n6791.n1818 0.0255
R19676 w_4660_n6791.n2126 w_4660_n6791.n1914 0.0255
R19677 w_4660_n6791.n1248 w_4660_n6791.n1118 0.0255
R19678 w_4660_n6791.n1351 w_4660_n6791.n1038 0.0255
R19679 w_4660_n6791.n1385 w_4660_n6791.n1006 0.0255
R19680 w_4660_n6791.n534 w_4660_n6791.n532 0.0255
R19681 w_4660_n6791.n820 w_4660_n6791.n629 0.0255
R19682 w_4660_n6791.n791 w_4660_n6791.n666 0.0255
R19683 w_4660_n6791.n1736 w_4660_n6791.n1542 0.0255
R19684 w_4660_n6791.n1707 w_4660_n6791.n1579 0.0255
R19685 w_4660_n6791.n2586 w_4660_n6791.n177 0.0255
R19686 w_4660_n6791.n2309 w_4660_n6791.n419 0.0255
R19687 w_4660_n6791.n2342 w_4660_n6791.n395 0.0255
R19688 w_4660_n6791.n2442 w_4660_n6791.n325 0.0255
R19689 w_4660_n6791.n2104 w_4660_n6791.n2103 0.0253227
R19690 w_4660_n6791.n2060 w_4660_n6791.n2059 0.0248794
R19691 w_4660_n6791.n1988 w_4660_n6791.n1982 0.0244362
R19692 w_4660_n6791.n2097 w_4660_n6791.n2096 0.0239929
R19693 w_4660_n6791.n2035 w_4660_n6791.n2034 0.0235496
R19694 w_4660_n6791.n2173 w_4660_n6791.n1864 0.0235
R19695 w_4660_n6791.n2169 w_4660_n6791.n1872 0.0235
R19696 w_4660_n6791.n1296 w_4660_n6791.n1080 0.0235
R19697 w_4660_n6791.n1300 w_4660_n6791.n1074 0.0235
R19698 w_4660_n6791.n868 w_4660_n6791.n578 0.0235
R19699 w_4660_n6791.n864 w_4660_n6791.n586 0.0235
R19700 w_4660_n6791.n2536 w_4660_n6791.n223 0.0235
R19701 w_4660_n6791.n2540 w_4660_n6791.n217 0.0235
R19702 w_4660_n6791.n2390 w_4660_n6791.n2389 0.0235
R19703 w_4660_n6791.n2398 w_4660_n6791.n2397 0.0235
R19704 w_4660_n6791.n458 w_4660_n6791.n455 0.0234167
R19705 w_4660_n6791.n2054 w_4660_n6791.n2053 0.0222199
R19706 w_4660_n6791.n2266 w_4660_n6791.n446 0.0217766
R19707 w_4660_n6791.n2241 w_4660_n6791.n1791 0.0215
R19708 w_4660_n6791.n2218 w_4660_n6791.n1814 0.0215
R19709 w_4660_n6791.n2112 w_4660_n6791.n1918 0.0215
R19710 w_4660_n6791.n1217 w_4660_n6791.n1216 0.0215
R19711 w_4660_n6791.n1244 w_4660_n6791.n1124 0.0215
R19712 w_4660_n6791.n1355 w_4660_n6791.n1032 0.0215
R19713 w_4660_n6791.n1381 w_4660_n6791.n1012 0.0215
R19714 w_4660_n6791.n934 w_4660_n6791.n505 0.0215
R19715 w_4660_n6791.n912 w_4660_n6791.n528 0.0215
R19716 w_4660_n6791.n635 w_4660_n6791.n633 0.0215
R19717 w_4660_n6791.n795 w_4660_n6791.n658 0.0215
R19718 w_4660_n6791.n1548 w_4660_n6791.n1546 0.0215
R19719 w_4660_n6791.n1711 w_4660_n6791.n1571 0.0215
R19720 w_4660_n6791.n2590 w_4660_n6791.n171 0.0215
R19721 w_4660_n6791.n2616 w_4660_n6791.n2615 0.0215
R19722 w_4660_n6791.n2313 w_4660_n6791.n417 0.0215
R19723 w_4660_n6791.n2338 w_4660_n6791.n397 0.0215
R19724 w_4660_n6791.n2446 w_4660_n6791.n323 0.0215
R19725 w_4660_n6791.n2469 w_4660_n6791.n303 0.0215
R19726 w_4660_n6791.n2041 w_4660_n6791.n2040 0.0204468
R19727 w_4660_n6791.n2674 w_4660_n6791.n81 0.0198531
R19728 w_4660_n6791.n2265 w_4660_n6791.n2264 0.0195
R19729 w_4660_n6791.n1841 w_4660_n6791.n1839 0.0195
R19730 w_4660_n6791.n2146 w_4660_n6791.n1894 0.0195
R19731 w_4660_n6791.n1270 w_4660_n6791.n1100 0.0195
R19732 w_4660_n6791.n1329 w_4660_n6791.n1056 0.0195
R19733 w_4660_n6791.n1408 w_4660_n6791.n987 0.0195
R19734 w_4660_n6791.n555 w_4660_n6791.n553 0.0195
R19735 w_4660_n6791.n840 w_4660_n6791.n609 0.0195
R19736 w_4660_n6791.n772 w_4660_n6791.n760 0.0195
R19737 w_4660_n6791.n1756 w_4660_n6791.n1523 0.0195
R19738 w_4660_n6791.n1688 w_4660_n6791.n1600 0.0195
R19739 w_4660_n6791.n2565 w_4660_n6791.n196 0.0195
R19740 w_4660_n6791.n2285 w_4660_n6791.n2284 0.0195
R19741 w_4660_n6791.n2364 w_4660_n6791.n375 0.0195
R19742 w_4660_n6791.n344 w_4660_n6791.n341 0.0195
R19743 w_4660_n6791.n2048 w_4660_n6791.n2047 0.019117
R19744 w_4660_n6791.n2047 w_4660_n6791.n2046 0.0177872
R19745 w_4660_n6791.n2100 w_4660_n6791.n2099 0.0175
R19746 w_4660_n6791.n2108 w_4660_n6791.n44 0.0175
R19747 w_4660_n6791.n2265 w_4660_n6791.n447 0.0175
R19748 w_4660_n6791.n2194 w_4660_n6791.n1841 0.0175
R19749 w_4660_n6791.n2149 w_4660_n6791.n1894 0.0175
R19750 w_4660_n6791.n1273 w_4660_n6791.n1100 0.0175
R19751 w_4660_n6791.n1326 w_4660_n6791.n1056 0.0175
R19752 w_4660_n6791.n1411 w_4660_n6791.n987 0.0175
R19753 w_4660_n6791.n888 w_4660_n6791.n555 0.0175
R19754 w_4660_n6791.n843 w_4660_n6791.n609 0.0175
R19755 w_4660_n6791.n769 w_4660_n6791.n760 0.0175
R19756 w_4660_n6791.n1758 w_4660_n6791.n1523 0.0175
R19757 w_4660_n6791.n1685 w_4660_n6791.n1600 0.0175
R19758 w_4660_n6791.n2562 w_4660_n6791.n196 0.0175
R19759 w_4660_n6791.n2287 w_4660_n6791.n2285 0.0175
R19760 w_4660_n6791.n2367 w_4660_n6791.n375 0.0175
R19761 w_4660_n6791.n2419 w_4660_n6791.n344 0.0175
R19762 w_4660_n6791.n2273 w_4660_n6791.n40 0.0171991
R19763 w_4660_n6791.n1415 w_4660_n6791.n939 0.0171667
R19764 w_4660_n6791.n78 w_4660_n6791.n64 0.017
R19765 w_4660_n6791.n2042 w_4660_n6791.n2041 0.0164574
R19766 w_4660_n6791.n2238 w_4660_n6791.n1791 0.0155
R19767 w_4660_n6791.n2221 w_4660_n6791.n1814 0.0155
R19768 w_4660_n6791.n2121 w_4660_n6791.n2112 0.0155
R19769 w_4660_n6791.n2683 w_4660_n6791.n64 0.0155
R19770 w_4660_n6791.n1221 w_4660_n6791.n1217 0.0155
R19771 w_4660_n6791.n1241 w_4660_n6791.n1124 0.0155
R19772 w_4660_n6791.n1358 w_4660_n6791.n1032 0.0155
R19773 w_4660_n6791.n1378 w_4660_n6791.n1012 0.0155
R19774 w_4660_n6791.n932 w_4660_n6791.n505 0.0155
R19775 w_4660_n6791.n915 w_4660_n6791.n528 0.0155
R19776 w_4660_n6791.n815 w_4660_n6791.n635 0.0155
R19777 w_4660_n6791.n658 w_4660_n6791.n656 0.0155
R19778 w_4660_n6791.n1731 w_4660_n6791.n1548 0.0155
R19779 w_4660_n6791.n1571 w_4660_n6791.n1569 0.0155
R19780 w_4660_n6791.n2593 w_4660_n6791.n171 0.0155
R19781 w_4660_n6791.n2615 w_4660_n6791.n147 0.0155
R19782 w_4660_n6791.n417 w_4660_n6791.n414 0.0155
R19783 w_4660_n6791.n2335 w_4660_n6791.n397 0.0155
R19784 w_4660_n6791.n323 w_4660_n6791.n320 0.0155
R19785 w_4660_n6791.n2467 w_4660_n6791.n303 0.0155
R19786 w_4660_n6791.n2267 w_4660_n6791.n2266 0.0151277
R19787 w_4660_n6791.n254 w_4660_n6791.n141 0.0150833
R19788 w_4660_n6791.n2076 w_4660_n6791.n1936 0.015
R19789 w_4660_n6791.n2053 w_4660_n6791.n2052 0.0146844
R19790 w_4660_n6791.n2016 w_4660_n6791.n2015 0.0143333
R19791 w_4660_n6791.n2269 w_4660_n6791.n2268 0.014
R19792 w_4660_n6791.n2268 w_4660_n6791.n34 0.014
R19793 w_4660_n6791.n35 w_4660_n6791.n34 0.014
R19794 w_4660_n6791.n1991 w_4660_n6791.n38 0.014
R19795 w_4660_n6791.n1993 w_4660_n6791.n1991 0.014
R19796 w_4660_n6791.n1997 w_4660_n6791.n0 0.014
R19797 w_4660_n6791.n2000 w_4660_n6791.n1997 0.014
R19798 w_4660_n6791.n2004 w_4660_n6791.n1976 0.014
R19799 w_4660_n6791.n2005 w_4660_n6791.n2004 0.014
R19800 w_4660_n6791.n2009 w_4660_n6791.n2008 0.014
R19801 w_4660_n6791.n2010 w_4660_n6791.n2009 0.014
R19802 w_4660_n6791.n2017 w_4660_n6791.n2016 0.014
R19803 w_4660_n6791.n2023 w_4660_n6791.n2022 0.014
R19804 w_4660_n6791.n2026 w_4660_n6791.n2023 0.014
R19805 w_4660_n6791.n2031 w_4660_n6791.n1962 0.014
R19806 w_4660_n6791.n2033 w_4660_n6791.n2032 0.014
R19807 w_4660_n6791.n2038 w_4660_n6791.n2037 0.014
R19808 w_4660_n6791.n2039 w_4660_n6791.n2038 0.014
R19809 w_4660_n6791.n2044 w_4660_n6791.n2043 0.014
R19810 w_4660_n6791.n2050 w_4660_n6791.n2049 0.014
R19811 w_4660_n6791.n2051 w_4660_n6791.n2050 0.014
R19812 w_4660_n6791.n2056 w_4660_n6791.n2055 0.014
R19813 w_4660_n6791.n2057 w_4660_n6791.n2056 0.014
R19814 w_4660_n6791.n2062 w_4660_n6791.n2061 0.014
R19815 w_4660_n6791.n2063 w_4660_n6791.n2062 0.014
R19816 w_4660_n6791.n2068 w_4660_n6791.n2067 0.014
R19817 w_4660_n6791.n2071 w_4660_n6791.n2068 0.014
R19818 w_4660_n6791.n4 w_4660_n6791.n2076 0.014
R19819 w_4660_n6791.n2080 w_4660_n6791.n3 0.014
R19820 w_4660_n6791.n2081 w_4660_n6791.n2080 0.014
R19821 w_4660_n6791.n2081 w_4660_n6791.n1932 0.014
R19822 w_4660_n6791.n2085 w_4660_n6791.n1932 0.014
R19823 w_4660_n6791.n2086 w_4660_n6791.n1929 0.014
R19824 w_4660_n6791.n2092 w_4660_n6791.n1929 0.014
R19825 w_4660_n6791.n2093 w_4660_n6791.n2092 0.014
R19826 w_4660_n6791.n2094 w_4660_n6791.n2093 0.014
R19827 w_4660_n6791.n2094 w_4660_n6791.n1926 0.014
R19828 w_4660_n6791.n2099 w_4660_n6791.n1926 0.014
R19829 w_4660_n6791.n2101 w_4660_n6791.n2100 0.014
R19830 w_4660_n6791.n2101 w_4660_n6791.n1923 0.014
R19831 w_4660_n6791.n2106 w_4660_n6791.n1923 0.014
R19832 w_4660_n6791.n2107 w_4660_n6791.n2106 0.014
R19833 w_4660_n6791.n2109 w_4660_n6791.n2107 0.014
R19834 w_4660_n6791.n2109 w_4660_n6791.n2108 0.014
R19835 w_4660_n6791.n2700 w_4660_n6791.n44 0.014
R19836 w_4660_n6791.n2701 w_4660_n6791.n2700 0.014
R19837 w_4660_n6791.n1987 w_4660_n6791.n38 0.014
R19838 w_4660_n6791.n1985 w_4660_n6791.n35 0.014
R19839 w_4660_n6791.n4 w_4660_n6791.n3 0.014
R19840 w_4660_n6791.n1993 w_4660_n6791.n0 0.014
R19841 w_4660_n6791.n1987 w_4660_n6791.n1985 0.0138333
R19842 w_4660_n6791.n2032 w_4660_n6791.n2031 0.0138333
R19843 w_4660_n6791.n2045 w_4660_n6791.n2044 0.0138333
R19844 w_4660_n6791.n2086 w_4660_n6791.n2085 0.0138333
R19845 w_4660_n6791.n1864 w_4660_n6791.n1862 0.0135
R19846 w_4660_n6791.n2166 w_4660_n6791.n1872 0.0135
R19847 w_4660_n6791.n1293 w_4660_n6791.n1080 0.0135
R19848 w_4660_n6791.n1303 w_4660_n6791.n1074 0.0135
R19849 w_4660_n6791.n578 w_4660_n6791.n576 0.0135
R19850 w_4660_n6791.n861 w_4660_n6791.n586 0.0135
R19851 w_4660_n6791.n2533 w_4660_n6791.n223 0.0135
R19852 w_4660_n6791.n2543 w_4660_n6791.n217 0.0135
R19853 w_4660_n6791.n2390 w_4660_n6791.n361 0.0135
R19854 w_4660_n6791.n2397 w_4660_n6791.n352 0.0135
R19855 w_4660_n6791.n2036 w_4660_n6791.n2035 0.0133546
R19856 w_4660_n6791.n2678 w_4660_n6791.n81 0.0132193
R19857 w_4660_n6791.n2098 w_4660_n6791.n2097 0.0129113
R19858 w_4660_n6791.n1984 w_4660_n6791.n1982 0.0120248
R19859 w_4660_n6791.n2059 w_4660_n6791.n2058 0.0115816
R19860 w_4660_n6791.n2103 w_4660_n6791.n2102 0.0115816
R19861 w_4660_n6791.n2000 w_4660_n6791.n1999 0.0115
R19862 w_4660_n6791.n1783 w_4660_n6791.n1781 0.0115
R19863 w_4660_n6791.n2213 w_4660_n6791.n1820 0.0115
R19864 w_4660_n6791.n2129 w_4660_n6791.n1914 0.0115
R19865 w_4660_n6791.n1251 w_4660_n6791.n1118 0.0115
R19866 w_4660_n6791.n1348 w_4660_n6791.n1038 0.0115
R19867 w_4660_n6791.n1388 w_4660_n6791.n1006 0.0115
R19868 w_4660_n6791.n907 w_4660_n6791.n534 0.0115
R19869 w_4660_n6791.n823 w_4660_n6791.n629 0.0115
R19870 w_4660_n6791.n788 w_4660_n6791.n666 0.0115
R19871 w_4660_n6791.n1739 w_4660_n6791.n1542 0.0115
R19872 w_4660_n6791.n1704 w_4660_n6791.n1579 0.0115
R19873 w_4660_n6791.n2583 w_4660_n6791.n177 0.0115
R19874 w_4660_n6791.n2306 w_4660_n6791.n419 0.0115
R19875 w_4660_n6791.n395 w_4660_n6791.n392 0.0115
R19876 w_4660_n6791.n2439 w_4660_n6791.n325 0.0115
R19877 w_4660_n6791.n2030 w_4660_n6791.n2029 0.010695
R19878 w_4660_n6791.n2070 w_4660_n6791.n1936 0.0106667
R19879 w_4660_n6791.n2005 w_4660_n6791.n1973 0.0105
R19880 w_4660_n6791.n2033 w_4660_n6791.n1959 0.0105
R19881 w_4660_n6791.n2090 w_4660_n6791.n1928 0.00980851
R19882 w_4660_n6791.n2270 w_4660_n6791.n40 0.00957195
R19883 w_4660_n6791.n2067 w_4660_n6791.n1940 0.0095
R19884 w_4660_n6791.n2257 w_4660_n6791.n1769 0.0095
R19885 w_4660_n6791.n2202 w_4660_n6791.n1834 0.0095
R19886 w_4660_n6791.n2141 w_4660_n6791.n1900 0.0095
R19887 w_4660_n6791.n1263 w_4660_n6791.n1106 0.0095
R19888 w_4660_n6791.n1054 w_4660_n6791.n1048 0.0095
R19889 w_4660_n6791.n1401 w_4660_n6791.n995 0.0095
R19890 w_4660_n6791.n896 w_4660_n6791.n548 0.0095
R19891 w_4660_n6791.n835 w_4660_n6791.n615 0.0095
R19892 w_4660_n6791.n680 w_4660_n6791.n678 0.0095
R19893 w_4660_n6791.n1751 w_4660_n6791.n1528 0.0095
R19894 w_4660_n6791.n1593 w_4660_n6791.n1591 0.0095
R19895 w_4660_n6791.n194 w_4660_n6791.n187 0.0095
R19896 w_4660_n6791.n2297 w_4660_n6791.n2296 0.0095
R19897 w_4660_n6791.n2359 w_4660_n6791.n2358 0.0095
R19898 w_4660_n6791.n2430 w_4660_n6791.n2429 0.0095
R19899 w_4660_n6791.n2271 w_4660_n6791.n2270 0.00940982
R19900 w_4660_n6791.n1990 w_4660_n6791.n1980 0.00936525
R19901 w_4660_n6791.n2010 w_4660_n6791.n1969 0.00933333
R19902 w_4660_n6791.n2039 w_4660_n6791.n1956 0.00933333
R19903 w_4660_n6791.n2065 w_4660_n6791.n2064 0.00892199
R19904 w_4660_n6791.n74 w_4660_n6791.n73 0.00862405
R19905 w_4660_n6791.n2474 w_4660_n6791.n2473 0.00862405
R19906 w_4660_n6791.n2111 w_4660_n6791.n1922 0.00847872
R19907 w_4660_n6791.n2045 w_4660_n6791.n1952 0.00833333
R19908 w_4660_n6791.n2061 w_4660_n6791.n1944 0.00833333
R19909 w_4660_n6791.n2017 w_4660_n6791.n1966 0.00783333
R19910 w_4660_n6791.n2025 w_4660_n6791.n1962 0.00783333
R19911 w_4660_n6791.n39 w_4660_n6791.n430 0.00773667
R19912 w_4660_n6791.n438 w_4660_n6791.n430 0.00773667
R19913 w_4660_n6791.n442 w_4660_n6791.n431 0.00773667
R19914 w_4660_n6791.n439 w_4660_n6791.n431 0.00773667
R19915 w_4660_n6791.n443 w_4660_n6791.n432 0.00773667
R19916 w_4660_n6791.n440 w_4660_n6791.n432 0.00773667
R19917 w_4660_n6791.n441 w_4660_n6791.n433 0.00773667
R19918 w_4660_n6791.n2269 w_4660_n6791.n434 0.00773667
R19919 w_4660_n6791.n445 w_4660_n6791.n441 0.00773667
R19920 w_4660_n6791.n440 w_4660_n6791.n435 0.00773667
R19921 w_4660_n6791.n439 w_4660_n6791.n436 0.00773667
R19922 w_4660_n6791.n438 w_4660_n6791.n437 0.00773667
R19923 w_4660_n6791.n443 w_4660_n6791.n436 0.00773667
R19924 w_4660_n6791.n442 w_4660_n6791.n437 0.00773667
R19925 w_4660_n6791.n2272 w_4660_n6791.n39 0.00773667
R19926 w_4660_n6791.n445 w_4660_n6791.n434 0.00773667
R19927 w_4660_n6791.n444 w_4660_n6791.n433 0.00765366
R19928 w_4660_n6791.n444 w_4660_n6791.n435 0.00765366
R19929 w_4660_n6791.n2020 w_4660_n6791.n1964 0.0075922
R19930 w_4660_n6791.n2187 w_4660_n6791.n1849 0.0075
R19931 w_4660_n6791.n1887 w_4660_n6791.n1885 0.0075
R19932 w_4660_n6791.n1098 w_4660_n6791.n1092 0.0075
R19933 w_4660_n6791.n1319 w_4660_n6791.n1062 0.0075
R19934 w_4660_n6791.n881 w_4660_n6791.n563 0.0075
R19935 w_4660_n6791.n601 w_4660_n6791.n598 0.0075
R19936 w_4660_n6791.n1680 w_4660_n6791.n1673 0.0075
R19937 w_4660_n6791.n2555 w_4660_n6791.n202 0.0075
R19938 w_4660_n6791.n373 w_4660_n6791.n370 0.0075
R19939 w_4660_n6791.n2412 w_4660_n6791.n346 0.0075
R19940 w_4660_n6791.n2055 w_4660_n6791.n1948 0.00733333
R19941 w_4660_n6791.n2051 w_4660_n6791.n1948 0.00716667
R19942 w_4660_n6791.n2087 w_4660_n6791.n1931 0.00670567
R19943 w_4660_n6791.n2022 w_4660_n6791.n1966 0.00666667
R19944 w_4660_n6791.n2026 w_4660_n6791.n2025 0.00666667
R19945 w_4660_n6791.n1996 w_4660_n6791.n1978 0.00626241
R19946 w_4660_n6791.n78 w_4660_n6791.n68 0.00620175
R19947 w_4660_n6791.n2049 w_4660_n6791.n1952 0.00616667
R19948 w_4660_n6791.n2057 w_4660_n6791.n1944 0.006
R19949 w_4660_n6791.n2073 w_4660_n6791.n2072 0.00581915
R19950 w_4660_n6791.n254 w_4660_n6791.n249 0.00570833
R19951 w_4660_n6791.n2233 w_4660_n6791.n1797 0.0055
R19952 w_4660_n6791.n1807 w_4660_n6791.n1805 0.0055
R19953 w_4660_n6791.n2696 w_4660_n6791.n2695 0.0055
R19954 w_4660_n6791.n55 w_4660_n6791.n42 0.0055
R19955 w_4660_n6791.n1215 w_4660_n6791.n1136 0.0055
R19956 w_4660_n6791.n1234 w_4660_n6791.n1130 0.0055
R19957 w_4660_n6791.n1030 w_4660_n6791.n1024 0.0055
R19958 w_4660_n6791.n1371 w_4660_n6791.n1018 0.0055
R19959 w_4660_n6791.n927 w_4660_n6791.n511 0.0055
R19960 w_4660_n6791.n521 w_4660_n6791.n519 0.0055
R19961 w_4660_n6791.n808 w_4660_n6791.n643 0.0055
R19962 w_4660_n6791.n803 w_4660_n6791.n651 0.0055
R19963 w_4660_n6791.n1724 w_4660_n6791.n1556 0.0055
R19964 w_4660_n6791.n1719 w_4660_n6791.n1564 0.0055
R19965 w_4660_n6791.n2600 w_4660_n6791.n165 0.0055
R19966 w_4660_n6791.n2612 w_4660_n6791.n153 0.0055
R19967 w_4660_n6791.n2324 w_4660_n6791.n2323 0.0055
R19968 w_4660_n6791.n2330 w_4660_n6791.n2329 0.0055
R19969 w_4660_n6791.n2457 w_4660_n6791.n2456 0.0055
R19970 w_4660_n6791.n2462 w_4660_n6791.n2461 0.0055
R19971 w_4660_n6791.n2015 w_4660_n6791.n1969 0.00516667
R19972 w_4660_n6791.n2043 w_4660_n6791.n1956 0.00516667
R19973 w_4660_n6791.n2063 w_4660_n6791.n1940 0.005
R19974 w_4660_n6791.n2698 w_4660_n6791.n2697 0.00493262
R19975 w_4660_n6791.n2013 w_4660_n6791.n1967 0.00448936
R19976 w_4660_n6791.n2082 w_4660_n6791.n1934 0.0040461
R19977 w_4660_n6791.n2008 w_4660_n6791.n1973 0.004
R19978 w_4660_n6791.n2037 w_4660_n6791.n1959 0.004
R19979 w_4660_n6791.n2071 w_4660_n6791.n2070 0.00383333
R19980 w_4660_n6791.n1419 w_4660_n6791.n939 0.003625
R19981 w_4660_n6791.n2003 w_4660_n6791.n1975 0.00360284
R19982 w_4660_n6791.n2181 w_4660_n6791.n1857 0.0035
R19983 w_4660_n6791.n2161 w_4660_n6791.n36 0.0035
R19984 w_4660_n6791.n1286 w_4660_n6791.n1086 0.0035
R19985 w_4660_n6791.n1311 w_4660_n6791.n1068 0.0035
R19986 w_4660_n6791.n876 w_4660_n6791.n571 0.0035
R19987 w_4660_n6791.n856 w_4660_n6791.n592 0.0035
R19988 w_4660_n6791.n2526 w_4660_n6791.n229 0.0035
R19989 w_4660_n6791.n215 w_4660_n6791.n208 0.0035
R19990 w_4660_n6791.n2380 w_4660_n6791.n368 0.0035
R19991 w_4660_n6791.n2407 w_4660_n6791.n350 0.0035
R19992 w_4660_n6791.n1999 w_4660_n6791.n1976 0.00283333
R19993 vin_p.n196 vin_p.t36 321.697
R19994 vin_p.n196 vin_p.t34 321.697
R19995 vin_p.n194 vin_p.t38 321.697
R19996 vin_p.n194 vin_p.t37 321.697
R19997 vin_p.n192 vin_p.t22 321.697
R19998 vin_p.n192 vin_p.t20 321.697
R19999 vin_p.n190 vin_p.t96 321.697
R20000 vin_p.n190 vin_p.t95 321.697
R20001 vin_p.n188 vin_p.t148 321.697
R20002 vin_p.n188 vin_p.t147 321.697
R20003 vin_p.n186 vin_p.t150 321.697
R20004 vin_p.n186 vin_p.t149 321.697
R20005 vin_p.n184 vin_p.t156 321.697
R20006 vin_p.n184 vin_p.t153 321.697
R20007 vin_p.n182 vin_p.t160 321.697
R20008 vin_p.n182 vin_p.t157 321.697
R20009 vin_p.n180 vin_p.t31 321.697
R20010 vin_p.n180 vin_p.t29 321.697
R20011 vin_p.n178 vin_p.t92 321.697
R20012 vin_p.n178 vin_p.t90 321.697
R20013 vin_p.n176 vin_p.t76 321.697
R20014 vin_p.n176 vin_p.t72 321.697
R20015 vin_p.n174 vin_p.t80 321.697
R20016 vin_p.n174 vin_p.t77 321.697
R20017 vin_p.n172 vin_p.t84 321.697
R20018 vin_p.n172 vin_p.t81 321.697
R20019 vin_p.n170 vin_p.t88 321.697
R20020 vin_p.n170 vin_p.t85 321.697
R20021 vin_p.n168 vin_p.t6 321.697
R20022 vin_p.n168 vin_p.t5 321.697
R20023 vin_p.n166 vin_p.t12 321.697
R20024 vin_p.n166 vin_p.t9 321.697
R20025 vin_p.n164 vin_p.t14 321.697
R20026 vin_p.n164 vin_p.t13 321.697
R20027 vin_p.n162 vin_p.t18 321.697
R20028 vin_p.n162 vin_p.t17 321.697
R20029 vin_p.n160 vin_p.t21 321.697
R20030 vin_p.n160 vin_p.t19 321.697
R20031 vin_p.n158 vin_p.t60 321.697
R20032 vin_p.n158 vin_p.t58 321.697
R20033 vin_p.n156 vin_p.t124 321.697
R20034 vin_p.n156 vin_p.t121 321.697
R20035 vin_p.n154 vin_p.t132 321.697
R20036 vin_p.n154 vin_p.t129 321.697
R20037 vin_p.n152 vin_p.t138 321.697
R20038 vin_p.n152 vin_p.t135 321.697
R20039 vin_p.n150 vin_p.t142 321.697
R20040 vin_p.n150 vin_p.t139 321.697
R20041 vin_p.n148 vin_p.t194 321.697
R20042 vin_p.n148 vin_p.t193 321.697
R20043 vin_p.n146 vin_p.t70 321.697
R20044 vin_p.n146 vin_p.t69 321.697
R20045 vin_p.n144 vin_p.t75 321.697
R20046 vin_p.n144 vin_p.t71 321.697
R20047 vin_p.n142 vin_p.t54 321.697
R20048 vin_p.n142 vin_p.t51 321.697
R20049 vin_p.n140 vin_p.t64 321.697
R20050 vin_p.n140 vin_p.t61 321.697
R20051 vin_p.n138 vin_p.t106 321.697
R20052 vin_p.n138 vin_p.t105 321.697
R20053 vin_p.n136 vin_p.t114 321.697
R20054 vin_p.n136 vin_p.t111 321.697
R20055 vin_p.n134 vin_p.t186 321.697
R20056 vin_p.n134 vin_p.t184 321.697
R20057 vin_p.n132 vin_p.t192 321.697
R20058 vin_p.n132 vin_p.t187 321.697
R20059 vin_p.n130 vin_p.t198 321.697
R20060 vin_p.n130 vin_p.t195 321.697
R20061 vin_p.n128 vin_p.t48 321.697
R20062 vin_p.n128 vin_p.t47 321.697
R20063 vin_p.n126 vin_p.t59 321.697
R20064 vin_p.n126 vin_p.t57 321.697
R20065 vin_p.n124 vin_p.t100 321.697
R20066 vin_p.n124 vin_p.t99 321.697
R20067 vin_p.n122 vin_p.t104 321.697
R20068 vin_p.n122 vin_p.t102 321.697
R20069 vin_p.n120 vin_p.t110 321.697
R20070 vin_p.n120 vin_p.t108 321.697
R20071 vin_p.n118 vin_p.t162 321.697
R20072 vin_p.n118 vin_p.t161 321.697
R20073 vin_p.n116 vin_p.t168 321.697
R20074 vin_p.n116 vin_p.t165 321.697
R20075 vin_p.n114 vin_p.t178 321.697
R20076 vin_p.n114 vin_p.t173 321.697
R20077 vin_p.n112 vin_p.t44 321.697
R20078 vin_p.n112 vin_p.t42 321.697
R20079 vin_p.n110 vin_p.t53 321.697
R20080 vin_p.n110 vin_p.t50 321.697
R20081 vin_p.n108 vin_p.t118 321.697
R20082 vin_p.n108 vin_p.t117 321.697
R20083 vin_p.n106 vin_p.t126 321.697
R20084 vin_p.n106 vin_p.t125 321.697
R20085 vin_p.n104 vin_p.t134 321.697
R20086 vin_p.n104 vin_p.t133 321.697
R20087 vin_p.n102 vin_p.t3 321.697
R20088 vin_p.n102 vin_p.t1 321.697
R20089 vin_p.n100 vin_p.t8 321.697
R20090 vin_p.n100 vin_p.t7 321.697
R20091 vin_p.n99 vin_p.t68 321.697
R20092 vin_p.n99 vin_p.t67 321.697
R20093 vin_p.n97 vin_p.t155 321.697
R20094 vin_p.n97 vin_p.t154 321.697
R20095 vin_p.n95 vin_p.t159 321.697
R20096 vin_p.n95 vin_p.t158 321.697
R20097 vin_p.n93 vin_p.t145 321.697
R20098 vin_p.n93 vin_p.t144 321.697
R20099 vin_p.n91 vin_p.t16 321.697
R20100 vin_p.n91 vin_p.t15 321.697
R20101 vin_p.n89 vin_p.t74 321.697
R20102 vin_p.n89 vin_p.t73 321.697
R20103 vin_p.n87 vin_p.t79 321.697
R20104 vin_p.n87 vin_p.t78 321.697
R20105 vin_p.n85 vin_p.t83 321.697
R20106 vin_p.n85 vin_p.t82 321.697
R20107 vin_p.n83 vin_p.t87 321.697
R20108 vin_p.n83 vin_p.t86 321.697
R20109 vin_p.n81 vin_p.t152 321.697
R20110 vin_p.n81 vin_p.t151 321.697
R20111 vin_p.n79 vin_p.t11 321.697
R20112 vin_p.n79 vin_p.t10 321.697
R20113 vin_p.n77 vin_p.t190 321.697
R20114 vin_p.n77 vin_p.t189 321.697
R20115 vin_p.n75 vin_p.t197 321.697
R20116 vin_p.n75 vin_p.t196 321.697
R20117 vin_p.n73 vin_p.t0 321.697
R20118 vin_p.n73 vin_p.t199 321.697
R20119 vin_p.n71 vin_p.t4 321.697
R20120 vin_p.n71 vin_p.t2 321.697
R20121 vin_p.n69 vin_p.t123 321.697
R20122 vin_p.n69 vin_p.t122 321.697
R20123 vin_p.n67 vin_p.t131 321.697
R20124 vin_p.n67 vin_p.t130 321.697
R20125 vin_p.n65 vin_p.t137 321.697
R20126 vin_p.n65 vin_p.t136 321.697
R20127 vin_p.n63 vin_p.t141 321.697
R20128 vin_p.n63 vin_p.t140 321.697
R20129 vin_p.n61 vin_p.t146 321.697
R20130 vin_p.n61 vin_p.t143 321.697
R20131 vin_p.n59 vin_p.t176 321.697
R20132 vin_p.n59 vin_p.t175 321.697
R20133 vin_p.n57 vin_p.t43 321.697
R20134 vin_p.n57 vin_p.t41 321.697
R20135 vin_p.n55 vin_p.t52 321.697
R20136 vin_p.n55 vin_p.t49 321.697
R20137 vin_p.n53 vin_p.t63 321.697
R20138 vin_p.n53 vin_p.t62 321.697
R20139 vin_p.n51 vin_p.t66 321.697
R20140 vin_p.n51 vin_p.t65 321.697
R20141 vin_p.n49 vin_p.t113 321.697
R20142 vin_p.n49 vin_p.t112 321.697
R20143 vin_p.n47 vin_p.t185 321.697
R20144 vin_p.n47 vin_p.t183 321.697
R20145 vin_p.n45 vin_p.t191 321.697
R20146 vin_p.n45 vin_p.t188 321.697
R20147 vin_p.n43 vin_p.t171 321.697
R20148 vin_p.n43 vin_p.t169 321.697
R20149 vin_p.n41 vin_p.t180 321.697
R20150 vin_p.n41 vin_p.t179 321.697
R20151 vin_p.n39 vin_p.t28 321.697
R20152 vin_p.n39 vin_p.t27 321.697
R20153 vin_p.n37 vin_p.t35 321.697
R20154 vin_p.n37 vin_p.t33 321.697
R20155 vin_p.n35 vin_p.t103 321.697
R20156 vin_p.n35 vin_p.t101 321.697
R20157 vin_p.n33 vin_p.t109 321.697
R20158 vin_p.n33 vin_p.t107 321.697
R20159 vin_p.n31 vin_p.t116 321.697
R20160 vin_p.n31 vin_p.t115 321.697
R20161 vin_p.n29 vin_p.t167 321.697
R20162 vin_p.n29 vin_p.t166 321.697
R20163 vin_p.n27 vin_p.t177 321.697
R20164 vin_p.n27 vin_p.t174 321.697
R20165 vin_p.n25 vin_p.t24 321.697
R20166 vin_p.n25 vin_p.t23 321.697
R20167 vin_p.n23 vin_p.t26 321.697
R20168 vin_p.n23 vin_p.t25 321.697
R20169 vin_p.n21 vin_p.t32 321.697
R20170 vin_p.n21 vin_p.t30 321.697
R20171 vin_p.n19 vin_p.t91 321.697
R20172 vin_p.n19 vin_p.t89 321.697
R20173 vin_p.n17 vin_p.t94 321.697
R20174 vin_p.n17 vin_p.t93 321.697
R20175 vin_p.n15 vin_p.t98 321.697
R20176 vin_p.n15 vin_p.t97 321.697
R20177 vin_p.n13 vin_p.t164 321.697
R20178 vin_p.n13 vin_p.t163 321.697
R20179 vin_p.n11 vin_p.t172 321.697
R20180 vin_p.n11 vin_p.t170 321.697
R20181 vin_p.n9 vin_p.t40 321.697
R20182 vin_p.n9 vin_p.t39 321.697
R20183 vin_p.n7 vin_p.t46 321.697
R20184 vin_p.n7 vin_p.t45 321.697
R20185 vin_p.n5 vin_p.t56 321.697
R20186 vin_p.n5 vin_p.t55 321.697
R20187 vin_p.n3 vin_p.t120 321.697
R20188 vin_p.n3 vin_p.t119 321.697
R20189 vin_p.n1 vin_p.t128 321.697
R20190 vin_p.n1 vin_p.t127 321.697
R20191 vin_p.n0 vin_p.t182 321.697
R20192 vin_p.n0 vin_p.t181 321.697
R20193 vin_p.n101 vin_p.n99 67.1865
R20194 vin_p.n2 vin_p.n0 67.1865
R20195 vin_p.n197 vin_p.n196 67.0982
R20196 vin_p.n195 vin_p.n194 67.0982
R20197 vin_p.n193 vin_p.n192 67.0982
R20198 vin_p.n191 vin_p.n190 67.0982
R20199 vin_p.n189 vin_p.n188 67.0982
R20200 vin_p.n187 vin_p.n186 67.0982
R20201 vin_p.n185 vin_p.n184 67.0982
R20202 vin_p.n183 vin_p.n182 67.0982
R20203 vin_p.n181 vin_p.n180 67.0982
R20204 vin_p.n179 vin_p.n178 67.0982
R20205 vin_p.n177 vin_p.n176 67.0982
R20206 vin_p.n175 vin_p.n174 67.0982
R20207 vin_p.n173 vin_p.n172 67.0982
R20208 vin_p.n171 vin_p.n170 67.0982
R20209 vin_p.n169 vin_p.n168 67.0982
R20210 vin_p.n167 vin_p.n166 67.0982
R20211 vin_p.n165 vin_p.n164 67.0982
R20212 vin_p.n163 vin_p.n162 67.0982
R20213 vin_p.n161 vin_p.n160 67.0982
R20214 vin_p.n159 vin_p.n158 67.0982
R20215 vin_p.n157 vin_p.n156 67.0982
R20216 vin_p.n155 vin_p.n154 67.0982
R20217 vin_p.n153 vin_p.n152 67.0982
R20218 vin_p.n151 vin_p.n150 67.0982
R20219 vin_p.n149 vin_p.n148 67.0982
R20220 vin_p.n147 vin_p.n146 67.0982
R20221 vin_p.n145 vin_p.n144 67.0982
R20222 vin_p.n143 vin_p.n142 67.0982
R20223 vin_p.n141 vin_p.n140 67.0982
R20224 vin_p.n139 vin_p.n138 67.0982
R20225 vin_p.n137 vin_p.n136 67.0982
R20226 vin_p.n135 vin_p.n134 67.0982
R20227 vin_p.n133 vin_p.n132 67.0982
R20228 vin_p.n131 vin_p.n130 67.0982
R20229 vin_p.n129 vin_p.n128 67.0982
R20230 vin_p.n127 vin_p.n126 67.0982
R20231 vin_p.n125 vin_p.n124 67.0982
R20232 vin_p.n123 vin_p.n122 67.0982
R20233 vin_p.n121 vin_p.n120 67.0982
R20234 vin_p.n119 vin_p.n118 67.0982
R20235 vin_p.n117 vin_p.n116 67.0982
R20236 vin_p.n115 vin_p.n114 67.0982
R20237 vin_p.n113 vin_p.n112 67.0982
R20238 vin_p.n111 vin_p.n110 67.0982
R20239 vin_p.n109 vin_p.n108 67.0982
R20240 vin_p.n107 vin_p.n106 67.0982
R20241 vin_p.n105 vin_p.n104 67.0982
R20242 vin_p.n103 vin_p.n102 67.0982
R20243 vin_p.n101 vin_p.n100 67.0982
R20244 vin_p.n98 vin_p.n97 67.0982
R20245 vin_p.n96 vin_p.n95 67.0982
R20246 vin_p.n94 vin_p.n93 67.0982
R20247 vin_p.n92 vin_p.n91 67.0982
R20248 vin_p.n90 vin_p.n89 67.0982
R20249 vin_p.n88 vin_p.n87 67.0982
R20250 vin_p.n86 vin_p.n85 67.0982
R20251 vin_p.n84 vin_p.n83 67.0982
R20252 vin_p.n82 vin_p.n81 67.0982
R20253 vin_p.n80 vin_p.n79 67.0982
R20254 vin_p.n78 vin_p.n77 67.0982
R20255 vin_p.n76 vin_p.n75 67.0982
R20256 vin_p.n74 vin_p.n73 67.0982
R20257 vin_p.n72 vin_p.n71 67.0982
R20258 vin_p.n70 vin_p.n69 67.0982
R20259 vin_p.n68 vin_p.n67 67.0982
R20260 vin_p.n66 vin_p.n65 67.0982
R20261 vin_p.n64 vin_p.n63 67.0982
R20262 vin_p.n62 vin_p.n61 67.0982
R20263 vin_p.n60 vin_p.n59 67.0982
R20264 vin_p.n58 vin_p.n57 67.0982
R20265 vin_p.n56 vin_p.n55 67.0982
R20266 vin_p.n54 vin_p.n53 67.0982
R20267 vin_p.n52 vin_p.n51 67.0982
R20268 vin_p.n50 vin_p.n49 67.0982
R20269 vin_p.n48 vin_p.n47 67.0982
R20270 vin_p.n46 vin_p.n45 67.0982
R20271 vin_p.n44 vin_p.n43 67.0982
R20272 vin_p.n42 vin_p.n41 67.0982
R20273 vin_p.n40 vin_p.n39 67.0982
R20274 vin_p.n38 vin_p.n37 67.0982
R20275 vin_p.n36 vin_p.n35 67.0982
R20276 vin_p.n34 vin_p.n33 67.0982
R20277 vin_p.n32 vin_p.n31 67.0982
R20278 vin_p.n30 vin_p.n29 67.0982
R20279 vin_p.n28 vin_p.n27 67.0982
R20280 vin_p.n26 vin_p.n25 67.0982
R20281 vin_p.n24 vin_p.n23 67.0982
R20282 vin_p.n22 vin_p.n21 67.0982
R20283 vin_p.n20 vin_p.n19 67.0982
R20284 vin_p.n18 vin_p.n17 67.0982
R20285 vin_p.n16 vin_p.n15 67.0982
R20286 vin_p.n14 vin_p.n13 67.0982
R20287 vin_p.n12 vin_p.n11 67.0982
R20288 vin_p.n10 vin_p.n9 67.0982
R20289 vin_p.n8 vin_p.n7 67.0982
R20290 vin_p.n6 vin_p.n5 67.0982
R20291 vin_p.n4 vin_p.n3 67.0982
R20292 vin_p.n2 vin_p.n1 67.0982
R20293 vin_p.n198 vin_p.n98 1.1048
R20294 vin_p.n198 vin_p.n197 1.10318
R20295 vin_p vin_p.n198 0.59929
R20296 vin_p.n103 vin_p.n101 0.0888234
R20297 vin_p.n105 vin_p.n103 0.0888234
R20298 vin_p.n107 vin_p.n105 0.0888234
R20299 vin_p.n109 vin_p.n107 0.0888234
R20300 vin_p.n111 vin_p.n109 0.0888234
R20301 vin_p.n113 vin_p.n111 0.0888234
R20302 vin_p.n115 vin_p.n113 0.0888234
R20303 vin_p.n117 vin_p.n115 0.0888234
R20304 vin_p.n119 vin_p.n117 0.0888234
R20305 vin_p.n121 vin_p.n119 0.0888234
R20306 vin_p.n123 vin_p.n121 0.0888234
R20307 vin_p.n125 vin_p.n123 0.0888234
R20308 vin_p.n127 vin_p.n125 0.0888234
R20309 vin_p.n129 vin_p.n127 0.0888234
R20310 vin_p.n131 vin_p.n129 0.0888234
R20311 vin_p.n133 vin_p.n131 0.0888234
R20312 vin_p.n135 vin_p.n133 0.0888234
R20313 vin_p.n137 vin_p.n135 0.0888234
R20314 vin_p.n139 vin_p.n137 0.0888234
R20315 vin_p.n141 vin_p.n139 0.0888234
R20316 vin_p.n143 vin_p.n141 0.0888234
R20317 vin_p.n145 vin_p.n143 0.0888234
R20318 vin_p.n147 vin_p.n145 0.0888234
R20319 vin_p.n149 vin_p.n147 0.0888234
R20320 vin_p.n151 vin_p.n149 0.0888234
R20321 vin_p.n153 vin_p.n151 0.0888234
R20322 vin_p.n155 vin_p.n153 0.0888234
R20323 vin_p.n157 vin_p.n155 0.0888234
R20324 vin_p.n159 vin_p.n157 0.0888234
R20325 vin_p.n161 vin_p.n159 0.0888234
R20326 vin_p.n163 vin_p.n161 0.0888234
R20327 vin_p.n165 vin_p.n163 0.0888234
R20328 vin_p.n167 vin_p.n165 0.0888234
R20329 vin_p.n169 vin_p.n167 0.0888234
R20330 vin_p.n171 vin_p.n169 0.0888234
R20331 vin_p.n173 vin_p.n171 0.0888234
R20332 vin_p.n175 vin_p.n173 0.0888234
R20333 vin_p.n177 vin_p.n175 0.0888234
R20334 vin_p.n179 vin_p.n177 0.0888234
R20335 vin_p.n181 vin_p.n179 0.0888234
R20336 vin_p.n183 vin_p.n181 0.0888234
R20337 vin_p.n185 vin_p.n183 0.0888234
R20338 vin_p.n187 vin_p.n185 0.0888234
R20339 vin_p.n189 vin_p.n187 0.0888234
R20340 vin_p.n191 vin_p.n189 0.0888234
R20341 vin_p.n193 vin_p.n191 0.0888234
R20342 vin_p.n4 vin_p.n2 0.0888234
R20343 vin_p.n6 vin_p.n4 0.0888234
R20344 vin_p.n8 vin_p.n6 0.0888234
R20345 vin_p.n10 vin_p.n8 0.0888234
R20346 vin_p.n12 vin_p.n10 0.0888234
R20347 vin_p.n14 vin_p.n12 0.0888234
R20348 vin_p.n16 vin_p.n14 0.0888234
R20349 vin_p.n18 vin_p.n16 0.0888234
R20350 vin_p.n20 vin_p.n18 0.0888234
R20351 vin_p.n22 vin_p.n20 0.0888234
R20352 vin_p.n24 vin_p.n22 0.0888234
R20353 vin_p.n26 vin_p.n24 0.0888234
R20354 vin_p.n28 vin_p.n26 0.0888234
R20355 vin_p.n30 vin_p.n28 0.0888234
R20356 vin_p.n32 vin_p.n30 0.0888234
R20357 vin_p.n34 vin_p.n32 0.0888234
R20358 vin_p.n36 vin_p.n34 0.0888234
R20359 vin_p.n38 vin_p.n36 0.0888234
R20360 vin_p.n40 vin_p.n38 0.0888234
R20361 vin_p.n42 vin_p.n40 0.0888234
R20362 vin_p.n44 vin_p.n42 0.0888234
R20363 vin_p.n46 vin_p.n44 0.0888234
R20364 vin_p.n48 vin_p.n46 0.0888234
R20365 vin_p.n50 vin_p.n48 0.0888234
R20366 vin_p.n52 vin_p.n50 0.0888234
R20367 vin_p.n54 vin_p.n52 0.0888234
R20368 vin_p.n56 vin_p.n54 0.0888234
R20369 vin_p.n58 vin_p.n56 0.0888234
R20370 vin_p.n60 vin_p.n58 0.0888234
R20371 vin_p.n62 vin_p.n60 0.0888234
R20372 vin_p.n64 vin_p.n62 0.0888234
R20373 vin_p.n66 vin_p.n64 0.0888234
R20374 vin_p.n68 vin_p.n66 0.0888234
R20375 vin_p.n70 vin_p.n68 0.0888234
R20376 vin_p.n72 vin_p.n70 0.0888234
R20377 vin_p.n74 vin_p.n72 0.0888234
R20378 vin_p.n76 vin_p.n74 0.0888234
R20379 vin_p.n78 vin_p.n76 0.0888234
R20380 vin_p.n80 vin_p.n78 0.0888234
R20381 vin_p.n82 vin_p.n80 0.0888234
R20382 vin_p.n84 vin_p.n82 0.0888234
R20383 vin_p.n86 vin_p.n84 0.0888234
R20384 vin_p.n88 vin_p.n86 0.0888234
R20385 vin_p.n90 vin_p.n88 0.0888234
R20386 vin_p.n92 vin_p.n90 0.0888234
R20387 vin_p.n94 vin_p.n92 0.0888234
R20388 vin_p.n96 vin_p.n94 0.0888234
R20389 vin_p.n98 vin_p.n96 0.0888234
R20390 vin_p.n195 vin_p.n193 0.088712
R20391 vin_p.n197 vin_p.n195 0.0882976
R20392 iref.n206 iref.t14 455.844
R20393 iref.n208 iref.t24 455.844
R20394 iref.n205 iref.t18 455.844
R20395 iref.n203 iref.t0 455.844
R20396 iref.n202 iref.t8 455.844
R20397 iref.n200 iref.t16 455.844
R20398 iref.n199 iref.t4 455.844
R20399 iref.n197 iref.t6 455.844
R20400 iref.n196 iref.t20 455.844
R20401 iref.n194 iref.t26 455.844
R20402 iref.n193 iref.t10 455.844
R20403 iref.n191 iref.t22 455.844
R20404 iref.n190 iref.t12 455.844
R20405 iref.n188 iref.t2 455.844
R20406 iref.n187 iref.t28 455.844
R20407 iref.n185 iref.t203 455.844
R20408 iref.n184 iref.t145 455.844
R20409 iref.n183 iref.t149 455.844
R20410 iref.n182 iref.t175 455.844
R20411 iref.n181 iref.t112 455.844
R20412 iref.n180 iref.t55 455.844
R20413 iref.n179 iref.t178 455.844
R20414 iref.n178 iref.t115 455.844
R20415 iref.n177 iref.t186 455.844
R20416 iref.n176 iref.t83 455.844
R20417 iref.n175 iref.t85 455.844
R20418 iref.n174 iref.t207 455.844
R20419 iref.n173 iref.t153 455.844
R20420 iref.n172 iref.t36 455.844
R20421 iref.n171 iref.t119 455.844
R20422 iref.n170 iref.t80 455.844
R20423 iref.n169 iref.t204 455.844
R20424 iref.n168 iref.t156 455.844
R20425 iref.n167 iref.t51 455.844
R20426 iref.n166 iref.t176 455.844
R20427 iref.n165 iref.t113 455.844
R20428 iref.n164 iref.t56 455.844
R20429 iref.n163 iref.t129 455.844
R20430 iref.n162 iref.t67 455.844
R20431 iref.n161 iref.t150 455.844
R20432 iref.n160 iref.t109 455.844
R20433 iref.n159 iref.t52 455.844
R20434 iref.n158 iref.t126 455.844
R20435 iref.n157 iref.t65 455.844
R20436 iref.n156 iref.t147 455.844
R20437 iref.n154 iref.t95 451.39
R20438 iref.n154 iref.t155 451.39
R20439 iref.n152 iref.t37 451.39
R20440 iref.n152 iref.t92 451.39
R20441 iref.n150 iref.t159 451.39
R20442 iref.n150 iref.t31 451.39
R20443 iref.n148 iref.t59 451.39
R20444 iref.n148 iref.t110 451.39
R20445 iref.n146 iref.t191 451.39
R20446 iref.n146 iref.t66 451.39
R20447 iref.n144 iref.t132 451.39
R20448 iref.n144 iref.t184 451.39
R20449 iref.n142 iref.t72 451.39
R20450 iref.n142 iref.t130 451.39
R20451 iref.n140 iref.t194 451.39
R20452 iref.n140 iref.t69 451.39
R20453 iref.n138 iref.t135 451.39
R20454 iref.n138 iref.t187 451.39
R20455 iref.n136 iref.t163 451.39
R20456 iref.n136 iref.t32 451.39
R20457 iref.n134 iref.t98 451.39
R20458 iref.n134 iref.t157 451.39
R20459 iref.n132 iref.t41 451.39
R20460 iref.n132 iref.t93 451.39
R20461 iref.n130 iref.t165 451.39
R20462 iref.n130 iref.t34 451.39
R20463 iref.n128 iref.t168 451.39
R20464 iref.n128 iref.t38 451.39
R20465 iref.n126 iref.t60 451.39
R20466 iref.n126 iref.t118 451.39
R20467 iref.n124 iref.t136 451.39
R20468 iref.n124 iref.t189 451.39
R20469 iref.n122 iref.t75 451.39
R20470 iref.n122 iref.t131 451.39
R20471 iref.n120 iref.t198 451.39
R20472 iref.n120 iref.t71 451.39
R20473 iref.n118 iref.t142 451.39
R20474 iref.n118 iref.t192 451.39
R20475 iref.n116 iref.t209 451.39
R20476 iref.n116 iref.t87 451.39
R20477 iref.n114 iref.t104 451.39
R20478 iref.n114 iref.t161 451.39
R20479 iref.n112 iref.t106 451.39
R20480 iref.n112 iref.t164 451.39
R20481 iref.n110 iref.t50 451.39
R20482 iref.n110 iref.t99 451.39
R20483 iref.n108 iref.t174 451.39
R20484 iref.n108 iref.t42 451.39
R20485 iref.n106 iref.t64 451.39
R20486 iref.n106 iref.t122 451.39
R20487 iref.n104 iref.t100 451.39
R20488 iref.n104 iref.t158 451.39
R20489 iref.n102 iref.t44 451.39
R20490 iref.n102 iref.t94 451.39
R20491 iref.n100 iref.t123 451.39
R20492 iref.n100 iref.t180 451.39
R20493 iref.n98 iref.t125 451.39
R20494 iref.n98 iref.t182 451.39
R20495 iref.n96 iref.t62 451.39
R20496 iref.n96 iref.t120 451.39
R20497 iref.n94 iref.t140 451.39
R20498 iref.n94 iref.t190 451.39
R20499 iref.n92 iref.t77 451.39
R20500 iref.n92 iref.t133 451.39
R20501 iref.n90 iref.t200 451.39
R20502 iref.n90 iref.t73 451.39
R20503 iref.n88 iref.t91 451.39
R20504 iref.n88 iref.t154 451.39
R20505 iref.n86 iref.t30 451.39
R20506 iref.n86 iref.t88 451.39
R20507 iref.n84 iref.t105 451.39
R20508 iref.n84 iref.t162 451.39
R20509 iref.n82 iref.t48 451.39
R20510 iref.n82 iref.t97 451.39
R20511 iref.n80 iref.t53 451.39
R20512 iref.n80 iref.t101 451.39
R20513 iref.n78 iref.t128 451.39
R20514 iref.n78 iref.t183 451.39
R20515 iref.n76 iref.t68 451.39
R20516 iref.n76 iref.t124 451.39
R20517 iref.n74 iref.t146 451.39
R20518 iref.n74 iref.t196 451.39
R20519 iref.n72 iref.t81 451.39
R20520 iref.n72 iref.t137 451.39
R20521 iref.n70 iref.t205 451.39
R20522 iref.n70 iref.t76 451.39
R20523 iref.n68 iref.t151 451.39
R20524 iref.n68 iref.t199 451.39
R20525 iref.n66 iref.t33 451.39
R20526 iref.n66 iref.t89 451.39
R20527 iref.n64 iref.t179 451.39
R20528 iref.n64 iref.t46 451.39
R20529 iref.n62 iref.t116 451.39
R20530 iref.n62 iref.t170 451.39
R20531 iref.n60 iref.t57 451.39
R20532 iref.n60 iref.t107 451.39
R20533 iref.n58 iref.t181 451.39
R20534 iref.n58 iref.t49 451.39
R20535 iref.n56 iref.t70 451.39
R20536 iref.n56 iref.t127 451.39
R20537 iref.n54 iref.t138 451.39
R20538 iref.n54 iref.t188 451.39
R20539 iref.n52 iref.t208 451.39
R20540 iref.n52 iref.t86 451.39
R20541 iref.n50 iref.t167 451.39
R20542 iref.n50 iref.t39 451.39
R20543 iref.n48 iref.t103 451.39
R20544 iref.n48 iref.t160 451.39
R20545 iref.n46 iref.t47 451.39
R20546 iref.n46 iref.t96 451.39
R20547 iref.n44 iref.t171 451.39
R20548 iref.n44 iref.t40 451.39
R20549 iref.n42 iref.t63 451.39
R20550 iref.n42 iref.t121 451.39
R20551 iref.n40 iref.t141 451.39
R20552 iref.n40 iref.t193 451.39
R20553 iref.n38 iref.t78 451.39
R20554 iref.n38 iref.t134 451.39
R20555 iref.n36 iref.t201 451.39
R20556 iref.n36 iref.t74 451.39
R20557 iref.n34 iref.t144 451.39
R20558 iref.n34 iref.t195 451.39
R20559 iref.n32 iref.t148 451.39
R20560 iref.n32 iref.t197 451.39
R20561 iref.n30 iref.t173 451.39
R20562 iref.n30 iref.t43 451.39
R20563 iref.n28 iref.t111 451.39
R20564 iref.n28 iref.t166 451.39
R20565 iref.n26 iref.t54 451.39
R20566 iref.n26 iref.t102 451.39
R20567 iref.n24 iref.t177 451.39
R20568 iref.n24 iref.t45 451.39
R20569 iref.n22 iref.t114 451.39
R20570 iref.n22 iref.t169 451.39
R20571 iref.n20 iref.t185 451.39
R20572 iref.n20 iref.t61 451.39
R20573 iref.n18 iref.t82 451.39
R20574 iref.n18 iref.t139 451.39
R20575 iref.n16 iref.t84 451.39
R20576 iref.n16 iref.t143 451.39
R20577 iref.n14 iref.t206 451.39
R20578 iref.n14 iref.t79 451.39
R20579 iref.n12 iref.t152 451.39
R20580 iref.n12 iref.t202 451.39
R20581 iref.n10 iref.t35 451.39
R20582 iref.n10 iref.t90 451.39
R20583 iref.n8 iref.t117 451.39
R20584 iref.n8 iref.t172 451.39
R20585 iref.n7 iref.t58 451.39
R20586 iref.n7 iref.t108 451.39
R20587 iref.n186 iref.t29 85.1726
R20588 iref.n189 iref.n6 75.651
R20589 iref.n192 iref.n5 75.651
R20590 iref.n195 iref.n4 75.651
R20591 iref.n198 iref.n3 75.651
R20592 iref.n201 iref.n2 75.651
R20593 iref.n204 iref.n1 75.651
R20594 iref.n207 iref.n0 75.651
R20595 iref.n6 iref.t3 9.52217
R20596 iref.n6 iref.t13 9.52217
R20597 iref.n5 iref.t23 9.52217
R20598 iref.n5 iref.t11 9.52217
R20599 iref.n4 iref.t27 9.52217
R20600 iref.n4 iref.t21 9.52217
R20601 iref.n3 iref.t7 9.52217
R20602 iref.n3 iref.t5 9.52217
R20603 iref.n2 iref.t17 9.52217
R20604 iref.n2 iref.t9 9.52217
R20605 iref.n1 iref.t1 9.52217
R20606 iref.n1 iref.t19 9.52217
R20607 iref.n0 iref.t15 9.52217
R20608 iref.n0 iref.t25 9.52217
R20609 iref.n9 iref.n7 2.33576
R20610 iref.n9 iref.n8 2.2505
R20611 iref.n11 iref.n10 2.2505
R20612 iref.n13 iref.n12 2.2505
R20613 iref.n15 iref.n14 2.2505
R20614 iref.n17 iref.n16 2.2505
R20615 iref.n19 iref.n18 2.2505
R20616 iref.n21 iref.n20 2.2505
R20617 iref.n23 iref.n22 2.2505
R20618 iref.n25 iref.n24 2.2505
R20619 iref.n27 iref.n26 2.2505
R20620 iref.n29 iref.n28 2.2505
R20621 iref.n31 iref.n30 2.2505
R20622 iref.n33 iref.n32 2.2505
R20623 iref.n35 iref.n34 2.2505
R20624 iref.n37 iref.n36 2.2505
R20625 iref.n39 iref.n38 2.2505
R20626 iref.n41 iref.n40 2.2505
R20627 iref.n43 iref.n42 2.2505
R20628 iref.n45 iref.n44 2.2505
R20629 iref.n47 iref.n46 2.2505
R20630 iref.n49 iref.n48 2.2505
R20631 iref.n51 iref.n50 2.2505
R20632 iref.n53 iref.n52 2.2505
R20633 iref.n55 iref.n54 2.2505
R20634 iref.n57 iref.n56 2.2505
R20635 iref.n59 iref.n58 2.2505
R20636 iref.n61 iref.n60 2.2505
R20637 iref.n63 iref.n62 2.2505
R20638 iref.n65 iref.n64 2.2505
R20639 iref.n67 iref.n66 2.2505
R20640 iref.n69 iref.n68 2.2505
R20641 iref.n71 iref.n70 2.2505
R20642 iref.n73 iref.n72 2.2505
R20643 iref.n75 iref.n74 2.2505
R20644 iref.n77 iref.n76 2.2505
R20645 iref.n79 iref.n78 2.2505
R20646 iref.n81 iref.n80 2.2505
R20647 iref.n83 iref.n82 2.2505
R20648 iref.n85 iref.n84 2.2505
R20649 iref.n87 iref.n86 2.2505
R20650 iref.n89 iref.n88 2.2505
R20651 iref.n91 iref.n90 2.2505
R20652 iref.n93 iref.n92 2.2505
R20653 iref.n95 iref.n94 2.2505
R20654 iref.n97 iref.n96 2.2505
R20655 iref.n99 iref.n98 2.2505
R20656 iref.n101 iref.n100 2.2505
R20657 iref.n103 iref.n102 2.2505
R20658 iref.n105 iref.n104 2.2505
R20659 iref.n107 iref.n106 2.2505
R20660 iref.n109 iref.n108 2.2505
R20661 iref.n111 iref.n110 2.2505
R20662 iref.n113 iref.n112 2.2505
R20663 iref.n115 iref.n114 2.2505
R20664 iref.n117 iref.n116 2.2505
R20665 iref.n119 iref.n118 2.2505
R20666 iref.n121 iref.n120 2.2505
R20667 iref.n123 iref.n122 2.2505
R20668 iref.n125 iref.n124 2.2505
R20669 iref.n127 iref.n126 2.2505
R20670 iref.n129 iref.n128 2.2505
R20671 iref.n131 iref.n130 2.2505
R20672 iref.n133 iref.n132 2.2505
R20673 iref.n135 iref.n134 2.2505
R20674 iref.n137 iref.n136 2.2505
R20675 iref.n139 iref.n138 2.2505
R20676 iref.n141 iref.n140 2.2505
R20677 iref.n143 iref.n142 2.2505
R20678 iref.n145 iref.n144 2.2505
R20679 iref.n147 iref.n146 2.2505
R20680 iref.n149 iref.n148 2.2505
R20681 iref.n151 iref.n150 2.2505
R20682 iref.n153 iref.n152 2.2505
R20683 iref.n155 iref.n154 2.2505
R20684 iref iref.n208 2.0359
R20685 iref.n156 iref.n155 1.47593
R20686 iref.n57 iref.n55 0.933303
R20687 iref.n107 iref.n105 0.933303
R20688 iref.n171 iref.n170 0.2505
R20689 iref.n186 iref.n185 0.20787
R20690 iref.n11 iref.n9 0.0857601
R20691 iref.n13 iref.n11 0.0857601
R20692 iref.n15 iref.n13 0.0857601
R20693 iref.n17 iref.n15 0.0857601
R20694 iref.n19 iref.n17 0.0857601
R20695 iref.n21 iref.n19 0.0857601
R20696 iref.n23 iref.n21 0.0857601
R20697 iref.n25 iref.n23 0.0857601
R20698 iref.n27 iref.n25 0.0857601
R20699 iref.n29 iref.n27 0.0857601
R20700 iref.n31 iref.n29 0.0857601
R20701 iref.n33 iref.n31 0.0857601
R20702 iref.n35 iref.n33 0.0857601
R20703 iref.n37 iref.n35 0.0857601
R20704 iref.n39 iref.n37 0.0857601
R20705 iref.n41 iref.n39 0.0857601
R20706 iref.n43 iref.n41 0.0857601
R20707 iref.n45 iref.n43 0.0857601
R20708 iref.n47 iref.n45 0.0857601
R20709 iref.n49 iref.n47 0.0857601
R20710 iref.n51 iref.n49 0.0857601
R20711 iref.n53 iref.n51 0.0857601
R20712 iref.n55 iref.n53 0.0857601
R20713 iref.n59 iref.n57 0.0857601
R20714 iref.n61 iref.n59 0.0857601
R20715 iref.n63 iref.n61 0.0857601
R20716 iref.n65 iref.n63 0.0857601
R20717 iref.n67 iref.n65 0.0857601
R20718 iref.n69 iref.n67 0.0857601
R20719 iref.n71 iref.n69 0.0857601
R20720 iref.n73 iref.n71 0.0857601
R20721 iref.n75 iref.n73 0.0857601
R20722 iref.n77 iref.n75 0.0857601
R20723 iref.n79 iref.n77 0.0857601
R20724 iref.n81 iref.n79 0.0857601
R20725 iref.n83 iref.n81 0.0857601
R20726 iref.n85 iref.n83 0.0857601
R20727 iref.n87 iref.n85 0.0857601
R20728 iref.n89 iref.n87 0.0857601
R20729 iref.n91 iref.n89 0.0857601
R20730 iref.n93 iref.n91 0.0857601
R20731 iref.n95 iref.n93 0.0857601
R20732 iref.n97 iref.n95 0.0857601
R20733 iref.n99 iref.n97 0.0857601
R20734 iref.n101 iref.n99 0.0857601
R20735 iref.n103 iref.n101 0.0857601
R20736 iref.n105 iref.n103 0.0857601
R20737 iref.n109 iref.n107 0.0857601
R20738 iref.n111 iref.n109 0.0857601
R20739 iref.n113 iref.n111 0.0857601
R20740 iref.n115 iref.n113 0.0857601
R20741 iref.n117 iref.n115 0.0857601
R20742 iref.n119 iref.n117 0.0857601
R20743 iref.n121 iref.n119 0.0857601
R20744 iref.n123 iref.n121 0.0857601
R20745 iref.n125 iref.n123 0.0857601
R20746 iref.n127 iref.n125 0.0857601
R20747 iref.n129 iref.n127 0.0857601
R20748 iref.n131 iref.n129 0.0857601
R20749 iref.n133 iref.n131 0.0857601
R20750 iref.n135 iref.n133 0.0857601
R20751 iref.n137 iref.n135 0.0857601
R20752 iref.n139 iref.n137 0.0857601
R20753 iref.n141 iref.n139 0.0857601
R20754 iref.n143 iref.n141 0.0857601
R20755 iref.n145 iref.n143 0.0857601
R20756 iref.n147 iref.n145 0.0857601
R20757 iref.n149 iref.n147 0.0857601
R20758 iref.n151 iref.n149 0.0857601
R20759 iref.n153 iref.n151 0.0857601
R20760 iref.n155 iref.n153 0.0857601
R20761 iref.n157 iref.n156 0.0857601
R20762 iref.n158 iref.n157 0.0857601
R20763 iref.n159 iref.n158 0.0857601
R20764 iref.n160 iref.n159 0.0857601
R20765 iref.n161 iref.n160 0.0857601
R20766 iref.n162 iref.n161 0.0857601
R20767 iref.n163 iref.n162 0.0857601
R20768 iref.n164 iref.n163 0.0857601
R20769 iref.n165 iref.n164 0.0857601
R20770 iref.n166 iref.n165 0.0857601
R20771 iref.n167 iref.n166 0.0857601
R20772 iref.n168 iref.n167 0.0857601
R20773 iref.n169 iref.n168 0.0857601
R20774 iref.n170 iref.n169 0.0857601
R20775 iref.n172 iref.n171 0.0857601
R20776 iref.n173 iref.n172 0.0857601
R20777 iref.n174 iref.n173 0.0857601
R20778 iref.n175 iref.n174 0.0857601
R20779 iref.n176 iref.n175 0.0857601
R20780 iref.n177 iref.n176 0.0857601
R20781 iref.n178 iref.n177 0.0857601
R20782 iref.n179 iref.n178 0.0857601
R20783 iref.n180 iref.n179 0.0857601
R20784 iref.n181 iref.n180 0.0857601
R20785 iref.n182 iref.n181 0.0857601
R20786 iref.n183 iref.n182 0.0857601
R20787 iref.n184 iref.n183 0.0857601
R20788 iref.n185 iref.n184 0.0857601
R20789 iref.n188 iref.n187 0.0857601
R20790 iref.n191 iref.n190 0.0857601
R20791 iref.n194 iref.n193 0.0857601
R20792 iref.n197 iref.n196 0.0857601
R20793 iref.n200 iref.n199 0.0857601
R20794 iref.n203 iref.n202 0.0857601
R20795 iref.n206 iref.n205 0.0857601
R20796 iref.n187 iref.n186 0.0431301
R20797 iref.n189 iref.n188 0.0431301
R20798 iref.n190 iref.n189 0.0431301
R20799 iref.n192 iref.n191 0.0431301
R20800 iref.n193 iref.n192 0.0431301
R20801 iref.n195 iref.n194 0.0431301
R20802 iref.n196 iref.n195 0.0431301
R20803 iref.n198 iref.n197 0.0431301
R20804 iref.n199 iref.n198 0.0431301
R20805 iref.n201 iref.n200 0.0431301
R20806 iref.n202 iref.n201 0.0431301
R20807 iref.n204 iref.n203 0.0431301
R20808 iref.n205 iref.n204 0.0431301
R20809 iref.n207 iref.n206 0.0431301
R20810 iref.n208 iref.n207 0.0431301
R20811 vdd.n2321 vdd.n312 21667.1
R20812 vdd.n1512 vdd.n311 21667.1
R20813 vdd.n2323 vdd.n238 8668.24
R20814 vdd.n2483 vdd.n238 8668.24
R20815 vdd.n2483 vdd.n239 8668.24
R20816 vdd.n2323 vdd.n239 8668.24
R20817 vdd.n1300 vdd.n308 8668.24
R20818 vdd.n2326 vdd.n308 8668.24
R20819 vdd.n1300 vdd.n309 8668.24
R20820 vdd.n2326 vdd.n309 8668.24
R20821 vdd.n1161 vdd.n618 8668.24
R20822 vdd.n1509 vdd.n618 8668.24
R20823 vdd.n1509 vdd.n619 8668.24
R20824 vdd.n1161 vdd.n619 8668.24
R20825 vdd.n2567 vdd.n237 5110.59
R20826 vdd.n2566 vdd.n237 5110.59
R20827 vdd.n2814 vdd.n136 5110.59
R20828 vdd.n2813 vdd.n136 5110.59
R20829 vdd.n2567 vdd.n144 3525.88
R20830 vdd.n2806 vdd.n144 3525.88
R20831 vdd.n2806 vdd.n135 3525.88
R20832 vdd.n2814 vdd.n135 3525.88
R20833 vdd.n2566 vdd.n140 3525.88
R20834 vdd.n2807 vdd.n140 3525.88
R20835 vdd.n2807 vdd.n137 3525.88
R20836 vdd.n2813 vdd.n137 3525.88
R20837 vdd.n142 vdd.n135 1584.71
R20838 vdd.n142 vdd.n137 1584.71
R20839 vdd.n2487 vdd.n144 1584.71
R20840 vdd.n2487 vdd.n140 1584.71
R20841 vdd.n2485 vdd.n2484 1205.7
R20842 vdd.n2565 vdd.n2564 545.13
R20843 vdd.n2812 vdd.n2811 545.13
R20844 vdd.n1510 vdd.n617 416.204
R20845 vdd.n2325 vdd.n2324 416.204
R20846 vdd.n2565 vdd.n139 376.094
R20847 vdd.n2808 vdd.n139 376.094
R20848 vdd.n2809 vdd.n2808 376.094
R20849 vdd.n2812 vdd.n2809 376.094
R20850 vdd.n2482 vdd.n2481 361.413
R20851 vdd.n2482 vdd.n240 353.507
R20852 vdd.n355 vdd.n294 326.401
R20853 vdd.n2346 vdd.n294 326.401
R20854 vdd.n1301 vdd.n525 326.401
R20855 vdd.n1302 vdd.n1301 326.401
R20856 vdd.n2327 vdd.n307 326.401
R20857 vdd.n2329 vdd.n2327 326.401
R20858 vdd.n1508 vdd.n526 326.401
R20859 vdd.n1508 vdd.n1507 326.401
R20860 vdd.n1162 vdd.n1160 326.401
R20861 vdd.n1163 vdd.n1162 326.401
R20862 vdd.n2179 vdd.t319 251.661
R20863 vdd.n2180 vdd.t318 251.661
R20864 vdd.n2181 vdd.t315 251.154
R20865 vdd.n2181 vdd.t320 251.153
R20866 vdd.n2180 vdd.t316 251.114
R20867 vdd.n2179 vdd.t317 251.114
R20868 vdd.n2811 vdd.n2810 196.142
R20869 vdd.n2685 vdd.n138 169.036
R20870 vdd.n2809 vdd.n138 169.036
R20871 vdd.n2564 vdd.n2563 169.036
R20872 vdd.n2486 vdd.n189 169.036
R20873 vdd.n2486 vdd.n139 169.036
R20874 vdd.t138 vdd.n136 141.232
R20875 vdd.t133 vdd.n2485 124.413
R20876 vdd.t254 vdd.n2488 124.413
R20877 vdd.n2488 vdd.t183 124.413
R20878 vdd.t20 vdd.n143 124.413
R20879 vdd.n143 vdd.t181 124.413
R20880 vdd.n1975 vdd.t227 85.6198
R20881 vdd.n370 vdd.t217 85.6198
R20882 vdd.n537 vdd.t148 85.6198
R20883 vdd.n623 vdd.t51 85.3025
R20884 vdd.n1373 vdd.t111 85.3025
R20885 vdd.n2479 vdd.t119 85.3025
R20886 vdd.n2855 vdd.t139 84.9754
R20887 vdd.n2767 vdd.t21 84.9754
R20888 vdd.n200 vdd.t255 84.9754
R20889 vdd.t269 vdd.t133 84.8605
R20890 vdd.t169 vdd.t269 84.8605
R20891 vdd.t291 vdd.t169 84.8605
R20892 vdd.t203 vdd.t291 84.8605
R20893 vdd.t124 vdd.t203 84.8605
R20894 vdd.t185 vdd.t124 84.8605
R20895 vdd.t164 vdd.t185 84.8605
R20896 vdd.t164 vdd.t281 84.8605
R20897 vdd.t281 vdd.t196 84.8605
R20898 vdd.t196 vdd.t74 84.8605
R20899 vdd.t74 vdd.t293 84.8605
R20900 vdd.t293 vdd.t116 84.8605
R20901 vdd.t116 vdd.t18 84.8605
R20902 vdd.t18 vdd.t254 84.8605
R20903 vdd.t183 vdd.t288 84.8605
R20904 vdd.t288 vdd.t122 84.8605
R20905 vdd.t122 vdd.t8 84.8605
R20906 vdd.t8 vdd.t223 84.8605
R20907 vdd.t223 vdd.t246 84.8605
R20908 vdd.t246 vdd.t4 84.8605
R20909 vdd.t191 vdd.t68 84.8605
R20910 vdd.t68 vdd.t283 84.8605
R20911 vdd.t283 vdd.t198 84.8605
R20912 vdd.t198 vdd.t76 84.8605
R20913 vdd.t76 vdd.t130 84.8605
R20914 vdd.t130 vdd.t136 84.8605
R20915 vdd.t136 vdd.t20 84.8605
R20916 vdd.t181 vdd.t2 84.8605
R20917 vdd.t2 vdd.t241 84.8605
R20918 vdd.t241 vdd.t126 84.8605
R20919 vdd.t126 vdd.t10 84.8605
R20920 vdd.t10 vdd.t14 84.8605
R20921 vdd.t14 vdd.t160 84.8605
R20922 vdd.t278 vdd.t160 84.8605
R20923 vdd.t278 vdd.t193 84.8605
R20924 vdd.t193 vdd.t70 84.8605
R20925 vdd.t70 vdd.t285 84.8605
R20926 vdd.t285 vdd.t112 84.8605
R20927 vdd.t112 vdd.t248 84.8605
R20928 vdd.t248 vdd.t252 84.8605
R20929 vdd.t252 vdd.t138 84.8605
R20930 vdd.n1161 vdd.t205 83.9026
R20931 vdd.t50 vdd.n1510 76.1943
R20932 vdd.n617 vdd.t167 76.1943
R20933 vdd.n2325 vdd.t110 76.1943
R20934 vdd.n2484 vdd.t118 76.1943
R20935 vdd.n460 vdd.n459 76.0981
R20936 vdd.n1119 vdd.n983 76.0981
R20937 vdd.n1970 vdd.n1969 76.0981
R20938 vdd.n1964 vdd.n1963 76.0981
R20939 vdd.n1958 vdd.n1957 76.0981
R20940 vdd.n1952 vdd.n1951 76.0981
R20941 vdd.n1946 vdd.n1945 76.0981
R20942 vdd.n1940 vdd.n1939 76.0981
R20943 vdd.n1934 vdd.n1933 76.0981
R20944 vdd.n1929 vdd.n1928 76.0981
R20945 vdd.n2295 vdd.n1923 76.0981
R20946 vdd.n2301 vdd.n1918 76.0981
R20947 vdd.n336 vdd.n335 76.0981
R20948 vdd.n1911 vdd.n338 76.0981
R20949 vdd.n1748 vdd.n1747 76.0981
R20950 vdd.n1745 vdd.n1744 76.0981
R20951 vdd.n1742 vdd.n1741 76.0981
R20952 vdd.n1739 vdd.n1738 76.0981
R20953 vdd.n1737 vdd.n1736 76.0981
R20954 vdd.n1779 vdd.n1733 76.0981
R20955 vdd.n1785 vdd.n1730 76.0981
R20956 vdd.n1725 vdd.n1724 76.0981
R20957 vdd.n480 vdd.n479 76.0981
R20958 vdd.n493 vdd.n492 76.0981
R20959 vdd.n1665 vdd.n1664 76.0981
R20960 vdd.n551 vdd.n550 76.0981
R20961 vdd.n564 vdd.n563 76.0981
R20962 vdd.n585 vdd.n584 76.0981
R20963 vdd.n588 vdd.n587 76.0981
R20964 vdd.n1526 vdd.n1525 76.0981
R20965 vdd.n979 vdd.n978 76.0981
R20966 vdd.n973 vdd.n972 76.0981
R20967 vdd.n967 vdd.n966 76.0981
R20968 vdd.n961 vdd.n960 76.0981
R20969 vdd.n955 vdd.n954 76.0981
R20970 vdd.n706 vdd.n705 76.0981
R20971 vdd.n1263 vdd.n637 75.7808
R20972 vdd.n1176 vdd.n682 75.7808
R20973 vdd.n1185 vdd.n677 75.7808
R20974 vdd.n1196 vdd.n672 75.7808
R20975 vdd.n1205 vdd.n667 75.7808
R20976 vdd.n1214 vdd.n662 75.7808
R20977 vdd.n1225 vdd.n657 75.7808
R20978 vdd.n1235 vdd.n652 75.7808
R20979 vdd.n1244 vdd.n647 75.7808
R20980 vdd.n1255 vdd.n642 75.7808
R20981 vdd.n633 vdd.n632 75.7808
R20982 vdd.n628 vdd.n627 75.7808
R20983 vdd.n1482 vdd.n1305 75.7808
R20984 vdd.n1473 vdd.n1311 75.7808
R20985 vdd.n1464 vdd.n1316 75.7808
R20986 vdd.n1454 vdd.n1321 75.7808
R20987 vdd.n1445 vdd.n1327 75.7808
R20988 vdd.n1436 vdd.n1332 75.7808
R20989 vdd.n1341 vdd.n1339 75.7808
R20990 vdd.n1347 vdd.n1346 75.7808
R20991 vdd.n1353 vdd.n1352 75.7808
R20992 vdd.n1360 vdd.n1359 75.7808
R20993 vdd.n1366 vdd.n1365 75.7808
R20994 vdd.n1372 vdd.n1371 75.7808
R20995 vdd.n2352 vdd.n2351 75.7808
R20996 vdd.n2364 vdd.n2363 75.7808
R20997 vdd.n2374 vdd.n2373 75.7808
R20998 vdd.n2384 vdd.n2383 75.7808
R20999 vdd.n2396 vdd.n2395 75.7808
R21000 vdd.n2406 vdd.n2405 75.7808
R21001 vdd.n2417 vdd.n2416 75.7808
R21002 vdd.n2429 vdd.n2428 75.7808
R21003 vdd.n2439 vdd.n2438 75.7808
R21004 vdd.n2449 vdd.n2448 75.7808
R21005 vdd.n2461 vdd.n2460 75.7808
R21006 vdd.n2470 vdd.n247 75.7808
R21007 vdd.n2722 vdd.n2721 75.5775
R21008 vdd.n2697 vdd.n2696 75.5775
R21009 vdd.n2631 vdd.n170 75.4538
R21010 vdd.n2845 vdd.n2844 75.4538
R21011 vdd.n117 vdd.n116 75.4538
R21012 vdd.n125 vdd.n124 75.4538
R21013 vdd.n2734 vdd.n2733 75.4538
R21014 vdd.n2705 vdd.n2704 75.4538
R21015 vdd.n2778 vdd.n2777 75.4538
R21016 vdd.n2789 vdd.n2788 75.4538
R21017 vdd.n2656 vdd.n2655 75.4538
R21018 vdd.n151 vdd.n150 75.4538
R21019 vdd.n162 vdd.n161 75.4538
R21020 vdd.n182 vdd.n181 75.4538
R21021 vdd.n206 vdd.n205 75.4538
R21022 vdd.n215 vdd.n214 75.4538
R21023 vdd.n2580 vdd.n2579 75.4538
R21024 vdd.n234 vdd.n233 75.4538
R21025 vdd.n2534 vdd.n2520 75.4538
R21026 vdd.n2545 vdd.n2544 75.4538
R21027 vdd.n2502 vdd.n2501 75.4538
R21028 vdd.n899 vdd.n814 62.1255
R21029 vdd.n466 vdd.n449 61.7417
R21030 vdd.n1797 vdd.n452 61.3652
R21031 vdd.n457 vdd.n454 61.3652
R21032 vdd.n1795 vdd.n1794 61.3652
R21033 vdd.t205 vdd.t82 51.9708
R21034 vdd.t82 vdd.t235 51.9708
R21035 vdd.t235 vdd.t22 51.9708
R21036 vdd.t22 vdd.t12 51.9708
R21037 vdd.t12 vdd.t141 51.9708
R21038 vdd.t141 vdd.t146 51.9708
R21039 vdd.t146 vdd.t54 51.9708
R21040 vdd.t54 vdd.t88 51.9708
R21041 vdd.t88 vdd.t72 51.9708
R21042 vdd.t72 vdd.t213 51.9708
R21043 vdd.t213 vdd.t94 51.9708
R21044 vdd.t94 vdd.t80 51.9708
R21045 vdd.t80 vdd.t32 51.9708
R21046 vdd.t32 vdd.t36 51.9708
R21047 vdd.t36 vdd.t24 51.9708
R21048 vdd.t24 vdd.t153 51.9708
R21049 vdd.t153 vdd.t40 51.9708
R21050 vdd.t177 vdd.t84 51.9708
R21051 vdd.t84 vdd.t225 51.9708
R21052 vdd.t225 vdd.t106 51.9708
R21053 vdd.t106 vdd.t92 51.9708
R21054 vdd.t92 vdd.t6 51.9708
R21055 vdd.t6 vdd.t50 51.9708
R21056 vdd.t167 vdd.t62 51.9708
R21057 vdd.t62 vdd.t207 51.9708
R21058 vdd.t207 vdd.t86 51.9708
R21059 vdd.t86 vdd.t66 51.9708
R21060 vdd.t66 vdd.t237 51.9708
R21061 vdd.t237 vdd.t28 51.9708
R21062 vdd.t28 vdd.t16 51.9708
R21063 vdd.t16 vdd.t149 51.9708
R21064 vdd.t149 vdd.t34 51.9708
R21065 vdd.t34 vdd.t172 51.9708
R21066 vdd.t172 vdd.t58 51.9708
R21067 vdd.t58 vdd.t215 51.9708
R21068 vdd.t215 vdd.t221 51.9708
R21069 vdd.t221 vdd.t102 51.9708
R21070 vdd.t102 vdd.t239 51.9708
R21071 vdd.t239 vdd.t120 51.9708
R21072 vdd.t120 vdd.t26 51.9708
R21073 vdd.t26 vdd.t155 51.9708
R21074 vdd.t155 vdd.t46 51.9708
R21075 vdd.t46 vdd.t179 51.9708
R21076 vdd.t179 vdd.t60 51.9708
R21077 vdd.t60 vdd.t64 51.9708
R21078 vdd.t64 vdd.t228 51.9708
R21079 vdd.t228 vdd.t110 51.9708
R21080 vdd.t175 vdd.t78 51.9708
R21081 vdd.t78 vdd.t218 51.9708
R21082 vdd.t218 vdd.t98 51.9708
R21083 vdd.t98 vdd.t104 51.9708
R21084 vdd.t104 vdd.t0 51.9708
R21085 vdd.t0 vdd.t42 51.9708
R21086 vdd.t42 vdd.t30 51.9708
R21087 vdd.t30 vdd.t158 51.9708
R21088 vdd.t158 vdd.t48 51.9708
R21089 vdd.t48 vdd.t187 51.9708
R21090 vdd.t187 vdd.t90 51.9708
R21091 vdd.t90 vdd.t96 51.9708
R21092 vdd.t96 vdd.t230 51.9708
R21093 vdd.t230 vdd.t114 51.9708
R21094 vdd.t114 vdd.t100 51.9708
R21095 vdd.t100 vdd.t52 51.9708
R21096 vdd.t52 vdd.t38 51.9708
R21097 vdd.t38 vdd.t162 51.9708
R21098 vdd.t162 vdd.t56 51.9708
R21099 vdd.t56 vdd.t44 51.9708
R21100 vdd.t44 vdd.t201 51.9708
R21101 vdd.t201 vdd.t108 51.9708
R21102 vdd.t108 vdd.t232 51.9708
R21103 vdd.t232 vdd.t118 51.9708
R21104 vdd.n2324 vdd.n2322 50.2091
R21105 vdd.t191 vdd.n141 48.1837
R21106 vdd.n899 vdd.n815 44.0005
R21107 vdd.n860 vdd.n841 41.7614
R21108 vdd.n875 vdd.n874 41.7614
R21109 vdd.n839 vdd.n835 41.7614
R21110 vdd.n881 vdd.n880 41.7614
R21111 vdd.n833 vdd.n829 41.7614
R21112 vdd.n887 vdd.n886 41.7614
R21113 vdd.n827 vdd.n820 41.7614
R21114 vdd.n893 vdd.n892 41.7614
R21115 vdd.n821 vdd.n816 41.7614
R21116 vdd.n898 vdd.n750 41.7614
R21117 vdd.n751 vdd.n747 41.7614
R21118 vdd.n906 vdd.n905 41.7614
R21119 vdd.n745 vdd.n742 41.7614
R21120 vdd.n744 vdd.n739 41.7614
R21121 vdd.n912 vdd.n911 41.7614
R21122 vdd.n737 vdd.n733 41.7614
R21123 vdd.n918 vdd.n917 41.7614
R21124 vdd.n731 vdd.n727 41.7614
R21125 vdd.n924 vdd.n923 41.7614
R21126 vdd.n755 vdd.n724 41.7614
R21127 vdd.t4 vdd.n141 36.6773
R21128 vdd.n2158 vdd.n2157 36.4064
R21129 vdd.n2158 vdd.n1977 36.4064
R21130 vdd.n2158 vdd.n1978 36.4064
R21131 vdd.n2560 vdd.n2490 36.4064
R21132 vdd.n2853 vdd.n97 36.4064
R21133 vdd.n2492 vdd.n2490 36.4064
R21134 vdd.n99 vdd.n97 36.4064
R21135 vdd.n2494 vdd.n2490 36.4064
R21136 vdd.n101 vdd.n97 36.4064
R21137 vdd.n868 vdd.n844 36.4064
R21138 vdd.n809 vdd.n762 34.5151
R21139 vdd.n774 vdd.n758 34.5141
R21140 vdd.n773 vdd.n760 34.5141
R21141 vdd.n813 vdd.n812 34.5141
R21142 vdd.n1506 vdd.n621 34.4388
R21143 vdd.n1658 vdd.n1657 34.4388
R21144 vdd.n1654 vdd.n1653 34.4388
R21145 vdd.n1634 vdd.n530 34.4388
R21146 vdd.n1639 vdd.n528 34.4388
R21147 vdd.n357 vdd.n356 34.4388
R21148 vdd.n1898 vdd.n1897 34.4388
R21149 vdd.n365 vdd.n354 34.4388
R21150 vdd.n1901 vdd.n1900 34.4388
R21151 vdd.n2345 vdd.n295 34.4338
R21152 vdd.n2328 vdd.n295 34.4289
R21153 vdd.n1639 vdd.n1638 34.4289
R21154 vdd.n1902 vdd.n1901 34.4289
R21155 vdd.n1635 vdd.n1634 34.4289
R21156 vdd.n365 vdd.n343 34.4289
R21157 vdd.n1653 vdd.n509 34.4289
R21158 vdd.n1897 vdd.n350 34.4289
R21159 vdd.n1511 vdd.t177 33.4729
R21160 vdd.n1302 vdd.n621 31.4171
R21161 vdd.n1658 vdd.n525 31.0406
R21162 vdd.n356 vdd.n355 30.6642
R21163 vdd.n2563 vdd.n2490 29.6299
R21164 vdd.n764 vdd.n758 27.1064
R21165 vdd.n785 vdd.n764 27.1064
R21166 vdd.n794 vdd.n785 27.1064
R21167 vdd.n795 vdd.n794 27.1064
R21168 vdd.n795 vdd.n718 27.1064
R21169 vdd.n718 vdd.n714 27.1064
R21170 vdd.n714 vdd.n713 27.1064
R21171 vdd.n713 vdd.n710 27.1064
R21172 vdd.n710 vdd.n693 27.1064
R21173 vdd.n698 vdd.n693 27.1064
R21174 vdd.n702 vdd.n698 27.1064
R21175 vdd.n1053 vdd.n702 27.1064
R21176 vdd.n1054 vdd.n1053 27.1064
R21177 vdd.n1054 vdd.n1028 27.1064
R21178 vdd.n1062 vdd.n1028 27.1064
R21179 vdd.n1063 vdd.n1062 27.1064
R21180 vdd.n1063 vdd.n1022 27.1064
R21181 vdd.n1071 vdd.n1022 27.1064
R21182 vdd.n1072 vdd.n1071 27.1064
R21183 vdd.n1072 vdd.n1016 27.1064
R21184 vdd.n1080 vdd.n1016 27.1064
R21185 vdd.n1081 vdd.n1080 27.1064
R21186 vdd.n1081 vdd.n1010 27.1064
R21187 vdd.n1089 vdd.n1010 27.1064
R21188 vdd.n1090 vdd.n1089 27.1064
R21189 vdd.n1090 vdd.n1004 27.1064
R21190 vdd.n1098 vdd.n1004 27.1064
R21191 vdd.n1099 vdd.n1098 27.1064
R21192 vdd.n1099 vdd.n1001 27.1064
R21193 vdd.n1001 vdd.n993 27.1064
R21194 vdd.n993 vdd.n992 27.1064
R21195 vdd.n992 vdd.n991 27.1064
R21196 vdd.n991 vdd.n990 27.1064
R21197 vdd.n990 vdd.n989 27.1064
R21198 vdd.n989 vdd.n609 27.1064
R21199 vdd.n609 vdd.n608 27.1064
R21200 vdd.n608 vdd.n607 27.1064
R21201 vdd.n607 vdd.n606 27.1064
R21202 vdd.n606 vdd.n605 27.1064
R21203 vdd.n582 vdd.n578 27.1064
R21204 vdd.n578 vdd.n573 27.1064
R21205 vdd.n573 vdd.n572 27.1064
R21206 vdd.n572 vdd.n571 27.1064
R21207 vdd.n571 vdd.n562 27.1064
R21208 vdd.n562 vdd.n558 27.1064
R21209 vdd.n558 vdd.n555 27.1064
R21210 vdd.n555 vdd.n549 27.1064
R21211 vdd.n549 vdd.n545 27.1064
R21212 vdd.n545 vdd.n542 27.1064
R21213 vdd.n542 vdd.n536 27.1064
R21214 vdd.n536 vdd.n533 27.1064
R21215 vdd.n533 vdd.n528 27.1064
R21216 vdd.n1638 vdd.n506 27.1064
R21217 vdd.n1676 vdd.n506 27.1064
R21218 vdd.n1677 vdd.n1676 27.1064
R21219 vdd.n1677 vdd.n498 27.1064
R21220 vdd.n1686 vdd.n498 27.1064
R21221 vdd.n1687 vdd.n1686 27.1064
R21222 vdd.n1687 vdd.n485 27.1064
R21223 vdd.n1699 vdd.n485 27.1064
R21224 vdd.n1700 vdd.n1699 27.1064
R21225 vdd.n1700 vdd.n469 27.1064
R21226 vdd.n1714 vdd.n469 27.1064
R21227 vdd.n1715 vdd.n1714 27.1064
R21228 vdd.n1716 vdd.n1715 27.1064
R21229 vdd.n1717 vdd.n1716 27.1064
R21230 vdd.n1717 vdd.n452 27.1064
R21231 vdd.n1798 vdd.n1797 27.1064
R21232 vdd.n1798 vdd.n443 27.1064
R21233 vdd.n1806 vdd.n443 27.1064
R21234 vdd.n1807 vdd.n1806 27.1064
R21235 vdd.n1807 vdd.n434 27.1064
R21236 vdd.n1816 vdd.n434 27.1064
R21237 vdd.n1817 vdd.n1816 27.1064
R21238 vdd.n1817 vdd.n424 27.1064
R21239 vdd.n1823 vdd.n424 27.1064
R21240 vdd.n1824 vdd.n1823 27.1064
R21241 vdd.n1824 vdd.n415 27.1064
R21242 vdd.n1832 vdd.n415 27.1064
R21243 vdd.n1833 vdd.n1832 27.1064
R21244 vdd.n1833 vdd.n406 27.1064
R21245 vdd.n1841 vdd.n406 27.1064
R21246 vdd.n1842 vdd.n1841 27.1064
R21247 vdd.n1842 vdd.n396 27.1064
R21248 vdd.n1848 vdd.n396 27.1064
R21249 vdd.n1849 vdd.n1848 27.1064
R21250 vdd.n1849 vdd.n387 27.1064
R21251 vdd.n1857 vdd.n387 27.1064
R21252 vdd.n1858 vdd.n1857 27.1064
R21253 vdd.n1858 vdd.n377 27.1064
R21254 vdd.n1866 vdd.n377 27.1064
R21255 vdd.n1867 vdd.n1866 27.1064
R21256 vdd.n1867 vdd.n352 27.1064
R21257 vdd.n1900 vdd.n352 27.1064
R21258 vdd.n1902 vdd.n313 27.1064
R21259 vdd.n2319 vdd.n314 27.1064
R21260 vdd.n2313 vdd.n314 27.1064
R21261 vdd.n2313 vdd.n2312 27.1064
R21262 vdd.n2312 vdd.n326 27.1064
R21263 vdd.n2059 vdd.n326 27.1064
R21264 vdd.n2060 vdd.n2059 27.1064
R21265 vdd.n2060 vdd.n2052 27.1064
R21266 vdd.n2068 vdd.n2052 27.1064
R21267 vdd.n2069 vdd.n2068 27.1064
R21268 vdd.n2069 vdd.n2043 27.1064
R21269 vdd.n2075 vdd.n2043 27.1064
R21270 vdd.n2076 vdd.n2075 27.1064
R21271 vdd.n2076 vdd.n2036 27.1064
R21272 vdd.n2084 vdd.n2036 27.1064
R21273 vdd.n2085 vdd.n2084 27.1064
R21274 vdd.n2085 vdd.n2030 27.1064
R21275 vdd.n2093 vdd.n2030 27.1064
R21276 vdd.n2094 vdd.n2093 27.1064
R21277 vdd.n2094 vdd.n2021 27.1064
R21278 vdd.n2100 vdd.n2021 27.1064
R21279 vdd.n2101 vdd.n2100 27.1064
R21280 vdd.n2101 vdd.n2015 27.1064
R21281 vdd.n2109 vdd.n2015 27.1064
R21282 vdd.n2110 vdd.n2109 27.1064
R21283 vdd.n2110 vdd.n2009 27.1064
R21284 vdd.n2118 vdd.n2009 27.1064
R21285 vdd.n2120 vdd.n2118 27.1064
R21286 vdd.n2120 vdd.n2119 27.1064
R21287 vdd.n2119 vdd.n2000 27.1064
R21288 vdd.n2129 vdd.n2000 27.1064
R21289 vdd.n2130 vdd.n2129 27.1064
R21290 vdd.n2130 vdd.n1994 27.1064
R21291 vdd.n2138 vdd.n1994 27.1064
R21292 vdd.n2139 vdd.n2138 27.1064
R21293 vdd.n2139 vdd.n1985 27.1064
R21294 vdd.n2147 vdd.n1985 27.1064
R21295 vdd.n2148 vdd.n2147 27.1064
R21296 vdd.n2149 vdd.n2148 27.1064
R21297 vdd.n2149 vdd.n1979 27.1064
R21298 vdd.n2157 vdd.n1979 27.1064
R21299 vdd.n806 vdd.n760 27.1064
R21300 vdd.n806 vdd.n805 27.1064
R21301 vdd.n805 vdd.n783 27.1064
R21302 vdd.n797 vdd.n783 27.1064
R21303 vdd.n797 vdd.n711 27.1064
R21304 vdd.n940 vdd.n711 27.1064
R21305 vdd.n941 vdd.n940 27.1064
R21306 vdd.n942 vdd.n941 27.1064
R21307 vdd.n942 vdd.n695 27.1064
R21308 vdd.n1153 vdd.n695 27.1064
R21309 vdd.n1153 vdd.n1152 27.1064
R21310 vdd.n1152 vdd.n700 27.1064
R21311 vdd.n1056 vdd.n700 27.1064
R21312 vdd.n1057 vdd.n1056 27.1064
R21313 vdd.n1057 vdd.n1026 27.1064
R21314 vdd.n1065 vdd.n1026 27.1064
R21315 vdd.n1066 vdd.n1065 27.1064
R21316 vdd.n1066 vdd.n1020 27.1064
R21317 vdd.n1074 vdd.n1020 27.1064
R21318 vdd.n1075 vdd.n1074 27.1064
R21319 vdd.n1075 vdd.n1014 27.1064
R21320 vdd.n1083 vdd.n1014 27.1064
R21321 vdd.n1084 vdd.n1083 27.1064
R21322 vdd.n1084 vdd.n1008 27.1064
R21323 vdd.n1092 vdd.n1008 27.1064
R21324 vdd.n1093 vdd.n1092 27.1064
R21325 vdd.n1093 vdd.n1002 27.1064
R21326 vdd.n1101 vdd.n1002 27.1064
R21327 vdd.n1102 vdd.n1101 27.1064
R21328 vdd.n1102 vdd.n998 27.1064
R21329 vdd.n998 vdd.n997 27.1064
R21330 vdd.n997 vdd.n996 27.1064
R21331 vdd.n996 vdd.n995 27.1064
R21332 vdd.n995 vdd.n994 27.1064
R21333 vdd.n994 vdd.n615 27.1064
R21334 vdd.n615 vdd.n614 27.1064
R21335 vdd.n614 vdd.n613 27.1064
R21336 vdd.n613 vdd.n612 27.1064
R21337 vdd.n612 vdd.n611 27.1064
R21338 vdd.n1551 vdd.n1550 27.1064
R21339 vdd.n1551 vdd.n575 27.1064
R21340 vdd.n575 vdd.n574 27.1064
R21341 vdd.n574 vdd.n560 27.1064
R21342 vdd.n1578 vdd.n560 27.1064
R21343 vdd.n1579 vdd.n1578 27.1064
R21344 vdd.n1579 vdd.n547 27.1064
R21345 vdd.n1591 vdd.n547 27.1064
R21346 vdd.n1592 vdd.n1591 27.1064
R21347 vdd.n1592 vdd.n534 27.1064
R21348 vdd.n1649 vdd.n534 27.1064
R21349 vdd.n1650 vdd.n1649 27.1064
R21350 vdd.n1650 vdd.n530 27.1064
R21351 vdd.n1635 vdd.n511 27.1064
R21352 vdd.n511 vdd.n503 27.1064
R21353 vdd.n1679 vdd.n503 27.1064
R21354 vdd.n1680 vdd.n1679 27.1064
R21355 vdd.n1680 vdd.n500 27.1064
R21356 vdd.n500 vdd.n497 27.1064
R21357 vdd.n497 vdd.n491 27.1064
R21358 vdd.n491 vdd.n487 27.1064
R21359 vdd.n487 vdd.n484 27.1064
R21360 vdd.n484 vdd.n478 27.1064
R21361 vdd.n478 vdd.n473 27.1064
R21362 vdd.n473 vdd.n472 27.1064
R21363 vdd.n472 vdd.n471 27.1064
R21364 vdd.n471 vdd.n468 27.1064
R21365 vdd.n468 vdd.n457 27.1064
R21366 vdd.n454 vdd.n451 27.1064
R21367 vdd.n451 vdd.n448 27.1064
R21368 vdd.n448 vdd.n445 27.1064
R21369 vdd.n445 vdd.n442 27.1064
R21370 vdd.n442 vdd.n439 27.1064
R21371 vdd.n439 vdd.n436 27.1064
R21372 vdd.n436 vdd.n430 27.1064
R21373 vdd.n430 vdd.n429 27.1064
R21374 vdd.n429 vdd.n426 27.1064
R21375 vdd.n426 vdd.n423 27.1064
R21376 vdd.n423 vdd.n420 27.1064
R21377 vdd.n420 vdd.n417 27.1064
R21378 vdd.n417 vdd.n414 27.1064
R21379 vdd.n414 vdd.n411 27.1064
R21380 vdd.n411 vdd.n408 27.1064
R21381 vdd.n408 vdd.n402 27.1064
R21382 vdd.n402 vdd.n401 27.1064
R21383 vdd.n401 vdd.n398 27.1064
R21384 vdd.n398 vdd.n395 27.1064
R21385 vdd.n395 vdd.n392 27.1064
R21386 vdd.n392 vdd.n389 27.1064
R21387 vdd.n389 vdd.n386 27.1064
R21388 vdd.n386 vdd.n383 27.1064
R21389 vdd.n383 vdd.n379 27.1064
R21390 vdd.n379 vdd.n373 27.1064
R21391 vdd.n373 vdd.n372 27.1064
R21392 vdd.n372 vdd.n354 27.1064
R21393 vdd.n346 vdd.n343 27.1064
R21394 vdd.n321 vdd.n316 27.1064
R21395 vdd.n323 vdd.n321 27.1064
R21396 vdd.n327 vdd.n323 27.1064
R21397 vdd.n331 vdd.n327 27.1064
R21398 vdd.n2057 vdd.n331 27.1064
R21399 vdd.n2058 vdd.n2057 27.1064
R21400 vdd.n2058 vdd.n2055 27.1064
R21401 vdd.n2055 vdd.n2053 27.1064
R21402 vdd.n2053 vdd.n2049 27.1064
R21403 vdd.n2049 vdd.n2048 27.1064
R21404 vdd.n2048 vdd.n2045 27.1064
R21405 vdd.n2045 vdd.n2042 27.1064
R21406 vdd.n2042 vdd.n2040 27.1064
R21407 vdd.n2040 vdd.n2038 27.1064
R21408 vdd.n2038 vdd.n2035 27.1064
R21409 vdd.n2035 vdd.n2033 27.1064
R21410 vdd.n2033 vdd.n2031 27.1064
R21411 vdd.n2031 vdd.n2026 27.1064
R21412 vdd.n2026 vdd.n2025 27.1064
R21413 vdd.n2025 vdd.n2023 27.1064
R21414 vdd.n2023 vdd.n2020 27.1064
R21415 vdd.n2020 vdd.n2018 27.1064
R21416 vdd.n2018 vdd.n2016 27.1064
R21417 vdd.n2016 vdd.n2014 27.1064
R21418 vdd.n2014 vdd.n2012 27.1064
R21419 vdd.n2012 vdd.n2010 27.1064
R21420 vdd.n2010 vdd.n2007 27.1064
R21421 vdd.n2007 vdd.n2006 27.1064
R21422 vdd.n2006 vdd.n2004 27.1064
R21423 vdd.n2004 vdd.n2001 27.1064
R21424 vdd.n2001 vdd.n1999 27.1064
R21425 vdd.n1999 vdd.n1997 27.1064
R21426 vdd.n1997 vdd.n1995 27.1064
R21427 vdd.n1995 vdd.n1993 27.1064
R21428 vdd.n1993 vdd.n1991 27.1064
R21429 vdd.n1991 vdd.n1987 27.1064
R21430 vdd.n1987 vdd.n1986 27.1064
R21431 vdd.n1986 vdd.n1984 27.1064
R21432 vdd.n1984 vdd.n1981 27.1064
R21433 vdd.n1981 vdd.n1977 27.1064
R21434 vdd.n809 vdd.n808 27.1064
R21435 vdd.n808 vdd.n763 27.1064
R21436 vdd.n786 vdd.n763 27.1064
R21437 vdd.n786 vdd.n716 27.1064
R21438 vdd.n936 vdd.n716 27.1064
R21439 vdd.n938 vdd.n936 27.1064
R21440 vdd.n938 vdd.n937 27.1064
R21441 vdd.n937 vdd.n696 27.1064
R21442 vdd.n1156 vdd.n696 27.1064
R21443 vdd.n1156 vdd.n1155 27.1064
R21444 vdd.n1155 vdd.n697 27.1064
R21445 vdd.n1051 vdd.n697 27.1064
R21446 vdd.n1051 vdd.n1030 27.1064
R21447 vdd.n1059 vdd.n1030 27.1064
R21448 vdd.n1060 vdd.n1059 27.1064
R21449 vdd.n1060 vdd.n1024 27.1064
R21450 vdd.n1068 vdd.n1024 27.1064
R21451 vdd.n1069 vdd.n1068 27.1064
R21452 vdd.n1069 vdd.n1018 27.1064
R21453 vdd.n1077 vdd.n1018 27.1064
R21454 vdd.n1078 vdd.n1077 27.1064
R21455 vdd.n1078 vdd.n1012 27.1064
R21456 vdd.n1086 vdd.n1012 27.1064
R21457 vdd.n1087 vdd.n1086 27.1064
R21458 vdd.n1087 vdd.n1006 27.1064
R21459 vdd.n1095 vdd.n1006 27.1064
R21460 vdd.n1096 vdd.n1095 27.1064
R21461 vdd.n1096 vdd.n999 27.1064
R21462 vdd.n1104 vdd.n999 27.1064
R21463 vdd.n1108 vdd.n1104 27.1064
R21464 vdd.n1108 vdd.n1107 27.1064
R21465 vdd.n1107 vdd.n1106 27.1064
R21466 vdd.n1106 vdd.n1105 27.1064
R21467 vdd.n1105 vdd.n616 27.1064
R21468 vdd.n1518 vdd.n616 27.1064
R21469 vdd.n1518 vdd.n1517 27.1064
R21470 vdd.n1517 vdd.n1516 27.1064
R21471 vdd.n1516 vdd.n1515 27.1064
R21472 vdd.n1515 vdd.n1514 27.1064
R21473 vdd.n1553 vdd.n576 27.1064
R21474 vdd.n1556 vdd.n1553 27.1064
R21475 vdd.n1556 vdd.n1555 27.1064
R21476 vdd.n1555 vdd.n1554 27.1064
R21477 vdd.n1554 vdd.n556 27.1064
R21478 vdd.n1581 vdd.n556 27.1064
R21479 vdd.n1582 vdd.n1581 27.1064
R21480 vdd.n1582 vdd.n543 27.1064
R21481 vdd.n1594 vdd.n543 27.1064
R21482 vdd.n1595 vdd.n1594 27.1064
R21483 vdd.n1595 vdd.n531 27.1064
R21484 vdd.n1652 vdd.n531 27.1064
R21485 vdd.n1654 vdd.n1652 27.1064
R21486 vdd.n1673 vdd.n509 27.1064
R21487 vdd.n1674 vdd.n1673 27.1064
R21488 vdd.n1674 vdd.n501 27.1064
R21489 vdd.n1683 vdd.n501 27.1064
R21490 vdd.n1684 vdd.n1683 27.1064
R21491 vdd.n1684 vdd.n489 27.1064
R21492 vdd.n1696 vdd.n489 27.1064
R21493 vdd.n1697 vdd.n1696 27.1064
R21494 vdd.n1697 vdd.n476 27.1064
R21495 vdd.n1709 vdd.n476 27.1064
R21496 vdd.n1712 vdd.n1709 27.1064
R21497 vdd.n1712 vdd.n1711 27.1064
R21498 vdd.n1711 vdd.n1710 27.1064
R21499 vdd.n1710 vdd.n455 27.1064
R21500 vdd.n1794 vdd.n455 27.1064
R21501 vdd.n1795 vdd.n446 27.1064
R21502 vdd.n1803 vdd.n446 27.1064
R21503 vdd.n1804 vdd.n1803 27.1064
R21504 vdd.n1804 vdd.n437 27.1064
R21505 vdd.n1813 vdd.n437 27.1064
R21506 vdd.n1814 vdd.n1813 27.1064
R21507 vdd.n1814 vdd.n433 27.1064
R21508 vdd.n433 vdd.n432 27.1064
R21509 vdd.n432 vdd.n421 27.1064
R21510 vdd.n1826 vdd.n421 27.1064
R21511 vdd.n1827 vdd.n1826 27.1064
R21512 vdd.n1827 vdd.n412 27.1064
R21513 vdd.n1835 vdd.n412 27.1064
R21514 vdd.n1836 vdd.n1835 27.1064
R21515 vdd.n1836 vdd.n399 27.1064
R21516 vdd.n1844 vdd.n399 27.1064
R21517 vdd.n1845 vdd.n1844 27.1064
R21518 vdd.n1846 vdd.n1845 27.1064
R21519 vdd.n1846 vdd.n390 27.1064
R21520 vdd.n1854 vdd.n390 27.1064
R21521 vdd.n1855 vdd.n1854 27.1064
R21522 vdd.n1855 vdd.n381 27.1064
R21523 vdd.n1863 vdd.n381 27.1064
R21524 vdd.n1864 vdd.n1863 27.1064
R21525 vdd.n1864 vdd.n376 27.1064
R21526 vdd.n376 vdd.n359 27.1064
R21527 vdd.n1898 vdd.n359 27.1064
R21528 vdd.n350 vdd.n349 27.1064
R21529 vdd.n2317 vdd.n2316 27.1064
R21530 vdd.n2316 vdd.n320 27.1064
R21531 vdd.n2310 vdd.n320 27.1064
R21532 vdd.n2310 vdd.n2309 27.1064
R21533 vdd.n2309 vdd.n330 27.1064
R21534 vdd.n2054 vdd.n330 27.1064
R21535 vdd.n2065 vdd.n2054 27.1064
R21536 vdd.n2066 vdd.n2065 27.1064
R21537 vdd.n2066 vdd.n2051 27.1064
R21538 vdd.n2051 vdd.n2050 27.1064
R21539 vdd.n2050 vdd.n2041 27.1064
R21540 vdd.n2078 vdd.n2041 27.1064
R21541 vdd.n2079 vdd.n2078 27.1064
R21542 vdd.n2079 vdd.n2034 27.1064
R21543 vdd.n2087 vdd.n2034 27.1064
R21544 vdd.n2088 vdd.n2087 27.1064
R21545 vdd.n2088 vdd.n2024 27.1064
R21546 vdd.n2096 vdd.n2024 27.1064
R21547 vdd.n2097 vdd.n2096 27.1064
R21548 vdd.n2098 vdd.n2097 27.1064
R21549 vdd.n2098 vdd.n2017 27.1064
R21550 vdd.n2106 vdd.n2017 27.1064
R21551 vdd.n2107 vdd.n2106 27.1064
R21552 vdd.n2107 vdd.n2011 27.1064
R21553 vdd.n2115 vdd.n2011 27.1064
R21554 vdd.n2116 vdd.n2115 27.1064
R21555 vdd.n2116 vdd.n2008 27.1064
R21556 vdd.n2008 vdd.n2002 27.1064
R21557 vdd.n2126 vdd.n2002 27.1064
R21558 vdd.n2127 vdd.n2126 27.1064
R21559 vdd.n2127 vdd.n1996 27.1064
R21560 vdd.n2135 vdd.n1996 27.1064
R21561 vdd.n2136 vdd.n2135 27.1064
R21562 vdd.n2136 vdd.n1990 27.1064
R21563 vdd.n2144 vdd.n1990 27.1064
R21564 vdd.n2145 vdd.n2144 27.1064
R21565 vdd.n2145 vdd.n1982 27.1064
R21566 vdd.n2151 vdd.n1982 27.1064
R21567 vdd.n2152 vdd.n2151 27.1064
R21568 vdd.n2152 vdd.n1978 27.1064
R21569 vdd.n2560 vdd.n2559 27.1064
R21570 vdd.n2559 vdd.n2558 27.1064
R21571 vdd.n2558 vdd.n2495 27.1064
R21572 vdd.n2551 vdd.n2495 27.1064
R21573 vdd.n2551 vdd.n2550 27.1064
R21574 vdd.n2550 vdd.n2507 27.1064
R21575 vdd.n2540 vdd.n2507 27.1064
R21576 vdd.n2540 vdd.n2539 27.1064
R21577 vdd.n2539 vdd.n2515 27.1064
R21578 vdd.n2532 vdd.n2515 27.1064
R21579 vdd.n2532 vdd.n2531 27.1064
R21580 vdd.n2531 vdd.n2523 27.1064
R21581 vdd.n2523 vdd.n230 27.1064
R21582 vdd.n2574 vdd.n230 27.1064
R21583 vdd.n2575 vdd.n2574 27.1064
R21584 vdd.n2575 vdd.n220 27.1064
R21585 vdd.n2585 vdd.n220 27.1064
R21586 vdd.n2586 vdd.n2585 27.1064
R21587 vdd.n2587 vdd.n2586 27.1064
R21588 vdd.n2587 vdd.n211 27.1064
R21589 vdd.n2595 vdd.n211 27.1064
R21590 vdd.n2596 vdd.n2595 27.1064
R21591 vdd.n2596 vdd.n202 27.1064
R21592 vdd.n2604 vdd.n202 27.1064
R21593 vdd.n2605 vdd.n2604 27.1064
R21594 vdd.n2605 vdd.n191 27.1064
R21595 vdd.n2611 vdd.n191 27.1064
R21596 vdd.n2612 vdd.n2611 27.1064
R21597 vdd.n2612 vdd.n184 27.1064
R21598 vdd.n2620 vdd.n184 27.1064
R21599 vdd.n2621 vdd.n2620 27.1064
R21600 vdd.n2621 vdd.n176 27.1064
R21601 vdd.n2629 vdd.n176 27.1064
R21602 vdd.n2630 vdd.n2629 27.1064
R21603 vdd.n2630 vdd.n166 27.1064
R21604 vdd.n2636 vdd.n166 27.1064
R21605 vdd.n2637 vdd.n2636 27.1064
R21606 vdd.n2637 vdd.n158 27.1064
R21607 vdd.n2645 vdd.n158 27.1064
R21608 vdd.n2646 vdd.n2645 27.1064
R21609 vdd.n2802 vdd.n2652 27.1064
R21610 vdd.n2802 vdd.n2801 27.1064
R21611 vdd.n2801 vdd.n2653 27.1064
R21612 vdd.n2795 vdd.n2653 27.1064
R21613 vdd.n2795 vdd.n2794 27.1064
R21614 vdd.n2794 vdd.n2663 27.1064
R21615 vdd.n2784 vdd.n2663 27.1064
R21616 vdd.n2784 vdd.n2783 27.1064
R21617 vdd.n2783 vdd.n2671 27.1064
R21618 vdd.n2773 vdd.n2671 27.1064
R21619 vdd.n2773 vdd.n2772 27.1064
R21620 vdd.n2772 vdd.n2677 27.1064
R21621 vdd.n2683 vdd.n2677 27.1064
R21622 vdd.n2686 vdd.n2683 27.1064
R21623 vdd.n2689 vdd.n2686 27.1064
R21624 vdd.n2756 vdd.n2689 27.1064
R21625 vdd.n2756 vdd.n2755 27.1064
R21626 vdd.n2755 vdd.n2694 27.1064
R21627 vdd.n2747 vdd.n2694 27.1064
R21628 vdd.n2747 vdd.n2746 27.1064
R21629 vdd.n2746 vdd.n2702 27.1064
R21630 vdd.n2740 vdd.n2702 27.1064
R21631 vdd.n2740 vdd.n2739 27.1064
R21632 vdd.n2739 vdd.n2712 27.1064
R21633 vdd.n2729 vdd.n2712 27.1064
R21634 vdd.n2729 vdd.n2728 27.1064
R21635 vdd.n2728 vdd.n2720 27.1064
R21636 vdd.n2720 vdd.n130 27.1064
R21637 vdd.n2821 vdd.n130 27.1064
R21638 vdd.n2822 vdd.n2821 27.1064
R21639 vdd.n2822 vdd.n121 27.1064
R21640 vdd.n2830 vdd.n121 27.1064
R21641 vdd.n2831 vdd.n2830 27.1064
R21642 vdd.n2831 vdd.n112 27.1064
R21643 vdd.n2839 vdd.n112 27.1064
R21644 vdd.n2840 vdd.n2839 27.1064
R21645 vdd.n2840 vdd.n102 27.1064
R21646 vdd.n2851 vdd.n102 27.1064
R21647 vdd.n2852 vdd.n2851 27.1064
R21648 vdd.n2853 vdd.n2852 27.1064
R21649 vdd.n2496 vdd.n2492 27.1064
R21650 vdd.n2497 vdd.n2496 27.1064
R21651 vdd.n2503 vdd.n2497 27.1064
R21652 vdd.n2505 vdd.n2503 27.1064
R21653 vdd.n2508 vdd.n2505 27.1064
R21654 vdd.n2511 vdd.n2508 27.1064
R21655 vdd.n2513 vdd.n2511 27.1064
R21656 vdd.n2516 vdd.n2513 27.1064
R21657 vdd.n2518 vdd.n2516 27.1064
R21658 vdd.n2521 vdd.n2518 27.1064
R21659 vdd.n2527 vdd.n2521 27.1064
R21660 vdd.n2527 vdd.n2526 27.1064
R21661 vdd.n2526 vdd.n235 27.1064
R21662 vdd.n235 vdd.n231 27.1064
R21663 vdd.n231 vdd.n229 27.1064
R21664 vdd.n229 vdd.n227 27.1064
R21665 vdd.n227 vdd.n223 27.1064
R21666 vdd.n223 vdd.n222 27.1064
R21667 vdd.n222 vdd.n219 27.1064
R21668 vdd.n219 vdd.n216 27.1064
R21669 vdd.n216 vdd.n212 27.1064
R21670 vdd.n212 vdd.n210 27.1064
R21671 vdd.n210 vdd.n207 27.1064
R21672 vdd.n207 vdd.n203 27.1064
R21673 vdd.n203 vdd.n197 27.1064
R21674 vdd.n197 vdd.n196 27.1064
R21675 vdd.n196 vdd.n193 27.1064
R21676 vdd.n193 vdd.n190 27.1064
R21677 vdd.n190 vdd.n188 27.1064
R21678 vdd.n188 vdd.n185 27.1064
R21679 vdd.n185 vdd.n183 27.1064
R21680 vdd.n183 vdd.n179 27.1064
R21681 vdd.n179 vdd.n177 27.1064
R21682 vdd.n177 vdd.n172 27.1064
R21683 vdd.n172 vdd.n171 27.1064
R21684 vdd.n171 vdd.n168 27.1064
R21685 vdd.n168 vdd.n165 27.1064
R21686 vdd.n165 vdd.n163 27.1064
R21687 vdd.n163 vdd.n159 27.1064
R21688 vdd.n159 vdd.n156 27.1064
R21689 vdd.n152 vdd.n147 27.1064
R21690 vdd.n2654 vdd.n147 27.1064
R21691 vdd.n2659 vdd.n2654 27.1064
R21692 vdd.n2661 vdd.n2659 27.1064
R21693 vdd.n2664 vdd.n2661 27.1064
R21694 vdd.n2667 vdd.n2664 27.1064
R21695 vdd.n2669 vdd.n2667 27.1064
R21696 vdd.n2672 vdd.n2669 27.1064
R21697 vdd.n2674 vdd.n2672 27.1064
R21698 vdd.n2676 vdd.n2674 27.1064
R21699 vdd.n2678 vdd.n2676 27.1064
R21700 vdd.n2681 vdd.n2678 27.1064
R21701 vdd.n2684 vdd.n2681 27.1064
R21702 vdd.n2762 vdd.n2684 27.1064
R21703 vdd.n2762 vdd.n2761 27.1064
R21704 vdd.n2761 vdd.n2688 27.1064
R21705 vdd.n2695 vdd.n2688 27.1064
R21706 vdd.n2699 vdd.n2695 27.1064
R21707 vdd.n2701 vdd.n2699 27.1064
R21708 vdd.n2703 vdd.n2701 27.1064
R21709 vdd.n2708 vdd.n2703 27.1064
R21710 vdd.n2710 vdd.n2708 27.1064
R21711 vdd.n2713 vdd.n2710 27.1064
R21712 vdd.n2716 vdd.n2713 27.1064
R21713 vdd.n2718 vdd.n2716 27.1064
R21714 vdd.n2725 vdd.n2718 27.1064
R21715 vdd.n2725 vdd.n2724 27.1064
R21716 vdd.n2724 vdd.n133 27.1064
R21717 vdd.n133 vdd.n131 27.1064
R21718 vdd.n131 vdd.n129 27.1064
R21719 vdd.n129 vdd.n126 27.1064
R21720 vdd.n126 vdd.n122 27.1064
R21721 vdd.n122 vdd.n120 27.1064
R21722 vdd.n120 vdd.n118 27.1064
R21723 vdd.n118 vdd.n114 27.1064
R21724 vdd.n114 vdd.n111 27.1064
R21725 vdd.n111 vdd.n109 27.1064
R21726 vdd.n109 vdd.n104 27.1064
R21727 vdd.n104 vdd.n103 27.1064
R21728 vdd.n103 vdd.n99 27.1064
R21729 vdd.n2499 vdd.n2494 27.1064
R21730 vdd.n2556 vdd.n2499 27.1064
R21731 vdd.n2556 vdd.n2555 27.1064
R21732 vdd.n2555 vdd.n2500 27.1064
R21733 vdd.n2548 vdd.n2500 27.1064
R21734 vdd.n2548 vdd.n2547 27.1064
R21735 vdd.n2547 vdd.n2510 27.1064
R21736 vdd.n2537 vdd.n2510 27.1064
R21737 vdd.n2537 vdd.n2536 27.1064
R21738 vdd.n2536 vdd.n2517 27.1064
R21739 vdd.n2529 vdd.n2517 27.1064
R21740 vdd.n2529 vdd.n232 27.1064
R21741 vdd.n2571 vdd.n232 27.1064
R21742 vdd.n2572 vdd.n2571 27.1064
R21743 vdd.n2572 vdd.n226 27.1064
R21744 vdd.n2582 vdd.n226 27.1064
R21745 vdd.n2583 vdd.n2582 27.1064
R21746 vdd.n2583 vdd.n217 27.1064
R21747 vdd.n2589 vdd.n217 27.1064
R21748 vdd.n2590 vdd.n2589 27.1064
R21749 vdd.n2590 vdd.n208 27.1064
R21750 vdd.n2598 vdd.n208 27.1064
R21751 vdd.n2599 vdd.n2598 27.1064
R21752 vdd.n2599 vdd.n195 27.1064
R21753 vdd.n2607 vdd.n195 27.1064
R21754 vdd.n2608 vdd.n2607 27.1064
R21755 vdd.n2609 vdd.n2608 27.1064
R21756 vdd.n2609 vdd.n187 27.1064
R21757 vdd.n2617 vdd.n187 27.1064
R21758 vdd.n2618 vdd.n2617 27.1064
R21759 vdd.n2618 vdd.n178 27.1064
R21760 vdd.n2626 vdd.n178 27.1064
R21761 vdd.n2627 vdd.n2626 27.1064
R21762 vdd.n2627 vdd.n175 27.1064
R21763 vdd.n175 vdd.n174 27.1064
R21764 vdd.n174 vdd.n164 27.1064
R21765 vdd.n2639 vdd.n164 27.1064
R21766 vdd.n2640 vdd.n2639 27.1064
R21767 vdd.n2640 vdd.n153 27.1064
R21768 vdd.n2648 vdd.n153 27.1064
R21769 vdd.n2650 vdd.n148 27.1064
R21770 vdd.n2799 vdd.n148 27.1064
R21771 vdd.n2799 vdd.n2798 27.1064
R21772 vdd.n2798 vdd.n2657 27.1064
R21773 vdd.n2792 vdd.n2657 27.1064
R21774 vdd.n2792 vdd.n2791 27.1064
R21775 vdd.n2791 vdd.n2666 27.1064
R21776 vdd.n2781 vdd.n2666 27.1064
R21777 vdd.n2781 vdd.n2780 27.1064
R21778 vdd.n2780 vdd.n2673 27.1064
R21779 vdd.n2770 vdd.n2673 27.1064
R21780 vdd.n2770 vdd.n2769 27.1064
R21781 vdd.n2769 vdd.n2680 27.1064
R21782 vdd.n2687 vdd.n2680 27.1064
R21783 vdd.n2690 vdd.n2687 27.1064
R21784 vdd.n2693 vdd.n2690 27.1064
R21785 vdd.n2753 vdd.n2693 27.1064
R21786 vdd.n2753 vdd.n2752 27.1064
R21787 vdd.n2752 vdd.n2698 27.1064
R21788 vdd.n2744 vdd.n2698 27.1064
R21789 vdd.n2744 vdd.n2743 27.1064
R21790 vdd.n2743 vdd.n2706 27.1064
R21791 vdd.n2737 vdd.n2706 27.1064
R21792 vdd.n2737 vdd.n2736 27.1064
R21793 vdd.n2736 vdd.n2715 27.1064
R21794 vdd.n2726 vdd.n2715 27.1064
R21795 vdd.n2726 vdd.n132 27.1064
R21796 vdd.n2818 vdd.n132 27.1064
R21797 vdd.n2819 vdd.n2818 27.1064
R21798 vdd.n2819 vdd.n123 27.1064
R21799 vdd.n2827 vdd.n123 27.1064
R21800 vdd.n2828 vdd.n2827 27.1064
R21801 vdd.n2828 vdd.n115 27.1064
R21802 vdd.n2836 vdd.n115 27.1064
R21803 vdd.n2837 vdd.n2836 27.1064
R21804 vdd.n2837 vdd.n108 27.1064
R21805 vdd.n2847 vdd.n108 27.1064
R21806 vdd.n2849 vdd.n2847 27.1064
R21807 vdd.n2849 vdd.n2848 27.1064
R21808 vdd.n2848 vdd.n101 27.1064
R21809 vdd.n2562 vdd.n2491 27.1064
R21810 vdd.n2498 vdd.n2491 27.1064
R21811 vdd.n2504 vdd.n2498 27.1064
R21812 vdd.n2506 vdd.n2504 27.1064
R21813 vdd.n2509 vdd.n2506 27.1064
R21814 vdd.n2543 vdd.n2509 27.1064
R21815 vdd.n2543 vdd.n2542 27.1064
R21816 vdd.n2542 vdd.n2512 27.1064
R21817 vdd.n2519 vdd.n2512 27.1064
R21818 vdd.n2522 vdd.n2519 27.1064
R21819 vdd.n2528 vdd.n2522 27.1064
R21820 vdd.n2528 vdd.n236 27.1064
R21821 vdd.n2569 vdd.n236 27.1064
R21822 vdd.n2577 vdd.n228 27.1064
R21823 vdd.n2578 vdd.n2577 27.1064
R21824 vdd.n2578 vdd.n225 27.1064
R21825 vdd.n225 vdd.n224 27.1064
R21826 vdd.n224 vdd.n213 27.1064
R21827 vdd.n2592 vdd.n213 27.1064
R21828 vdd.n2593 vdd.n2592 27.1064
R21829 vdd.n2593 vdd.n204 27.1064
R21830 vdd.n2601 vdd.n204 27.1064
R21831 vdd.n2602 vdd.n2601 27.1064
R21832 vdd.n2602 vdd.n199 27.1064
R21833 vdd.n199 vdd.n198 27.1064
R21834 vdd.n198 vdd.n194 27.1064
R21835 vdd.n2615 vdd.n2614 27.1064
R21836 vdd.n2615 vdd.n180 27.1064
R21837 vdd.n2623 vdd.n180 27.1064
R21838 vdd.n2624 vdd.n2623 27.1064
R21839 vdd.n2624 vdd.n169 27.1064
R21840 vdd.n2632 vdd.n169 27.1064
R21841 vdd.n2633 vdd.n2632 27.1064
R21842 vdd.n2634 vdd.n2633 27.1064
R21843 vdd.n2634 vdd.n160 27.1064
R21844 vdd.n2642 vdd.n160 27.1064
R21845 vdd.n2643 vdd.n2642 27.1064
R21846 vdd.n2643 vdd.n157 27.1064
R21847 vdd.n157 vdd.n145 27.1064
R21848 vdd.n2804 vdd.n146 27.1064
R21849 vdd.n2660 vdd.n146 27.1064
R21850 vdd.n2662 vdd.n2660 27.1064
R21851 vdd.n2665 vdd.n2662 27.1064
R21852 vdd.n2787 vdd.n2665 27.1064
R21853 vdd.n2787 vdd.n2786 27.1064
R21854 vdd.n2786 vdd.n2668 27.1064
R21855 vdd.n2776 vdd.n2668 27.1064
R21856 vdd.n2776 vdd.n2775 27.1064
R21857 vdd.n2775 vdd.n2675 27.1064
R21858 vdd.n2682 vdd.n2675 27.1064
R21859 vdd.n2765 vdd.n2682 27.1064
R21860 vdd.n2765 vdd.n2764 27.1064
R21861 vdd.n2759 vdd.n2758 27.1064
R21862 vdd.n2758 vdd.n2691 27.1064
R21863 vdd.n2750 vdd.n2691 27.1064
R21864 vdd.n2750 vdd.n2749 27.1064
R21865 vdd.n2749 vdd.n2700 27.1064
R21866 vdd.n2709 vdd.n2700 27.1064
R21867 vdd.n2711 vdd.n2709 27.1064
R21868 vdd.n2714 vdd.n2711 27.1064
R21869 vdd.n2732 vdd.n2714 27.1064
R21870 vdd.n2732 vdd.n2731 27.1064
R21871 vdd.n2731 vdd.n2717 27.1064
R21872 vdd.n2717 vdd.n134 27.1064
R21873 vdd.n2816 vdd.n134 27.1064
R21874 vdd.n2824 vdd.n127 27.1064
R21875 vdd.n2825 vdd.n2824 27.1064
R21876 vdd.n2825 vdd.n119 27.1064
R21877 vdd.n2833 vdd.n119 27.1064
R21878 vdd.n2834 vdd.n2833 27.1064
R21879 vdd.n2834 vdd.n110 27.1064
R21880 vdd.n2842 vdd.n110 27.1064
R21881 vdd.n2843 vdd.n2842 27.1064
R21882 vdd.n2843 vdd.n106 27.1064
R21883 vdd.n106 vdd.n105 27.1064
R21884 vdd.n105 vdd.n100 27.1064
R21885 vdd.n2810 vdd.n100 27.1064
R21886 vdd.n812 vdd.n756 27.1064
R21887 vdd.n788 vdd.n756 27.1064
R21888 vdd.n801 vdd.n788 27.1064
R21889 vdd.n801 vdd.n800 27.1064
R21890 vdd.n800 vdd.n792 27.1064
R21891 vdd.n792 vdd.n791 27.1064
R21892 vdd.n791 vdd.n790 27.1064
R21893 vdd.n790 vdd.n690 27.1064
R21894 vdd.n1159 vdd.n691 27.1064
R21895 vdd.n1032 vdd.n691 27.1064
R21896 vdd.n1033 vdd.n1032 27.1064
R21897 vdd.n1049 vdd.n1033 27.1064
R21898 vdd.n1049 vdd.n1048 27.1064
R21899 vdd.n1048 vdd.n1047 27.1064
R21900 vdd.n1047 vdd.n1046 27.1064
R21901 vdd.n1046 vdd.n1045 27.1064
R21902 vdd.n1045 vdd.n1044 27.1064
R21903 vdd.n1044 vdd.n1043 27.1064
R21904 vdd.n1043 vdd.n1042 27.1064
R21905 vdd.n1042 vdd.n1041 27.1064
R21906 vdd.n1041 vdd.n1040 27.1064
R21907 vdd.n1040 vdd.n1039 27.1064
R21908 vdd.n1039 vdd.n1038 27.1064
R21909 vdd.n1038 vdd.n1037 27.1064
R21910 vdd.n1037 vdd.n1036 27.1064
R21911 vdd.n1036 vdd.n1035 27.1064
R21912 vdd.n1035 vdd.n1034 27.1064
R21913 vdd.n1034 vdd.n988 27.1064
R21914 vdd.n1111 vdd.n988 27.1064
R21915 vdd.n1115 vdd.n1114 27.1064
R21916 vdd.n1115 vdd.n601 27.1064
R21917 vdd.n1522 vdd.n601 27.1064
R21918 vdd.n1522 vdd.n1521 27.1064
R21919 vdd.n1521 vdd.n602 27.1064
R21920 vdd.n602 vdd.n592 27.1064
R21921 vdd.n1535 vdd.n592 27.1064
R21922 vdd.n1538 vdd.n1535 27.1064
R21923 vdd.n1538 vdd.n1537 27.1064
R21924 vdd.n1537 vdd.n1536 27.1064
R21925 vdd.n1536 vdd.n569 27.1064
R21926 vdd.n1560 vdd.n569 27.1064
R21927 vdd.n1569 vdd.n1560 27.1064
R21928 vdd.n1569 vdd.n1568 27.1064
R21929 vdd.n1568 vdd.n1567 27.1064
R21930 vdd.n1567 vdd.n1566 27.1064
R21931 vdd.n1566 vdd.n1565 27.1064
R21932 vdd.n1565 vdd.n1564 27.1064
R21933 vdd.n1564 vdd.n1563 27.1064
R21934 vdd.n1563 vdd.n1562 27.1064
R21935 vdd.n1562 vdd.n1561 27.1064
R21936 vdd.n1632 vdd.n1631 27.1064
R21937 vdd.n1631 vdd.n1630 27.1064
R21938 vdd.n1630 vdd.n1629 27.1064
R21939 vdd.n1629 vdd.n1628 27.1064
R21940 vdd.n1628 vdd.n1627 27.1064
R21941 vdd.n1627 vdd.n1626 27.1064
R21942 vdd.n1626 vdd.n1625 27.1064
R21943 vdd.n1625 vdd.n1624 27.1064
R21944 vdd.n1624 vdd.n1623 27.1064
R21945 vdd.n1623 vdd.n1622 27.1064
R21946 vdd.n1622 vdd.n1621 27.1064
R21947 vdd.n1621 vdd.n465 27.1064
R21948 vdd.n1721 vdd.n465 27.1064
R21949 vdd.n1721 vdd.n1720 27.1064
R21950 vdd.n1720 vdd.n466 27.1064
R21951 vdd.n1800 vdd.n449 27.1064
R21952 vdd.n1801 vdd.n1800 27.1064
R21953 vdd.n1801 vdd.n440 27.1064
R21954 vdd.n1809 vdd.n440 27.1064
R21955 vdd.n1811 vdd.n427 27.1064
R21956 vdd.n1819 vdd.n427 27.1064
R21957 vdd.n1820 vdd.n1819 27.1064
R21958 vdd.n1821 vdd.n1820 27.1064
R21959 vdd.n1821 vdd.n418 27.1064
R21960 vdd.n1829 vdd.n418 27.1064
R21961 vdd.n1830 vdd.n1829 27.1064
R21962 vdd.n1830 vdd.n409 27.1064
R21963 vdd.n1838 vdd.n409 27.1064
R21964 vdd.n1839 vdd.n1838 27.1064
R21965 vdd.n1839 vdd.n404 27.1064
R21966 vdd.n404 vdd.n403 27.1064
R21967 vdd.n403 vdd.n393 27.1064
R21968 vdd.n1851 vdd.n393 27.1064
R21969 vdd.n1852 vdd.n1851 27.1064
R21970 vdd.n1852 vdd.n384 27.1064
R21971 vdd.n1860 vdd.n384 27.1064
R21972 vdd.n1861 vdd.n1860 27.1064
R21973 vdd.n1861 vdd.n380 27.1064
R21974 vdd.n380 vdd.n375 27.1064
R21975 vdd.n375 vdd.n374 27.1064
R21976 vdd.n347 vdd.n344 27.1064
R21977 vdd.n347 vdd.n317 27.1064
R21978 vdd.n322 vdd.n317 27.1064
R21979 vdd.n324 vdd.n322 27.1064
R21980 vdd.n328 vdd.n324 27.1064
R21981 vdd.n332 vdd.n328 27.1064
R21982 vdd.n2056 vdd.n332 27.1064
R21983 vdd.n2062 vdd.n2056 27.1064
R21984 vdd.n2063 vdd.n2062 27.1064
R21985 vdd.n2063 vdd.n2046 27.1064
R21986 vdd.n2071 vdd.n2046 27.1064
R21987 vdd.n2072 vdd.n2071 27.1064
R21988 vdd.n2073 vdd.n2072 27.1064
R21989 vdd.n2073 vdd.n2039 27.1064
R21990 vdd.n2081 vdd.n2039 27.1064
R21991 vdd.n2082 vdd.n2081 27.1064
R21992 vdd.n2082 vdd.n2032 27.1064
R21993 vdd.n2090 vdd.n2032 27.1064
R21994 vdd.n2091 vdd.n2090 27.1064
R21995 vdd.n2091 vdd.n2029 27.1064
R21996 vdd.n2029 vdd.n2028 27.1064
R21997 vdd.n2103 vdd.n2019 27.1064
R21998 vdd.n2104 vdd.n2103 27.1064
R21999 vdd.n2104 vdd.n2013 27.1064
R22000 vdd.n2112 vdd.n2013 27.1064
R22001 vdd.n2113 vdd.n2112 27.1064
R22002 vdd.n2113 vdd.n2005 27.1064
R22003 vdd.n2122 vdd.n2005 27.1064
R22004 vdd.n2123 vdd.n2122 27.1064
R22005 vdd.n2124 vdd.n2123 27.1064
R22006 vdd.n2124 vdd.n1998 27.1064
R22007 vdd.n2132 vdd.n1998 27.1064
R22008 vdd.n2133 vdd.n2132 27.1064
R22009 vdd.n2133 vdd.n1992 27.1064
R22010 vdd.n2141 vdd.n1992 27.1064
R22011 vdd.n2142 vdd.n2141 27.1064
R22012 vdd.n2142 vdd.n1989 27.1064
R22013 vdd.n1989 vdd.n1988 27.1064
R22014 vdd.n1988 vdd.n1980 27.1064
R22015 vdd.n2154 vdd.n1980 27.1064
R22016 vdd.n2155 vdd.n2154 27.1064
R22017 vdd.n2155 vdd.n240 27.1064
R22018 vdd.n868 vdd.n867 27.1064
R22019 vdd.n867 vdd.n846 27.1064
R22020 vdd.n858 vdd.n846 27.1064
R22021 vdd.n858 vdd.n857 27.1064
R22022 vdd.n857 vdd.n850 27.1064
R22023 vdd.n850 vdd.n689 27.1064
R22024 vdd.n1164 vdd.n689 27.1064
R22025 vdd.n1171 vdd.n685 27.1064
R22026 vdd.n1172 vdd.n1171 27.1064
R22027 vdd.n1172 vdd.n680 27.1064
R22028 vdd.n1180 vdd.n680 27.1064
R22029 vdd.n1181 vdd.n1180 27.1064
R22030 vdd.n1181 vdd.n675 27.1064
R22031 vdd.n1190 vdd.n675 27.1064
R22032 vdd.n1191 vdd.n1190 27.1064
R22033 vdd.n1192 vdd.n1191 27.1064
R22034 vdd.n1192 vdd.n670 27.1064
R22035 vdd.n1200 vdd.n670 27.1064
R22036 vdd.n1201 vdd.n1200 27.1064
R22037 vdd.n1201 vdd.n665 27.1064
R22038 vdd.n1209 vdd.n665 27.1064
R22039 vdd.n1210 vdd.n1209 27.1064
R22040 vdd.n1210 vdd.n660 27.1064
R22041 vdd.n1219 vdd.n660 27.1064
R22042 vdd.n1220 vdd.n1219 27.1064
R22043 vdd.n1221 vdd.n1220 27.1064
R22044 vdd.n1221 vdd.n655 27.1064
R22045 vdd.n1229 vdd.n655 27.1064
R22046 vdd.n1231 vdd.n650 27.1064
R22047 vdd.n1239 vdd.n650 27.1064
R22048 vdd.n1240 vdd.n1239 27.1064
R22049 vdd.n1240 vdd.n645 27.1064
R22050 vdd.n1249 vdd.n645 27.1064
R22051 vdd.n1250 vdd.n1249 27.1064
R22052 vdd.n1251 vdd.n1250 27.1064
R22053 vdd.n1251 vdd.n640 27.1064
R22054 vdd.n1259 vdd.n640 27.1064
R22055 vdd.n1260 vdd.n1259 27.1064
R22056 vdd.n1260 vdd.n635 27.1064
R22057 vdd.n1268 vdd.n635 27.1064
R22058 vdd.n1269 vdd.n1268 27.1064
R22059 vdd.n1269 vdd.n630 27.1064
R22060 vdd.n1278 vdd.n630 27.1064
R22061 vdd.n1279 vdd.n1278 27.1064
R22062 vdd.n1280 vdd.n1279 27.1064
R22063 vdd.n1280 vdd.n625 27.1064
R22064 vdd.n1288 vdd.n625 27.1064
R22065 vdd.n1289 vdd.n1288 27.1064
R22066 vdd.n1289 vdd.n620 27.1064
R22067 vdd.n1488 vdd.n1487 27.1064
R22068 vdd.n1487 vdd.n1303 27.1064
R22069 vdd.n1308 vdd.n1303 27.1064
R22070 vdd.n1478 vdd.n1308 27.1064
R22071 vdd.n1478 vdd.n1477 27.1064
R22072 vdd.n1477 vdd.n1309 27.1064
R22073 vdd.n1469 vdd.n1309 27.1064
R22074 vdd.n1469 vdd.n1468 27.1064
R22075 vdd.n1468 vdd.n1314 27.1064
R22076 vdd.n1460 vdd.n1314 27.1064
R22077 vdd.n1460 vdd.n1459 27.1064
R22078 vdd.n1459 vdd.n1319 27.1064
R22079 vdd.n1324 vdd.n1319 27.1064
R22080 vdd.n1450 vdd.n1324 27.1064
R22081 vdd.n1450 vdd.n1449 27.1064
R22082 vdd.n1449 vdd.n1325 27.1064
R22083 vdd.n1441 vdd.n1325 27.1064
R22084 vdd.n1441 vdd.n1440 27.1064
R22085 vdd.n1440 vdd.n1330 27.1064
R22086 vdd.n1432 vdd.n1330 27.1064
R22087 vdd.n1432 vdd.n1431 27.1064
R22088 vdd.n1428 vdd.n1427 27.1064
R22089 vdd.n1427 vdd.n1337 27.1064
R22090 vdd.n1420 vdd.n1337 27.1064
R22091 vdd.n1420 vdd.n1419 27.1064
R22092 vdd.n1419 vdd.n1344 27.1064
R22093 vdd.n1412 vdd.n1344 27.1064
R22094 vdd.n1412 vdd.n1411 27.1064
R22095 vdd.n1411 vdd.n1350 27.1064
R22096 vdd.n1404 vdd.n1350 27.1064
R22097 vdd.n1404 vdd.n1403 27.1064
R22098 vdd.n1403 vdd.n1402 27.1064
R22099 vdd.n1402 vdd.n1356 27.1064
R22100 vdd.n1395 vdd.n1356 27.1064
R22101 vdd.n1395 vdd.n1394 27.1064
R22102 vdd.n1394 vdd.n1363 27.1064
R22103 vdd.n1387 vdd.n1363 27.1064
R22104 vdd.n1387 vdd.n1386 27.1064
R22105 vdd.n1386 vdd.n1369 27.1064
R22106 vdd.n1379 vdd.n1369 27.1064
R22107 vdd.n1379 vdd.n1378 27.1064
R22108 vdd.n1378 vdd.n306 27.1064
R22109 vdd.n2330 vdd.n306 27.1064
R22110 vdd.n2347 vdd.n290 27.1064
R22111 vdd.n2357 vdd.n290 27.1064
R22112 vdd.n2358 vdd.n2357 27.1064
R22113 vdd.n2359 vdd.n2358 27.1064
R22114 vdd.n2359 vdd.n286 27.1064
R22115 vdd.n2368 vdd.n286 27.1064
R22116 vdd.n2369 vdd.n2368 27.1064
R22117 vdd.n2369 vdd.n282 27.1064
R22118 vdd.n2378 vdd.n282 27.1064
R22119 vdd.n2379 vdd.n2378 27.1064
R22120 vdd.n2379 vdd.n278 27.1064
R22121 vdd.n2389 vdd.n278 27.1064
R22122 vdd.n2390 vdd.n2389 27.1064
R22123 vdd.n2391 vdd.n2390 27.1064
R22124 vdd.n2391 vdd.n274 27.1064
R22125 vdd.n2400 vdd.n274 27.1064
R22126 vdd.n2401 vdd.n2400 27.1064
R22127 vdd.n2401 vdd.n270 27.1064
R22128 vdd.n2410 vdd.n270 27.1064
R22129 vdd.n2412 vdd.n2410 27.1064
R22130 vdd.n2412 vdd.n2411 27.1064
R22131 vdd.n2423 vdd.n2422 27.1064
R22132 vdd.n2424 vdd.n2423 27.1064
R22133 vdd.n2424 vdd.n262 27.1064
R22134 vdd.n2433 vdd.n262 27.1064
R22135 vdd.n2434 vdd.n2433 27.1064
R22136 vdd.n2434 vdd.n258 27.1064
R22137 vdd.n2443 vdd.n258 27.1064
R22138 vdd.n2444 vdd.n2443 27.1064
R22139 vdd.n2444 vdd.n254 27.1064
R22140 vdd.n2454 vdd.n254 27.1064
R22141 vdd.n2455 vdd.n2454 27.1064
R22142 vdd.n2456 vdd.n2455 27.1064
R22143 vdd.n2456 vdd.n250 27.1064
R22144 vdd.n2465 vdd.n250 27.1064
R22145 vdd.n2466 vdd.n2465 27.1064
R22146 vdd.n2466 vdd.n245 27.1064
R22147 vdd.n2474 vdd.n245 27.1064
R22148 vdd.n2475 vdd.n2474 27.1064
R22149 vdd.n2475 vdd.n241 27.1064
R22150 vdd.n2481 vdd.n241 27.1064
R22151 vdd.n2329 vdd.n2328 26.3534
R22152 vdd.n2322 vdd.t175 25.9857
R22153 vdd.n1431 vdd.n1335 25.977
R22154 vdd.n2028 vdd.n2027 25.224
R22155 vdd.n2815 vdd.n127 23.7181
R22156 vdd.n2347 vdd.n2346 22.9652
R22157 vdd.n2422 vdd.n266 21.0829
R22158 vdd.n1507 vdd.n620 20.7064
R22159 vdd.n2759 vdd.n2685 20.3299
R22160 vdd.n1561 vdd.n526 20.3299
R22161 vdd.n374 vdd.n307 19.9534
R22162 vdd.n1230 vdd.n1229 18.824
R22163 vdd.n1511 vdd.t40 18.4984
R22164 vdd.n1112 vdd.n1111 18.4476
R22165 vdd.n1810 vdd.n1809 18.0711
R22166 vdd.n2569 vdd.n2568 16.9417
R22167 vdd.n2805 vdd.n2804 16.9417
R22168 vdd.n1164 vdd.n1163 16.9417
R22169 vdd.n2487 vdd.n2486 16.8187
R22170 vdd.n2488 vdd.n2487 16.8187
R22171 vdd.n142 vdd.n138 16.8187
R22172 vdd.n143 vdd.n142 16.8187
R22173 vdd.n2811 vdd.n136 16.8187
R22174 vdd.n2564 vdd.n237 16.8187
R22175 vdd.n2485 vdd.n237 16.8187
R22176 vdd.n1160 vdd.n690 16.5652
R22177 vdd.n604 vdd.n582 15.0593
R22178 vdd.n2320 vdd.n2319 15.0593
R22179 vdd.n1550 vdd.n580 15.0593
R22180 vdd.n316 vdd.n310 15.0593
R22181 vdd.n1513 vdd.n576 15.0593
R22182 vdd.n2317 vdd.n319 15.0593
R22183 vdd.n2652 vdd.n149 15.0593
R22184 vdd.n155 vdd.n152 15.0593
R22185 vdd.n2650 vdd.n2649 15.0593
R22186 vdd.n194 vdd.n189 13.5534
R22187 vdd.n2614 vdd.n189 13.5534
R22188 vdd.n2343 vdd.n296 13.2536
R22189 vdd.n605 vdd.n604 12.0476
R22190 vdd.n2320 vdd.n313 12.0476
R22191 vdd.n611 vdd.n580 12.0476
R22192 vdd.n346 vdd.n310 12.0476
R22193 vdd.n1514 vdd.n1513 12.0476
R22194 vdd.n349 vdd.n319 12.0476
R22195 vdd.n2646 vdd.n149 12.0476
R22196 vdd.n156 vdd.n155 12.0476
R22197 vdd.n2649 vdd.n2648 12.0476
R22198 vdd.n1160 vdd.n1159 10.5417
R22199 vdd.n1490 vdd.n524 10.4005
R22200 vdd.n1504 vdd.n524 10.388
R22201 vdd.n2568 vdd.n228 10.1652
R22202 vdd.n2805 vdd.n145 10.1652
R22203 vdd.n1163 vdd.n685 10.1652
R22204 vdd.n459 vdd.t251 9.52217
R22205 vdd.n459 vdd.t135 9.52217
R22206 vdd.n983 vdd.t81 9.52217
R22207 vdd.n983 vdd.t132 9.52217
R22208 vdd.n637 vdd.t178 9.52217
R22209 vdd.n637 vdd.t305 9.52217
R22210 vdd.n170 vdd.t123 9.52217
R22211 vdd.n170 vdd.t9 9.52217
R22212 vdd.n1969 vdd.t109 9.52217
R22213 vdd.n1969 vdd.t308 9.52217
R22214 vdd.n1963 vdd.t45 9.52217
R22215 vdd.n1963 vdd.t276 9.52217
R22216 vdd.n1957 vdd.t263 9.52217
R22217 vdd.n1957 vdd.t157 9.52217
R22218 vdd.n1951 vdd.t152 9.52217
R22219 vdd.n1951 vdd.t39 9.52217
R22220 vdd.n1945 vdd.t220 9.52217
R22221 vdd.n1945 vdd.t101 9.52217
R22222 vdd.n1939 vdd.t97 9.52217
R22223 vdd.n1939 vdd.t304 9.52217
R22224 vdd.n1933 vdd.t275 9.52217
R22225 vdd.n1933 vdd.t91 9.52217
R22226 vdd.n1928 vdd.t260 9.52217
R22227 vdd.n1928 vdd.t151 9.52217
R22228 vdd.n1923 vdd.t143 9.52217
R22229 vdd.n1923 vdd.t31 9.52217
R22230 vdd.n1918 vdd.t211 9.52217
R22231 vdd.n1918 vdd.t1 9.52217
R22232 vdd.n335 vdd.t295 9.52217
R22233 vdd.n335 vdd.t209 9.52217
R22234 vdd.n338 vdd.t271 9.52217
R22235 vdd.n338 vdd.t79 9.52217
R22236 vdd.n1747 vdd.t174 9.52217
R22237 vdd.n1747 vdd.t301 9.52217
R22238 vdd.n1744 vdd.t273 9.52217
R22239 vdd.n1744 vdd.t171 9.52217
R22240 vdd.n1741 vdd.t258 9.52217
R22241 vdd.n1741 vdd.t145 9.52217
R22242 vdd.n1738 vdd.t234 9.52217
R22243 vdd.n1738 vdd.t27 9.52217
R22244 vdd.n1736 vdd.t210 9.52217
R22245 vdd.n1736 vdd.t314 9.52217
R22246 vdd.n1733 vdd.t290 9.52217
R22247 vdd.n1733 vdd.t297 9.52217
R22248 vdd.n1730 vdd.t267 9.52217
R22249 vdd.n1730 vdd.t166 9.52217
R22250 vdd.n1724 vdd.t129 9.52217
R22251 vdd.n1724 vdd.t17 9.52217
R22252 vdd.n479 vdd.t67 9.52217
R22253 vdd.n479 vdd.t311 9.52217
R22254 vdd.n492 vdd.t280 9.52217
R22255 vdd.n492 vdd.t190 9.52217
R22256 vdd.n1664 vdd.t265 9.52217
R22257 vdd.n1664 vdd.t63 9.52217
R22258 vdd.n550 vdd.t93 9.52217
R22259 vdd.n550 vdd.t7 9.52217
R22260 vdd.n563 vdd.t298 9.52217
R22261 vdd.n563 vdd.t212 9.52217
R22262 vdd.n584 vdd.t272 9.52217
R22263 vdd.n584 vdd.t85 9.52217
R22264 vdd.n587 vdd.t257 9.52217
R22265 vdd.n587 vdd.t144 9.52217
R22266 vdd.n1525 vdd.t140 9.52217
R22267 vdd.n1525 vdd.t25 9.52217
R22268 vdd.n978 vdd.t287 9.52217
R22269 vdd.n978 vdd.t200 9.52217
R22270 vdd.n972 vdd.t195 9.52217
R22271 vdd.n972 vdd.t73 9.52217
R22272 vdd.n966 vdd.t250 9.52217
R22273 vdd.n966 vdd.t55 9.52217
R22274 vdd.n960 vdd.t13 9.52217
R22275 vdd.n960 vdd.t245 9.52217
R22276 vdd.n954 vdd.t309 9.52217
R22277 vdd.n954 vdd.t128 9.52217
R22278 vdd.n705 vdd.t277 9.52217
R22279 vdd.n705 vdd.t189 9.52217
R22280 vdd.n2844 vdd.t249 9.52217
R22281 vdd.n2844 vdd.t253 9.52217
R22282 vdd.n116 vdd.t286 9.52217
R22283 vdd.n116 vdd.t113 9.52217
R22284 vdd.n124 vdd.t194 9.52217
R22285 vdd.n124 vdd.t71 9.52217
R22286 vdd.n2721 vdd.t161 9.52217
R22287 vdd.n2721 vdd.t279 9.52217
R22288 vdd.n2733 vdd.t11 9.52217
R22289 vdd.n2733 vdd.t15 9.52217
R22290 vdd.n2704 vdd.t242 9.52217
R22291 vdd.n2704 vdd.t127 9.52217
R22292 vdd.n2696 vdd.t182 9.52217
R22293 vdd.n2696 vdd.t3 9.52217
R22294 vdd.n2777 vdd.t131 9.52217
R22295 vdd.n2777 vdd.t137 9.52217
R22296 vdd.n2788 vdd.t199 9.52217
R22297 vdd.n2788 vdd.t77 9.52217
R22298 vdd.n2655 vdd.t69 9.52217
R22299 vdd.n2655 vdd.t284 9.52217
R22300 vdd.n150 vdd.t5 9.52217
R22301 vdd.n150 vdd.t192 9.52217
R22302 vdd.n161 vdd.t224 9.52217
R22303 vdd.n161 vdd.t247 9.52217
R22304 vdd.n181 vdd.t184 9.52217
R22305 vdd.n181 vdd.t289 9.52217
R22306 vdd.n205 vdd.t117 9.52217
R22307 vdd.n205 vdd.t19 9.52217
R22308 vdd.n214 vdd.t75 9.52217
R22309 vdd.n214 vdd.t294 9.52217
R22310 vdd.n2579 vdd.t282 9.52217
R22311 vdd.n2579 vdd.t197 9.52217
R22312 vdd.n233 vdd.t186 9.52217
R22313 vdd.n233 vdd.t165 9.52217
R22314 vdd.n2520 vdd.t204 9.52217
R22315 vdd.n2520 vdd.t125 9.52217
R22316 vdd.n2544 vdd.t170 9.52217
R22317 vdd.n2544 vdd.t292 9.52217
R22318 vdd.n2501 vdd.t134 9.52217
R22319 vdd.n2501 vdd.t270 9.52217
R22320 vdd.n682 vdd.t206 9.52217
R22321 vdd.n682 vdd.t83 9.52217
R22322 vdd.n677 vdd.t236 9.52217
R22323 vdd.n677 vdd.t23 9.52217
R22324 vdd.n672 vdd.t256 9.52217
R22325 vdd.n672 vdd.t142 9.52217
R22326 vdd.n667 vdd.t147 9.52217
R22327 vdd.n667 vdd.t274 9.52217
R22328 vdd.n662 vdd.t89 9.52217
R22329 vdd.n662 vdd.t300 9.52217
R22330 vdd.n657 vdd.t214 9.52217
R22331 vdd.n657 vdd.t95 9.52217
R22332 vdd.n652 vdd.t302 9.52217
R22333 vdd.n652 vdd.t33 9.52217
R22334 vdd.n647 vdd.t37 9.52217
R22335 vdd.n647 vdd.t261 9.52217
R22336 vdd.n642 vdd.t154 9.52217
R22337 vdd.n642 vdd.t41 9.52217
R22338 vdd.n632 vdd.t226 9.52217
R22339 vdd.n632 vdd.t107 9.52217
R22340 vdd.n627 vdd.t306 9.52217
R22341 vdd.n627 vdd.t244 9.52217
R22342 vdd.n1305 vdd.t168 9.52217
R22343 vdd.n1305 vdd.t296 9.52217
R22344 vdd.n1311 vdd.t208 9.52217
R22345 vdd.n1311 vdd.t87 9.52217
R22346 vdd.n1316 vdd.t299 9.52217
R22347 vdd.n1316 vdd.t238 9.52217
R22348 vdd.n1321 vdd.t29 9.52217
R22349 vdd.n1321 vdd.t259 9.52217
R22350 vdd.n1327 vdd.t150 9.52217
R22351 vdd.n1327 vdd.t35 9.52217
R22352 vdd.n1332 vdd.t173 9.52217
R22353 vdd.n1332 vdd.t59 9.52217
R22354 vdd.n1339 vdd.t216 9.52217
R22355 vdd.n1339 vdd.t222 9.52217
R22356 vdd.n1346 vdd.t103 9.52217
R22357 vdd.n1346 vdd.t240 9.52217
R22358 vdd.n1352 vdd.t121 9.52217
R22359 vdd.n1352 vdd.t262 9.52217
R22360 vdd.n1359 vdd.t156 9.52217
R22361 vdd.n1359 vdd.t47 9.52217
R22362 vdd.n1365 vdd.t180 9.52217
R22363 vdd.n1365 vdd.t61 9.52217
R22364 vdd.n1371 vdd.t65 9.52217
R22365 vdd.n1371 vdd.t229 9.52217
R22366 vdd.n2351 vdd.t176 9.52217
R22367 vdd.n2351 vdd.t303 9.52217
R22368 vdd.n2363 vdd.t219 9.52217
R22369 vdd.n2363 vdd.t99 9.52217
R22370 vdd.n2373 vdd.t105 9.52217
R22371 vdd.n2373 vdd.t243 9.52217
R22372 vdd.n2383 vdd.t43 9.52217
R22373 vdd.n2383 vdd.t264 9.52217
R22374 vdd.n2395 vdd.t159 9.52217
R22375 vdd.n2395 vdd.t49 9.52217
R22376 vdd.n2405 vdd.t188 9.52217
R22377 vdd.n2405 vdd.t307 9.52217
R22378 vdd.n2416 vdd.t310 9.52217
R22379 vdd.n2416 vdd.t231 9.52217
R22380 vdd.n2428 vdd.t115 9.52217
R22381 vdd.n2428 vdd.t312 9.52217
R22382 vdd.n2438 vdd.t53 9.52217
R22383 vdd.n2438 vdd.t266 9.52217
R22384 vdd.n2448 vdd.t163 9.52217
R22385 vdd.n2448 vdd.t57 9.52217
R22386 vdd.n2460 vdd.t268 9.52217
R22387 vdd.n2460 vdd.t202 9.52217
R22388 vdd.n247 vdd.t313 9.52217
R22389 vdd.n247 vdd.t233 9.52217
R22390 vdd.n2481 vdd.n2480 9.31222
R22391 vdd.n943 vdd.n942 9.3005
R22392 vdd.n1157 vdd.n695 9.3005
R22393 vdd.n1154 vdd.n1153 9.3005
R22394 vdd.n1152 vdd.n1151 9.3005
R22395 vdd.n1052 vdd.n700 9.3005
R22396 vdd.n1056 vdd.n1055 9.3005
R22397 vdd.n1058 vdd.n1057 9.3005
R22398 vdd.n1061 vdd.n1026 9.3005
R22399 vdd.n1065 vdd.n1064 9.3005
R22400 vdd.n1067 vdd.n1066 9.3005
R22401 vdd.n1070 vdd.n1020 9.3005
R22402 vdd.n1074 vdd.n1073 9.3005
R22403 vdd.n1076 vdd.n1075 9.3005
R22404 vdd.n1079 vdd.n1014 9.3005
R22405 vdd.n1083 vdd.n1082 9.3005
R22406 vdd.n1085 vdd.n1084 9.3005
R22407 vdd.n1088 vdd.n1008 9.3005
R22408 vdd.n1092 vdd.n1091 9.3005
R22409 vdd.n1094 vdd.n1093 9.3005
R22410 vdd.n1097 vdd.n1002 9.3005
R22411 vdd.n1101 vdd.n1100 9.3005
R22412 vdd.n1103 vdd.n1102 9.3005
R22413 vdd.n1109 vdd.n998 9.3005
R22414 vdd.n997 vdd.n984 9.3005
R22415 vdd.n996 vdd.n987 9.3005
R22416 vdd.n995 vdd.n599 9.3005
R22417 vdd.n994 vdd.n600 9.3005
R22418 vdd.n1519 vdd.n615 9.3005
R22419 vdd.n614 vdd.n596 9.3005
R22420 vdd.n613 vdd.n593 9.3005
R22421 vdd.n612 vdd.n589 9.3005
R22422 vdd.n611 vdd.n591 9.3005
R22423 vdd.n1550 vdd.n1549 9.3005
R22424 vdd.n1552 vdd.n1551 9.3005
R22425 vdd.n1557 vdd.n575 9.3005
R22426 vdd.n574 vdd.n567 9.3005
R22427 vdd.n568 vdd.n560 9.3005
R22428 vdd.n1578 vdd.n1577 9.3005
R22429 vdd.n1580 vdd.n1579 9.3005
R22430 vdd.n1583 vdd.n547 9.3005
R22431 vdd.n1591 vdd.n1590 9.3005
R22432 vdd.n1593 vdd.n1592 9.3005
R22433 vdd.n1596 vdd.n534 9.3005
R22434 vdd.n1649 vdd.n1648 9.3005
R22435 vdd.n1651 vdd.n1650 9.3005
R22436 vdd.n1655 vdd.n530 9.3005
R22437 vdd.n943 vdd.n710 9.3005
R22438 vdd.n1157 vdd.n693 9.3005
R22439 vdd.n1154 vdd.n698 9.3005
R22440 vdd.n1151 vdd.n702 9.3005
R22441 vdd.n1053 vdd.n1052 9.3005
R22442 vdd.n1055 vdd.n1054 9.3005
R22443 vdd.n1058 vdd.n1028 9.3005
R22444 vdd.n1062 vdd.n1061 9.3005
R22445 vdd.n1064 vdd.n1063 9.3005
R22446 vdd.n1067 vdd.n1022 9.3005
R22447 vdd.n1071 vdd.n1070 9.3005
R22448 vdd.n1073 vdd.n1072 9.3005
R22449 vdd.n1076 vdd.n1016 9.3005
R22450 vdd.n1080 vdd.n1079 9.3005
R22451 vdd.n1082 vdd.n1081 9.3005
R22452 vdd.n1085 vdd.n1010 9.3005
R22453 vdd.n1089 vdd.n1088 9.3005
R22454 vdd.n1091 vdd.n1090 9.3005
R22455 vdd.n1094 vdd.n1004 9.3005
R22456 vdd.n1098 vdd.n1097 9.3005
R22457 vdd.n1100 vdd.n1099 9.3005
R22458 vdd.n1103 vdd.n1001 9.3005
R22459 vdd.n1109 vdd.n993 9.3005
R22460 vdd.n992 vdd.n984 9.3005
R22461 vdd.n991 vdd.n987 9.3005
R22462 vdd.n990 vdd.n599 9.3005
R22463 vdd.n989 vdd.n600 9.3005
R22464 vdd.n1519 vdd.n609 9.3005
R22465 vdd.n608 vdd.n596 9.3005
R22466 vdd.n607 vdd.n593 9.3005
R22467 vdd.n606 vdd.n589 9.3005
R22468 vdd.n605 vdd.n591 9.3005
R22469 vdd.n1549 vdd.n582 9.3005
R22470 vdd.n1552 vdd.n578 9.3005
R22471 vdd.n1557 vdd.n573 9.3005
R22472 vdd.n572 vdd.n567 9.3005
R22473 vdd.n571 vdd.n568 9.3005
R22474 vdd.n1577 vdd.n562 9.3005
R22475 vdd.n1580 vdd.n558 9.3005
R22476 vdd.n1583 vdd.n555 9.3005
R22477 vdd.n1590 vdd.n549 9.3005
R22478 vdd.n1593 vdd.n545 9.3005
R22479 vdd.n1596 vdd.n542 9.3005
R22480 vdd.n1648 vdd.n536 9.3005
R22481 vdd.n1651 vdd.n533 9.3005
R22482 vdd.n1655 vdd.n528 9.3005
R22483 vdd.n810 vdd.n760 9.3005
R22484 vdd.n807 vdd.n806 9.3005
R22485 vdd.n805 vdd.n804 9.3005
R22486 vdd.n787 vdd.n783 9.3005
R22487 vdd.n798 vdd.n797 9.3005
R22488 vdd.n935 vdd.n711 9.3005
R22489 vdd.n940 vdd.n939 9.3005
R22490 vdd.n941 vdd.n709 9.3005
R22491 vdd.n810 vdd.n758 9.3005
R22492 vdd.n807 vdd.n764 9.3005
R22493 vdd.n804 vdd.n785 9.3005
R22494 vdd.n794 vdd.n787 9.3005
R22495 vdd.n798 vdd.n795 9.3005
R22496 vdd.n935 vdd.n718 9.3005
R22497 vdd.n939 vdd.n714 9.3005
R22498 vdd.n713 vdd.n709 9.3005
R22499 vdd.n810 vdd.n809 9.3005
R22500 vdd.n808 vdd.n807 9.3005
R22501 vdd.n804 vdd.n763 9.3005
R22502 vdd.n787 vdd.n786 9.3005
R22503 vdd.n798 vdd.n716 9.3005
R22504 vdd.n936 vdd.n935 9.3005
R22505 vdd.n939 vdd.n938 9.3005
R22506 vdd.n937 vdd.n709 9.3005
R22507 vdd.n943 vdd.n696 9.3005
R22508 vdd.n1157 vdd.n1156 9.3005
R22509 vdd.n1155 vdd.n1154 9.3005
R22510 vdd.n1151 vdd.n697 9.3005
R22511 vdd.n1052 vdd.n1051 9.3005
R22512 vdd.n1055 vdd.n1030 9.3005
R22513 vdd.n1059 vdd.n1058 9.3005
R22514 vdd.n1061 vdd.n1060 9.3005
R22515 vdd.n1064 vdd.n1024 9.3005
R22516 vdd.n1068 vdd.n1067 9.3005
R22517 vdd.n1070 vdd.n1069 9.3005
R22518 vdd.n1073 vdd.n1018 9.3005
R22519 vdd.n1077 vdd.n1076 9.3005
R22520 vdd.n1079 vdd.n1078 9.3005
R22521 vdd.n1082 vdd.n1012 9.3005
R22522 vdd.n1086 vdd.n1085 9.3005
R22523 vdd.n1088 vdd.n1087 9.3005
R22524 vdd.n1091 vdd.n1006 9.3005
R22525 vdd.n1095 vdd.n1094 9.3005
R22526 vdd.n1097 vdd.n1096 9.3005
R22527 vdd.n1100 vdd.n999 9.3005
R22528 vdd.n1104 vdd.n1103 9.3005
R22529 vdd.n1109 vdd.n1108 9.3005
R22530 vdd.n1107 vdd.n984 9.3005
R22531 vdd.n1106 vdd.n987 9.3005
R22532 vdd.n1105 vdd.n599 9.3005
R22533 vdd.n616 vdd.n600 9.3005
R22534 vdd.n1519 vdd.n1518 9.3005
R22535 vdd.n1517 vdd.n596 9.3005
R22536 vdd.n1516 vdd.n593 9.3005
R22537 vdd.n1515 vdd.n589 9.3005
R22538 vdd.n1514 vdd.n591 9.3005
R22539 vdd.n1549 vdd.n576 9.3005
R22540 vdd.n1553 vdd.n1552 9.3005
R22541 vdd.n1557 vdd.n1556 9.3005
R22542 vdd.n1555 vdd.n567 9.3005
R22543 vdd.n1554 vdd.n568 9.3005
R22544 vdd.n1577 vdd.n556 9.3005
R22545 vdd.n1581 vdd.n1580 9.3005
R22546 vdd.n1583 vdd.n1582 9.3005
R22547 vdd.n1590 vdd.n543 9.3005
R22548 vdd.n1594 vdd.n1593 9.3005
R22549 vdd.n1596 vdd.n1595 9.3005
R22550 vdd.n1648 vdd.n531 9.3005
R22551 vdd.n1652 vdd.n1651 9.3005
R22552 vdd.n1655 vdd.n1654 9.3005
R22553 vdd.n812 vdd.n811 9.3005
R22554 vdd.n759 vdd.n756 9.3005
R22555 vdd.n788 vdd.n784 9.3005
R22556 vdd.n802 vdd.n801 9.3005
R22557 vdd.n800 vdd.n799 9.3005
R22558 vdd.n792 vdd.n717 9.3005
R22559 vdd.n791 vdd.n712 9.3005
R22560 vdd.n790 vdd.n789 9.3005
R22561 vdd.n944 vdd.n690 9.3005
R22562 vdd.n1159 vdd.n1158 9.3005
R22563 vdd.n694 vdd.n691 9.3005
R22564 vdd.n1032 vdd.n701 9.3005
R22565 vdd.n1033 vdd.n703 9.3005
R22566 vdd.n1050 vdd.n1049 9.3005
R22567 vdd.n1048 vdd.n1031 9.3005
R22568 vdd.n1047 vdd.n1029 9.3005
R22569 vdd.n1046 vdd.n1027 9.3005
R22570 vdd.n1045 vdd.n1025 9.3005
R22571 vdd.n1044 vdd.n1023 9.3005
R22572 vdd.n1043 vdd.n1021 9.3005
R22573 vdd.n1042 vdd.n1019 9.3005
R22574 vdd.n1041 vdd.n1017 9.3005
R22575 vdd.n1040 vdd.n1015 9.3005
R22576 vdd.n1039 vdd.n1013 9.3005
R22577 vdd.n1038 vdd.n1011 9.3005
R22578 vdd.n1037 vdd.n1009 9.3005
R22579 vdd.n1036 vdd.n1007 9.3005
R22580 vdd.n1035 vdd.n1005 9.3005
R22581 vdd.n1034 vdd.n1003 9.3005
R22582 vdd.n1000 vdd.n988 9.3005
R22583 vdd.n1111 vdd.n1110 9.3005
R22584 vdd.n1114 vdd.n1113 9.3005
R22585 vdd.n1116 vdd.n1115 9.3005
R22586 vdd.n985 vdd.n601 9.3005
R22587 vdd.n1523 vdd.n1522 9.3005
R22588 vdd.n1521 vdd.n1520 9.3005
R22589 vdd.n610 vdd.n602 9.3005
R22590 vdd.n595 vdd.n592 9.3005
R22591 vdd.n1535 vdd.n1534 9.3005
R22592 vdd.n1539 vdd.n1538 9.3005
R22593 vdd.n1537 vdd.n581 9.3005
R22594 vdd.n1536 vdd.n577 9.3005
R22595 vdd.n570 vdd.n569 9.3005
R22596 vdd.n1560 vdd.n1559 9.3005
R22597 vdd.n1570 vdd.n1569 9.3005
R22598 vdd.n1568 vdd.n561 9.3005
R22599 vdd.n1567 vdd.n557 9.3005
R22600 vdd.n1566 vdd.n554 9.3005
R22601 vdd.n1565 vdd.n548 9.3005
R22602 vdd.n1564 vdd.n544 9.3005
R22603 vdd.n1563 vdd.n541 9.3005
R22604 vdd.n1562 vdd.n535 9.3005
R22605 vdd.n1561 vdd.n532 9.3005
R22606 vdd.n1657 vdd.n1656 9.3005
R22607 vdd.n1171 vdd.n1170 9.3005
R22608 vdd.n1173 vdd.n1172 9.3005
R22609 vdd.n681 vdd.n680 9.3005
R22610 vdd.n1180 vdd.n1179 9.3005
R22611 vdd.n1182 vdd.n1181 9.3005
R22612 vdd.n676 vdd.n675 9.3005
R22613 vdd.n1190 vdd.n1189 9.3005
R22614 vdd.n1191 vdd.n674 9.3005
R22615 vdd.n1193 vdd.n1192 9.3005
R22616 vdd.n671 vdd.n670 9.3005
R22617 vdd.n1200 vdd.n1199 9.3005
R22618 vdd.n1202 vdd.n1201 9.3005
R22619 vdd.n666 vdd.n665 9.3005
R22620 vdd.n1209 vdd.n1208 9.3005
R22621 vdd.n1211 vdd.n1210 9.3005
R22622 vdd.n661 vdd.n660 9.3005
R22623 vdd.n1219 vdd.n1218 9.3005
R22624 vdd.n1220 vdd.n659 9.3005
R22625 vdd.n1222 vdd.n1221 9.3005
R22626 vdd.n656 vdd.n655 9.3005
R22627 vdd.n1229 vdd.n1228 9.3005
R22628 vdd.n1232 vdd.n1231 9.3005
R22629 vdd.n651 vdd.n650 9.3005
R22630 vdd.n1239 vdd.n1238 9.3005
R22631 vdd.n1241 vdd.n1240 9.3005
R22632 vdd.n646 vdd.n645 9.3005
R22633 vdd.n1249 vdd.n1248 9.3005
R22634 vdd.n1250 vdd.n644 9.3005
R22635 vdd.n1252 vdd.n1251 9.3005
R22636 vdd.n641 vdd.n640 9.3005
R22637 vdd.n1259 vdd.n1258 9.3005
R22638 vdd.n1261 vdd.n1260 9.3005
R22639 vdd.n636 vdd.n635 9.3005
R22640 vdd.n1268 vdd.n1267 9.3005
R22641 vdd.n1270 vdd.n1269 9.3005
R22642 vdd.n1271 vdd.n630 9.3005
R22643 vdd.n1278 vdd.n1277 9.3005
R22644 vdd.n1279 vdd.n629 9.3005
R22645 vdd.n1281 vdd.n1280 9.3005
R22646 vdd.n626 vdd.n625 9.3005
R22647 vdd.n1288 vdd.n1287 9.3005
R22648 vdd.n1290 vdd.n1289 9.3005
R22649 vdd.n686 vdd.n685 9.3005
R22650 vdd.n869 vdd.n868 9.3005
R22651 vdd.n867 vdd.n866 9.3005
R22652 vdd.n847 vdd.n846 9.3005
R22653 vdd.n859 vdd.n858 9.3005
R22654 vdd.n857 vdd.n856 9.3005
R22655 vdd.n852 vdd.n850 9.3005
R22656 vdd.n689 vdd.n688 9.3005
R22657 vdd.n1165 vdd.n1164 9.3005
R22658 vdd.n1291 vdd.n620 9.3005
R22659 vdd.n1506 vdd.n1505 9.3005
R22660 vdd.n1485 vdd.n1303 9.3005
R22661 vdd.n1308 vdd.n1304 9.3005
R22662 vdd.n1479 vdd.n1478 9.3005
R22663 vdd.n1477 vdd.n1476 9.3005
R22664 vdd.n1310 vdd.n1309 9.3005
R22665 vdd.n1470 vdd.n1469 9.3005
R22666 vdd.n1468 vdd.n1467 9.3005
R22667 vdd.n1315 vdd.n1314 9.3005
R22668 vdd.n1461 vdd.n1460 9.3005
R22669 vdd.n1459 vdd.n1458 9.3005
R22670 vdd.n1457 vdd.n1319 9.3005
R22671 vdd.n1324 vdd.n1320 9.3005
R22672 vdd.n1451 vdd.n1450 9.3005
R22673 vdd.n1449 vdd.n1448 9.3005
R22674 vdd.n1326 vdd.n1325 9.3005
R22675 vdd.n1442 vdd.n1441 9.3005
R22676 vdd.n1440 vdd.n1439 9.3005
R22677 vdd.n1331 vdd.n1330 9.3005
R22678 vdd.n1433 vdd.n1432 9.3005
R22679 vdd.n1431 vdd.n1430 9.3005
R22680 vdd.n1429 vdd.n1428 9.3005
R22681 vdd.n1427 vdd.n1426 9.3005
R22682 vdd.n1338 vdd.n1337 9.3005
R22683 vdd.n1421 vdd.n1420 9.3005
R22684 vdd.n1419 vdd.n1418 9.3005
R22685 vdd.n1345 vdd.n1344 9.3005
R22686 vdd.n1413 vdd.n1412 9.3005
R22687 vdd.n1411 vdd.n1410 9.3005
R22688 vdd.n1351 vdd.n1350 9.3005
R22689 vdd.n1405 vdd.n1404 9.3005
R22690 vdd.n1403 vdd.n1355 9.3005
R22691 vdd.n1402 vdd.n1401 9.3005
R22692 vdd.n1358 vdd.n1356 9.3005
R22693 vdd.n1396 vdd.n1395 9.3005
R22694 vdd.n1394 vdd.n1393 9.3005
R22695 vdd.n1364 vdd.n1363 9.3005
R22696 vdd.n1388 vdd.n1387 9.3005
R22697 vdd.n1386 vdd.n1385 9.3005
R22698 vdd.n1370 vdd.n1369 9.3005
R22699 vdd.n1380 vdd.n1379 9.3005
R22700 vdd.n1378 vdd.n1377 9.3005
R22701 vdd.n1487 vdd.n1486 9.3005
R22702 vdd.n1489 vdd.n1488 9.3005
R22703 vdd.n2328 vdd.n296 9.3005
R22704 vdd.n2331 vdd.n2330 9.3005
R22705 vdd.n1375 vdd.n306 9.3005
R22706 vdd.n1633 vdd.n1632 9.3005
R22707 vdd.n1631 vdd.n510 9.3005
R22708 vdd.n1630 vdd.n507 9.3005
R22709 vdd.n1629 vdd.n504 9.3005
R22710 vdd.n1628 vdd.n502 9.3005
R22711 vdd.n1627 vdd.n499 9.3005
R22712 vdd.n1626 vdd.n496 9.3005
R22713 vdd.n1625 vdd.n490 9.3005
R22714 vdd.n1624 vdd.n486 9.3005
R22715 vdd.n1623 vdd.n483 9.3005
R22716 vdd.n1622 vdd.n477 9.3005
R22717 vdd.n1621 vdd.n470 9.3005
R22718 vdd.n474 vdd.n465 9.3005
R22719 vdd.n1722 vdd.n1721 9.3005
R22720 vdd.n1720 vdd.n1719 9.3005
R22721 vdd.n466 vdd.n456 9.3005
R22722 vdd.n1637 vdd.n509 9.3005
R22723 vdd.n1673 vdd.n1672 9.3005
R22724 vdd.n1675 vdd.n1674 9.3005
R22725 vdd.n1678 vdd.n501 9.3005
R22726 vdd.n1683 vdd.n1682 9.3005
R22727 vdd.n1685 vdd.n1684 9.3005
R22728 vdd.n1688 vdd.n489 9.3005
R22729 vdd.n1696 vdd.n1695 9.3005
R22730 vdd.n1698 vdd.n1697 9.3005
R22731 vdd.n1701 vdd.n476 9.3005
R22732 vdd.n1709 vdd.n1708 9.3005
R22733 vdd.n1713 vdd.n1712 9.3005
R22734 vdd.n1711 vdd.n463 9.3005
R22735 vdd.n1710 vdd.n464 9.3005
R22736 vdd.n1718 vdd.n455 9.3005
R22737 vdd.n1637 vdd.n1635 9.3005
R22738 vdd.n1672 vdd.n511 9.3005
R22739 vdd.n1675 vdd.n503 9.3005
R22740 vdd.n1679 vdd.n1678 9.3005
R22741 vdd.n1682 vdd.n1680 9.3005
R22742 vdd.n1685 vdd.n500 9.3005
R22743 vdd.n1688 vdd.n497 9.3005
R22744 vdd.n1695 vdd.n491 9.3005
R22745 vdd.n1698 vdd.n487 9.3005
R22746 vdd.n1701 vdd.n484 9.3005
R22747 vdd.n1708 vdd.n478 9.3005
R22748 vdd.n1713 vdd.n473 9.3005
R22749 vdd.n472 vdd.n463 9.3005
R22750 vdd.n471 vdd.n464 9.3005
R22751 vdd.n1718 vdd.n468 9.3005
R22752 vdd.n1638 vdd.n1637 9.3005
R22753 vdd.n1672 vdd.n506 9.3005
R22754 vdd.n1676 vdd.n1675 9.3005
R22755 vdd.n1678 vdd.n1677 9.3005
R22756 vdd.n1682 vdd.n498 9.3005
R22757 vdd.n1686 vdd.n1685 9.3005
R22758 vdd.n1688 vdd.n1687 9.3005
R22759 vdd.n1695 vdd.n485 9.3005
R22760 vdd.n1699 vdd.n1698 9.3005
R22761 vdd.n1701 vdd.n1700 9.3005
R22762 vdd.n1708 vdd.n469 9.3005
R22763 vdd.n1714 vdd.n1713 9.3005
R22764 vdd.n1715 vdd.n463 9.3005
R22765 vdd.n1716 vdd.n464 9.3005
R22766 vdd.n1718 vdd.n1717 9.3005
R22767 vdd.n1794 vdd.n1793 9.3005
R22768 vdd.n1793 vdd.n457 9.3005
R22769 vdd.n1793 vdd.n452 9.3005
R22770 vdd.n2562 vdd.n2561 9.3005
R22771 vdd.n2493 vdd.n2491 9.3005
R22772 vdd.n2557 vdd.n2498 9.3005
R22773 vdd.n2554 vdd.n2504 9.3005
R22774 vdd.n2552 vdd.n2506 9.3005
R22775 vdd.n2549 vdd.n2509 9.3005
R22776 vdd.n2546 vdd.n2543 9.3005
R22777 vdd.n2542 vdd.n2541 9.3005
R22778 vdd.n2538 vdd.n2512 9.3005
R22779 vdd.n2535 vdd.n2519 9.3005
R22780 vdd.n2533 vdd.n2522 9.3005
R22781 vdd.n2530 vdd.n2528 9.3005
R22782 vdd.n2525 vdd.n236 9.3005
R22783 vdd.n2570 vdd.n2569 9.3005
R22784 vdd.n2573 vdd.n228 9.3005
R22785 vdd.n2577 vdd.n2576 9.3005
R22786 vdd.n2581 vdd.n2578 9.3005
R22787 vdd.n2584 vdd.n225 9.3005
R22788 vdd.n224 vdd.n218 9.3005
R22789 vdd.n2588 vdd.n213 9.3005
R22790 vdd.n2592 vdd.n2591 9.3005
R22791 vdd.n2594 vdd.n2593 9.3005
R22792 vdd.n2597 vdd.n204 9.3005
R22793 vdd.n2601 vdd.n2600 9.3005
R22794 vdd.n2603 vdd.n2602 9.3005
R22795 vdd.n2606 vdd.n199 9.3005
R22796 vdd.n198 vdd.n192 9.3005
R22797 vdd.n2610 vdd.n194 9.3005
R22798 vdd.n2614 vdd.n2613 9.3005
R22799 vdd.n2616 vdd.n2615 9.3005
R22800 vdd.n2619 vdd.n180 9.3005
R22801 vdd.n2623 vdd.n2622 9.3005
R22802 vdd.n2625 vdd.n2624 9.3005
R22803 vdd.n2628 vdd.n169 9.3005
R22804 vdd.n2632 vdd.n2631 9.3005
R22805 vdd.n2633 vdd.n167 9.3005
R22806 vdd.n2635 vdd.n2634 9.3005
R22807 vdd.n2638 vdd.n160 9.3005
R22808 vdd.n2642 vdd.n2641 9.3005
R22809 vdd.n2644 vdd.n2643 9.3005
R22810 vdd.n2647 vdd.n157 9.3005
R22811 vdd.n2651 vdd.n145 9.3005
R22812 vdd.n2804 vdd.n2803 9.3005
R22813 vdd.n2800 vdd.n146 9.3005
R22814 vdd.n2797 vdd.n2660 9.3005
R22815 vdd.n2796 vdd.n2662 9.3005
R22816 vdd.n2793 vdd.n2665 9.3005
R22817 vdd.n2790 vdd.n2787 9.3005
R22818 vdd.n2786 vdd.n2785 9.3005
R22819 vdd.n2782 vdd.n2668 9.3005
R22820 vdd.n2779 vdd.n2776 9.3005
R22821 vdd.n2775 vdd.n2774 9.3005
R22822 vdd.n2771 vdd.n2675 9.3005
R22823 vdd.n2768 vdd.n2682 9.3005
R22824 vdd.n2758 vdd.n2757 9.3005
R22825 vdd.n2754 vdd.n2691 9.3005
R22826 vdd.n2751 vdd.n2750 9.3005
R22827 vdd.n2749 vdd.n2748 9.3005
R22828 vdd.n2745 vdd.n2700 9.3005
R22829 vdd.n2742 vdd.n2709 9.3005
R22830 vdd.n2741 vdd.n2711 9.3005
R22831 vdd.n2738 vdd.n2714 9.3005
R22832 vdd.n2735 vdd.n2732 9.3005
R22833 vdd.n2731 vdd.n2730 9.3005
R22834 vdd.n2727 vdd.n2717 9.3005
R22835 vdd.n2723 vdd.n134 9.3005
R22836 vdd.n2817 vdd.n2816 9.3005
R22837 vdd.n2820 vdd.n127 9.3005
R22838 vdd.n2824 vdd.n2823 9.3005
R22839 vdd.n2826 vdd.n2825 9.3005
R22840 vdd.n2829 vdd.n119 9.3005
R22841 vdd.n2833 vdd.n2832 9.3005
R22842 vdd.n2835 vdd.n2834 9.3005
R22843 vdd.n2838 vdd.n110 9.3005
R22844 vdd.n2842 vdd.n2841 9.3005
R22845 vdd.n2846 vdd.n2843 9.3005
R22846 vdd.n2850 vdd.n106 9.3005
R22847 vdd.n105 vdd.n98 9.3005
R22848 vdd.n2854 vdd.n100 9.3005
R22849 vdd.n2561 vdd.n2494 9.3005
R22850 vdd.n2499 vdd.n2493 9.3005
R22851 vdd.n2557 vdd.n2556 9.3005
R22852 vdd.n2555 vdd.n2554 9.3005
R22853 vdd.n2552 vdd.n2500 9.3005
R22854 vdd.n2549 vdd.n2548 9.3005
R22855 vdd.n2547 vdd.n2546 9.3005
R22856 vdd.n2541 vdd.n2510 9.3005
R22857 vdd.n2538 vdd.n2537 9.3005
R22858 vdd.n2536 vdd.n2535 9.3005
R22859 vdd.n2533 vdd.n2517 9.3005
R22860 vdd.n2530 vdd.n2529 9.3005
R22861 vdd.n2525 vdd.n232 9.3005
R22862 vdd.n2571 vdd.n2570 9.3005
R22863 vdd.n2573 vdd.n2572 9.3005
R22864 vdd.n2576 vdd.n226 9.3005
R22865 vdd.n2582 vdd.n2581 9.3005
R22866 vdd.n2584 vdd.n2583 9.3005
R22867 vdd.n218 vdd.n217 9.3005
R22868 vdd.n2589 vdd.n2588 9.3005
R22869 vdd.n2591 vdd.n2590 9.3005
R22870 vdd.n2594 vdd.n208 9.3005
R22871 vdd.n2598 vdd.n2597 9.3005
R22872 vdd.n2600 vdd.n2599 9.3005
R22873 vdd.n2603 vdd.n195 9.3005
R22874 vdd.n2607 vdd.n2606 9.3005
R22875 vdd.n2608 vdd.n192 9.3005
R22876 vdd.n2610 vdd.n2609 9.3005
R22877 vdd.n2613 vdd.n187 9.3005
R22878 vdd.n2617 vdd.n2616 9.3005
R22879 vdd.n2619 vdd.n2618 9.3005
R22880 vdd.n2622 vdd.n178 9.3005
R22881 vdd.n2626 vdd.n2625 9.3005
R22882 vdd.n2628 vdd.n2627 9.3005
R22883 vdd.n2631 vdd.n175 9.3005
R22884 vdd.n174 vdd.n167 9.3005
R22885 vdd.n2635 vdd.n164 9.3005
R22886 vdd.n2639 vdd.n2638 9.3005
R22887 vdd.n2641 vdd.n2640 9.3005
R22888 vdd.n2644 vdd.n153 9.3005
R22889 vdd.n2648 vdd.n2647 9.3005
R22890 vdd.n2651 vdd.n2650 9.3005
R22891 vdd.n2803 vdd.n148 9.3005
R22892 vdd.n2800 vdd.n2799 9.3005
R22893 vdd.n2798 vdd.n2797 9.3005
R22894 vdd.n2796 vdd.n2657 9.3005
R22895 vdd.n2793 vdd.n2792 9.3005
R22896 vdd.n2791 vdd.n2790 9.3005
R22897 vdd.n2785 vdd.n2666 9.3005
R22898 vdd.n2782 vdd.n2781 9.3005
R22899 vdd.n2780 vdd.n2779 9.3005
R22900 vdd.n2774 vdd.n2673 9.3005
R22901 vdd.n2771 vdd.n2770 9.3005
R22902 vdd.n2769 vdd.n2768 9.3005
R22903 vdd.n2766 vdd.n2680 9.3005
R22904 vdd.n2763 vdd.n2687 9.3005
R22905 vdd.n2760 vdd.n2690 9.3005
R22906 vdd.n2757 vdd.n2693 9.3005
R22907 vdd.n2754 vdd.n2753 9.3005
R22908 vdd.n2752 vdd.n2751 9.3005
R22909 vdd.n2748 vdd.n2698 9.3005
R22910 vdd.n2745 vdd.n2744 9.3005
R22911 vdd.n2743 vdd.n2742 9.3005
R22912 vdd.n2741 vdd.n2706 9.3005
R22913 vdd.n2738 vdd.n2737 9.3005
R22914 vdd.n2736 vdd.n2735 9.3005
R22915 vdd.n2730 vdd.n2715 9.3005
R22916 vdd.n2727 vdd.n2726 9.3005
R22917 vdd.n2723 vdd.n132 9.3005
R22918 vdd.n2818 vdd.n2817 9.3005
R22919 vdd.n2820 vdd.n2819 9.3005
R22920 vdd.n2823 vdd.n123 9.3005
R22921 vdd.n2827 vdd.n2826 9.3005
R22922 vdd.n2829 vdd.n2828 9.3005
R22923 vdd.n2832 vdd.n115 9.3005
R22924 vdd.n2836 vdd.n2835 9.3005
R22925 vdd.n2838 vdd.n2837 9.3005
R22926 vdd.n2841 vdd.n108 9.3005
R22927 vdd.n2847 vdd.n2846 9.3005
R22928 vdd.n2850 vdd.n2849 9.3005
R22929 vdd.n2848 vdd.n98 9.3005
R22930 vdd.n2854 vdd.n101 9.3005
R22931 vdd.n2561 vdd.n2492 9.3005
R22932 vdd.n2496 vdd.n2493 9.3005
R22933 vdd.n2557 vdd.n2497 9.3005
R22934 vdd.n2554 vdd.n2503 9.3005
R22935 vdd.n2552 vdd.n2505 9.3005
R22936 vdd.n2549 vdd.n2508 9.3005
R22937 vdd.n2546 vdd.n2511 9.3005
R22938 vdd.n2541 vdd.n2513 9.3005
R22939 vdd.n2538 vdd.n2516 9.3005
R22940 vdd.n2535 vdd.n2518 9.3005
R22941 vdd.n2533 vdd.n2521 9.3005
R22942 vdd.n2530 vdd.n2527 9.3005
R22943 vdd.n2526 vdd.n2525 9.3005
R22944 vdd.n2570 vdd.n235 9.3005
R22945 vdd.n2573 vdd.n231 9.3005
R22946 vdd.n2576 vdd.n229 9.3005
R22947 vdd.n2581 vdd.n227 9.3005
R22948 vdd.n2584 vdd.n223 9.3005
R22949 vdd.n222 vdd.n218 9.3005
R22950 vdd.n2588 vdd.n219 9.3005
R22951 vdd.n2591 vdd.n216 9.3005
R22952 vdd.n2594 vdd.n212 9.3005
R22953 vdd.n2597 vdd.n210 9.3005
R22954 vdd.n2600 vdd.n207 9.3005
R22955 vdd.n2603 vdd.n203 9.3005
R22956 vdd.n2606 vdd.n197 9.3005
R22957 vdd.n196 vdd.n192 9.3005
R22958 vdd.n2610 vdd.n193 9.3005
R22959 vdd.n2613 vdd.n190 9.3005
R22960 vdd.n2616 vdd.n188 9.3005
R22961 vdd.n2619 vdd.n185 9.3005
R22962 vdd.n2622 vdd.n183 9.3005
R22963 vdd.n2625 vdd.n179 9.3005
R22964 vdd.n2628 vdd.n177 9.3005
R22965 vdd.n2631 vdd.n172 9.3005
R22966 vdd.n171 vdd.n167 9.3005
R22967 vdd.n2635 vdd.n168 9.3005
R22968 vdd.n2638 vdd.n165 9.3005
R22969 vdd.n2641 vdd.n163 9.3005
R22970 vdd.n2644 vdd.n159 9.3005
R22971 vdd.n2647 vdd.n156 9.3005
R22972 vdd.n2651 vdd.n152 9.3005
R22973 vdd.n2803 vdd.n147 9.3005
R22974 vdd.n2800 vdd.n2654 9.3005
R22975 vdd.n2797 vdd.n2659 9.3005
R22976 vdd.n2796 vdd.n2661 9.3005
R22977 vdd.n2793 vdd.n2664 9.3005
R22978 vdd.n2790 vdd.n2667 9.3005
R22979 vdd.n2785 vdd.n2669 9.3005
R22980 vdd.n2782 vdd.n2672 9.3005
R22981 vdd.n2779 vdd.n2674 9.3005
R22982 vdd.n2774 vdd.n2676 9.3005
R22983 vdd.n2771 vdd.n2678 9.3005
R22984 vdd.n2768 vdd.n2681 9.3005
R22985 vdd.n2766 vdd.n2684 9.3005
R22986 vdd.n2763 vdd.n2762 9.3005
R22987 vdd.n2761 vdd.n2760 9.3005
R22988 vdd.n2757 vdd.n2688 9.3005
R22989 vdd.n2754 vdd.n2695 9.3005
R22990 vdd.n2751 vdd.n2699 9.3005
R22991 vdd.n2748 vdd.n2701 9.3005
R22992 vdd.n2745 vdd.n2703 9.3005
R22993 vdd.n2742 vdd.n2708 9.3005
R22994 vdd.n2741 vdd.n2710 9.3005
R22995 vdd.n2738 vdd.n2713 9.3005
R22996 vdd.n2735 vdd.n2716 9.3005
R22997 vdd.n2730 vdd.n2718 9.3005
R22998 vdd.n2727 vdd.n2725 9.3005
R22999 vdd.n2724 vdd.n2723 9.3005
R23000 vdd.n2817 vdd.n133 9.3005
R23001 vdd.n2820 vdd.n131 9.3005
R23002 vdd.n2823 vdd.n129 9.3005
R23003 vdd.n2826 vdd.n126 9.3005
R23004 vdd.n2829 vdd.n122 9.3005
R23005 vdd.n2832 vdd.n120 9.3005
R23006 vdd.n2835 vdd.n118 9.3005
R23007 vdd.n2838 vdd.n114 9.3005
R23008 vdd.n2841 vdd.n111 9.3005
R23009 vdd.n2846 vdd.n109 9.3005
R23010 vdd.n2850 vdd.n104 9.3005
R23011 vdd.n103 vdd.n98 9.3005
R23012 vdd.n2854 vdd.n99 9.3005
R23013 vdd.n2561 vdd.n2560 9.3005
R23014 vdd.n2559 vdd.n2493 9.3005
R23015 vdd.n2558 vdd.n2557 9.3005
R23016 vdd.n2554 vdd.n2495 9.3005
R23017 vdd.n2552 vdd.n2551 9.3005
R23018 vdd.n2550 vdd.n2549 9.3005
R23019 vdd.n2546 vdd.n2507 9.3005
R23020 vdd.n2541 vdd.n2540 9.3005
R23021 vdd.n2539 vdd.n2538 9.3005
R23022 vdd.n2535 vdd.n2515 9.3005
R23023 vdd.n2533 vdd.n2532 9.3005
R23024 vdd.n2531 vdd.n2530 9.3005
R23025 vdd.n2525 vdd.n2523 9.3005
R23026 vdd.n2570 vdd.n230 9.3005
R23027 vdd.n2574 vdd.n2573 9.3005
R23028 vdd.n2576 vdd.n2575 9.3005
R23029 vdd.n2581 vdd.n220 9.3005
R23030 vdd.n2585 vdd.n2584 9.3005
R23031 vdd.n2586 vdd.n218 9.3005
R23032 vdd.n2588 vdd.n2587 9.3005
R23033 vdd.n2591 vdd.n211 9.3005
R23034 vdd.n2595 vdd.n2594 9.3005
R23035 vdd.n2597 vdd.n2596 9.3005
R23036 vdd.n2600 vdd.n202 9.3005
R23037 vdd.n2604 vdd.n2603 9.3005
R23038 vdd.n2606 vdd.n2605 9.3005
R23039 vdd.n192 vdd.n191 9.3005
R23040 vdd.n2611 vdd.n2610 9.3005
R23041 vdd.n2613 vdd.n2612 9.3005
R23042 vdd.n2616 vdd.n184 9.3005
R23043 vdd.n2620 vdd.n2619 9.3005
R23044 vdd.n2622 vdd.n2621 9.3005
R23045 vdd.n2625 vdd.n176 9.3005
R23046 vdd.n2629 vdd.n2628 9.3005
R23047 vdd.n2631 vdd.n2630 9.3005
R23048 vdd.n167 vdd.n166 9.3005
R23049 vdd.n2636 vdd.n2635 9.3005
R23050 vdd.n2638 vdd.n2637 9.3005
R23051 vdd.n2641 vdd.n158 9.3005
R23052 vdd.n2645 vdd.n2644 9.3005
R23053 vdd.n2647 vdd.n2646 9.3005
R23054 vdd.n2652 vdd.n2651 9.3005
R23055 vdd.n2803 vdd.n2802 9.3005
R23056 vdd.n2801 vdd.n2800 9.3005
R23057 vdd.n2797 vdd.n2653 9.3005
R23058 vdd.n2796 vdd.n2795 9.3005
R23059 vdd.n2794 vdd.n2793 9.3005
R23060 vdd.n2790 vdd.n2663 9.3005
R23061 vdd.n2785 vdd.n2784 9.3005
R23062 vdd.n2783 vdd.n2782 9.3005
R23063 vdd.n2779 vdd.n2671 9.3005
R23064 vdd.n2774 vdd.n2773 9.3005
R23065 vdd.n2772 vdd.n2771 9.3005
R23066 vdd.n2768 vdd.n2677 9.3005
R23067 vdd.n2766 vdd.n2683 9.3005
R23068 vdd.n2763 vdd.n2686 9.3005
R23069 vdd.n2760 vdd.n2689 9.3005
R23070 vdd.n2757 vdd.n2756 9.3005
R23071 vdd.n2755 vdd.n2754 9.3005
R23072 vdd.n2751 vdd.n2694 9.3005
R23073 vdd.n2748 vdd.n2747 9.3005
R23074 vdd.n2746 vdd.n2745 9.3005
R23075 vdd.n2742 vdd.n2702 9.3005
R23076 vdd.n2741 vdd.n2740 9.3005
R23077 vdd.n2739 vdd.n2738 9.3005
R23078 vdd.n2735 vdd.n2712 9.3005
R23079 vdd.n2730 vdd.n2729 9.3005
R23080 vdd.n2728 vdd.n2727 9.3005
R23081 vdd.n2723 vdd.n2720 9.3005
R23082 vdd.n2817 vdd.n130 9.3005
R23083 vdd.n2821 vdd.n2820 9.3005
R23084 vdd.n2823 vdd.n2822 9.3005
R23085 vdd.n2826 vdd.n121 9.3005
R23086 vdd.n2830 vdd.n2829 9.3005
R23087 vdd.n2832 vdd.n2831 9.3005
R23088 vdd.n2835 vdd.n112 9.3005
R23089 vdd.n2839 vdd.n2838 9.3005
R23090 vdd.n2841 vdd.n2840 9.3005
R23091 vdd.n2846 vdd.n102 9.3005
R23092 vdd.n2851 vdd.n2850 9.3005
R23093 vdd.n2852 vdd.n98 9.3005
R23094 vdd.n2854 vdd.n2853 9.3005
R23095 vdd.n2760 vdd.n2759 9.3005
R23096 vdd.n2764 vdd.n2763 9.3005
R23097 vdd.n2766 vdd.n2765 9.3005
R23098 vdd.n2810 vdd.n97 9.3005
R23099 vdd.n1903 vdd.n344 9.3005
R23100 vdd.n348 vdd.n347 9.3005
R23101 vdd.n2318 vdd.n317 9.3005
R23102 vdd.n2315 vdd.n322 9.3005
R23103 vdd.n2314 vdd.n324 9.3005
R23104 vdd.n2311 vdd.n328 9.3005
R23105 vdd.n2308 vdd.n332 9.3005
R23106 vdd.n2056 vdd.n333 9.3005
R23107 vdd.n2062 vdd.n2061 9.3005
R23108 vdd.n2064 vdd.n2063 9.3005
R23109 vdd.n2067 vdd.n2046 9.3005
R23110 vdd.n2071 vdd.n2070 9.3005
R23111 vdd.n2072 vdd.n2044 9.3005
R23112 vdd.n2074 vdd.n2073 9.3005
R23113 vdd.n2077 vdd.n2039 9.3005
R23114 vdd.n2081 vdd.n2080 9.3005
R23115 vdd.n2083 vdd.n2082 9.3005
R23116 vdd.n2086 vdd.n2032 9.3005
R23117 vdd.n2090 vdd.n2089 9.3005
R23118 vdd.n2092 vdd.n2091 9.3005
R23119 vdd.n2095 vdd.n2029 9.3005
R23120 vdd.n2028 vdd.n2022 9.3005
R23121 vdd.n2099 vdd.n2019 9.3005
R23122 vdd.n2103 vdd.n2102 9.3005
R23123 vdd.n2105 vdd.n2104 9.3005
R23124 vdd.n2108 vdd.n2013 9.3005
R23125 vdd.n2112 vdd.n2111 9.3005
R23126 vdd.n2114 vdd.n2113 9.3005
R23127 vdd.n2117 vdd.n2005 9.3005
R23128 vdd.n2122 vdd.n2121 9.3005
R23129 vdd.n2123 vdd.n2003 9.3005
R23130 vdd.n2125 vdd.n2124 9.3005
R23131 vdd.n2128 vdd.n1998 9.3005
R23132 vdd.n2132 vdd.n2131 9.3005
R23133 vdd.n2134 vdd.n2133 9.3005
R23134 vdd.n2137 vdd.n1992 9.3005
R23135 vdd.n2141 vdd.n2140 9.3005
R23136 vdd.n2143 vdd.n2142 9.3005
R23137 vdd.n2146 vdd.n1989 9.3005
R23138 vdd.n1988 vdd.n1983 9.3005
R23139 vdd.n2150 vdd.n1980 9.3005
R23140 vdd.n2154 vdd.n2153 9.3005
R23141 vdd.n2156 vdd.n2155 9.3005
R23142 vdd.n1903 vdd.n350 9.3005
R23143 vdd.n349 vdd.n348 9.3005
R23144 vdd.n2318 vdd.n2317 9.3005
R23145 vdd.n2316 vdd.n2315 9.3005
R23146 vdd.n2314 vdd.n320 9.3005
R23147 vdd.n2311 vdd.n2310 9.3005
R23148 vdd.n2309 vdd.n2308 9.3005
R23149 vdd.n333 vdd.n330 9.3005
R23150 vdd.n2061 vdd.n2054 9.3005
R23151 vdd.n2065 vdd.n2064 9.3005
R23152 vdd.n2067 vdd.n2066 9.3005
R23153 vdd.n2070 vdd.n2051 9.3005
R23154 vdd.n2050 vdd.n2044 9.3005
R23155 vdd.n2074 vdd.n2041 9.3005
R23156 vdd.n2078 vdd.n2077 9.3005
R23157 vdd.n2080 vdd.n2079 9.3005
R23158 vdd.n2083 vdd.n2034 9.3005
R23159 vdd.n2087 vdd.n2086 9.3005
R23160 vdd.n2089 vdd.n2088 9.3005
R23161 vdd.n2092 vdd.n2024 9.3005
R23162 vdd.n2096 vdd.n2095 9.3005
R23163 vdd.n2097 vdd.n2022 9.3005
R23164 vdd.n2099 vdd.n2098 9.3005
R23165 vdd.n2102 vdd.n2017 9.3005
R23166 vdd.n2106 vdd.n2105 9.3005
R23167 vdd.n2108 vdd.n2107 9.3005
R23168 vdd.n2111 vdd.n2011 9.3005
R23169 vdd.n2115 vdd.n2114 9.3005
R23170 vdd.n2117 vdd.n2116 9.3005
R23171 vdd.n2121 vdd.n2008 9.3005
R23172 vdd.n2003 vdd.n2002 9.3005
R23173 vdd.n2126 vdd.n2125 9.3005
R23174 vdd.n2128 vdd.n2127 9.3005
R23175 vdd.n2131 vdd.n1996 9.3005
R23176 vdd.n2135 vdd.n2134 9.3005
R23177 vdd.n2137 vdd.n2136 9.3005
R23178 vdd.n2140 vdd.n1990 9.3005
R23179 vdd.n2144 vdd.n2143 9.3005
R23180 vdd.n2146 vdd.n2145 9.3005
R23181 vdd.n1983 vdd.n1982 9.3005
R23182 vdd.n2151 vdd.n2150 9.3005
R23183 vdd.n2153 vdd.n2152 9.3005
R23184 vdd.n2156 vdd.n1978 9.3005
R23185 vdd.n1903 vdd.n343 9.3005
R23186 vdd.n348 vdd.n346 9.3005
R23187 vdd.n2318 vdd.n316 9.3005
R23188 vdd.n2315 vdd.n321 9.3005
R23189 vdd.n2314 vdd.n323 9.3005
R23190 vdd.n2311 vdd.n327 9.3005
R23191 vdd.n2308 vdd.n331 9.3005
R23192 vdd.n2057 vdd.n333 9.3005
R23193 vdd.n2061 vdd.n2058 9.3005
R23194 vdd.n2064 vdd.n2055 9.3005
R23195 vdd.n2067 vdd.n2053 9.3005
R23196 vdd.n2070 vdd.n2049 9.3005
R23197 vdd.n2048 vdd.n2044 9.3005
R23198 vdd.n2074 vdd.n2045 9.3005
R23199 vdd.n2077 vdd.n2042 9.3005
R23200 vdd.n2080 vdd.n2040 9.3005
R23201 vdd.n2083 vdd.n2038 9.3005
R23202 vdd.n2086 vdd.n2035 9.3005
R23203 vdd.n2089 vdd.n2033 9.3005
R23204 vdd.n2092 vdd.n2031 9.3005
R23205 vdd.n2095 vdd.n2026 9.3005
R23206 vdd.n2025 vdd.n2022 9.3005
R23207 vdd.n2099 vdd.n2023 9.3005
R23208 vdd.n2102 vdd.n2020 9.3005
R23209 vdd.n2105 vdd.n2018 9.3005
R23210 vdd.n2108 vdd.n2016 9.3005
R23211 vdd.n2111 vdd.n2014 9.3005
R23212 vdd.n2114 vdd.n2012 9.3005
R23213 vdd.n2117 vdd.n2010 9.3005
R23214 vdd.n2121 vdd.n2007 9.3005
R23215 vdd.n2006 vdd.n2003 9.3005
R23216 vdd.n2125 vdd.n2004 9.3005
R23217 vdd.n2128 vdd.n2001 9.3005
R23218 vdd.n2131 vdd.n1999 9.3005
R23219 vdd.n2134 vdd.n1997 9.3005
R23220 vdd.n2137 vdd.n1995 9.3005
R23221 vdd.n2140 vdd.n1993 9.3005
R23222 vdd.n2143 vdd.n1991 9.3005
R23223 vdd.n2146 vdd.n1987 9.3005
R23224 vdd.n1986 vdd.n1983 9.3005
R23225 vdd.n2150 vdd.n1984 9.3005
R23226 vdd.n2153 vdd.n1981 9.3005
R23227 vdd.n2156 vdd.n1977 9.3005
R23228 vdd.n1903 vdd.n1902 9.3005
R23229 vdd.n348 vdd.n313 9.3005
R23230 vdd.n2319 vdd.n2318 9.3005
R23231 vdd.n2315 vdd.n314 9.3005
R23232 vdd.n2314 vdd.n2313 9.3005
R23233 vdd.n2312 vdd.n2311 9.3005
R23234 vdd.n2308 vdd.n326 9.3005
R23235 vdd.n2059 vdd.n333 9.3005
R23236 vdd.n2061 vdd.n2060 9.3005
R23237 vdd.n2064 vdd.n2052 9.3005
R23238 vdd.n2068 vdd.n2067 9.3005
R23239 vdd.n2070 vdd.n2069 9.3005
R23240 vdd.n2044 vdd.n2043 9.3005
R23241 vdd.n2075 vdd.n2074 9.3005
R23242 vdd.n2077 vdd.n2076 9.3005
R23243 vdd.n2080 vdd.n2036 9.3005
R23244 vdd.n2084 vdd.n2083 9.3005
R23245 vdd.n2086 vdd.n2085 9.3005
R23246 vdd.n2089 vdd.n2030 9.3005
R23247 vdd.n2093 vdd.n2092 9.3005
R23248 vdd.n2095 vdd.n2094 9.3005
R23249 vdd.n2022 vdd.n2021 9.3005
R23250 vdd.n2100 vdd.n2099 9.3005
R23251 vdd.n2102 vdd.n2101 9.3005
R23252 vdd.n2105 vdd.n2015 9.3005
R23253 vdd.n2109 vdd.n2108 9.3005
R23254 vdd.n2111 vdd.n2110 9.3005
R23255 vdd.n2114 vdd.n2009 9.3005
R23256 vdd.n2118 vdd.n2117 9.3005
R23257 vdd.n2121 vdd.n2120 9.3005
R23258 vdd.n2119 vdd.n2003 9.3005
R23259 vdd.n2125 vdd.n2000 9.3005
R23260 vdd.n2129 vdd.n2128 9.3005
R23261 vdd.n2131 vdd.n2130 9.3005
R23262 vdd.n2134 vdd.n1994 9.3005
R23263 vdd.n2138 vdd.n2137 9.3005
R23264 vdd.n2140 vdd.n2139 9.3005
R23265 vdd.n2143 vdd.n1985 9.3005
R23266 vdd.n2147 vdd.n2146 9.3005
R23267 vdd.n2148 vdd.n1983 9.3005
R23268 vdd.n2150 vdd.n2149 9.3005
R23269 vdd.n2153 vdd.n1979 9.3005
R23270 vdd.n2157 vdd.n2156 9.3005
R23271 vdd.n2158 vdd.n240 9.3005
R23272 vdd.n1796 vdd.n449 9.3005
R23273 vdd.n1800 vdd.n1799 9.3005
R23274 vdd.n1802 vdd.n1801 9.3005
R23275 vdd.n1805 vdd.n440 9.3005
R23276 vdd.n1809 vdd.n1808 9.3005
R23277 vdd.n1812 vdd.n1811 9.3005
R23278 vdd.n1815 vdd.n427 9.3005
R23279 vdd.n1819 vdd.n1818 9.3005
R23280 vdd.n1820 vdd.n425 9.3005
R23281 vdd.n1822 vdd.n1821 9.3005
R23282 vdd.n1825 vdd.n418 9.3005
R23283 vdd.n1829 vdd.n1828 9.3005
R23284 vdd.n1831 vdd.n1830 9.3005
R23285 vdd.n1834 vdd.n409 9.3005
R23286 vdd.n1838 vdd.n1837 9.3005
R23287 vdd.n1840 vdd.n1839 9.3005
R23288 vdd.n1843 vdd.n404 9.3005
R23289 vdd.n403 vdd.n397 9.3005
R23290 vdd.n1847 vdd.n393 9.3005
R23291 vdd.n1851 vdd.n1850 9.3005
R23292 vdd.n1853 vdd.n1852 9.3005
R23293 vdd.n1856 vdd.n384 9.3005
R23294 vdd.n1860 vdd.n1859 9.3005
R23295 vdd.n1862 vdd.n1861 9.3005
R23296 vdd.n1865 vdd.n380 9.3005
R23297 vdd.n1868 vdd.n375 9.3005
R23298 vdd.n374 vdd.n353 9.3005
R23299 vdd.n1899 vdd.n357 9.3005
R23300 vdd.n1799 vdd.n446 9.3005
R23301 vdd.n1803 vdd.n1802 9.3005
R23302 vdd.n1805 vdd.n1804 9.3005
R23303 vdd.n1808 vdd.n437 9.3005
R23304 vdd.n1813 vdd.n1812 9.3005
R23305 vdd.n1815 vdd.n1814 9.3005
R23306 vdd.n1818 vdd.n433 9.3005
R23307 vdd.n432 vdd.n425 9.3005
R23308 vdd.n1822 vdd.n421 9.3005
R23309 vdd.n1826 vdd.n1825 9.3005
R23310 vdd.n1828 vdd.n1827 9.3005
R23311 vdd.n1831 vdd.n412 9.3005
R23312 vdd.n1835 vdd.n1834 9.3005
R23313 vdd.n1837 vdd.n1836 9.3005
R23314 vdd.n1840 vdd.n399 9.3005
R23315 vdd.n1844 vdd.n1843 9.3005
R23316 vdd.n1845 vdd.n397 9.3005
R23317 vdd.n1847 vdd.n1846 9.3005
R23318 vdd.n1850 vdd.n390 9.3005
R23319 vdd.n1854 vdd.n1853 9.3005
R23320 vdd.n1856 vdd.n1855 9.3005
R23321 vdd.n1859 vdd.n381 9.3005
R23322 vdd.n1863 vdd.n1862 9.3005
R23323 vdd.n1865 vdd.n1864 9.3005
R23324 vdd.n1868 vdd.n376 9.3005
R23325 vdd.n359 vdd.n353 9.3005
R23326 vdd.n1899 vdd.n1898 9.3005
R23327 vdd.n1799 vdd.n451 9.3005
R23328 vdd.n1802 vdd.n448 9.3005
R23329 vdd.n1805 vdd.n445 9.3005
R23330 vdd.n1808 vdd.n442 9.3005
R23331 vdd.n1812 vdd.n439 9.3005
R23332 vdd.n1815 vdd.n436 9.3005
R23333 vdd.n1818 vdd.n430 9.3005
R23334 vdd.n429 vdd.n425 9.3005
R23335 vdd.n1822 vdd.n426 9.3005
R23336 vdd.n1825 vdd.n423 9.3005
R23337 vdd.n1828 vdd.n420 9.3005
R23338 vdd.n1831 vdd.n417 9.3005
R23339 vdd.n1834 vdd.n414 9.3005
R23340 vdd.n1837 vdd.n411 9.3005
R23341 vdd.n1840 vdd.n408 9.3005
R23342 vdd.n1843 vdd.n402 9.3005
R23343 vdd.n401 vdd.n397 9.3005
R23344 vdd.n1847 vdd.n398 9.3005
R23345 vdd.n1850 vdd.n395 9.3005
R23346 vdd.n1853 vdd.n392 9.3005
R23347 vdd.n1856 vdd.n389 9.3005
R23348 vdd.n1859 vdd.n386 9.3005
R23349 vdd.n1862 vdd.n383 9.3005
R23350 vdd.n1865 vdd.n379 9.3005
R23351 vdd.n1868 vdd.n373 9.3005
R23352 vdd.n372 vdd.n353 9.3005
R23353 vdd.n1899 vdd.n354 9.3005
R23354 vdd.n1799 vdd.n1798 9.3005
R23355 vdd.n1802 vdd.n443 9.3005
R23356 vdd.n1806 vdd.n1805 9.3005
R23357 vdd.n1808 vdd.n1807 9.3005
R23358 vdd.n1812 vdd.n434 9.3005
R23359 vdd.n1816 vdd.n1815 9.3005
R23360 vdd.n1818 vdd.n1817 9.3005
R23361 vdd.n425 vdd.n424 9.3005
R23362 vdd.n1823 vdd.n1822 9.3005
R23363 vdd.n1825 vdd.n1824 9.3005
R23364 vdd.n1828 vdd.n415 9.3005
R23365 vdd.n1832 vdd.n1831 9.3005
R23366 vdd.n1834 vdd.n1833 9.3005
R23367 vdd.n1837 vdd.n406 9.3005
R23368 vdd.n1841 vdd.n1840 9.3005
R23369 vdd.n1843 vdd.n1842 9.3005
R23370 vdd.n397 vdd.n396 9.3005
R23371 vdd.n1848 vdd.n1847 9.3005
R23372 vdd.n1850 vdd.n1849 9.3005
R23373 vdd.n1853 vdd.n387 9.3005
R23374 vdd.n1857 vdd.n1856 9.3005
R23375 vdd.n1859 vdd.n1858 9.3005
R23376 vdd.n1862 vdd.n377 9.3005
R23377 vdd.n1866 vdd.n1865 9.3005
R23378 vdd.n1868 vdd.n1867 9.3005
R23379 vdd.n353 vdd.n352 9.3005
R23380 vdd.n1900 vdd.n1899 9.3005
R23381 vdd.n1796 vdd.n1795 9.3005
R23382 vdd.n1796 vdd.n454 9.3005
R23383 vdd.n1797 vdd.n1796 9.3005
R23384 vdd.n291 vdd.n290 9.3005
R23385 vdd.n2357 vdd.n2356 9.3005
R23386 vdd.n2358 vdd.n289 9.3005
R23387 vdd.n2360 vdd.n2359 9.3005
R23388 vdd.n287 vdd.n286 9.3005
R23389 vdd.n2368 vdd.n2367 9.3005
R23390 vdd.n2370 vdd.n2369 9.3005
R23391 vdd.n283 vdd.n282 9.3005
R23392 vdd.n2378 vdd.n2377 9.3005
R23393 vdd.n2380 vdd.n2379 9.3005
R23394 vdd.n279 vdd.n278 9.3005
R23395 vdd.n2389 vdd.n2388 9.3005
R23396 vdd.n2390 vdd.n277 9.3005
R23397 vdd.n2392 vdd.n2391 9.3005
R23398 vdd.n275 vdd.n274 9.3005
R23399 vdd.n2400 vdd.n2399 9.3005
R23400 vdd.n2402 vdd.n2401 9.3005
R23401 vdd.n271 vdd.n270 9.3005
R23402 vdd.n2410 vdd.n2409 9.3005
R23403 vdd.n2413 vdd.n2412 9.3005
R23404 vdd.n2411 vdd.n267 9.3005
R23405 vdd.n2422 vdd.n2421 9.3005
R23406 vdd.n2423 vdd.n265 9.3005
R23407 vdd.n2425 vdd.n2424 9.3005
R23408 vdd.n263 vdd.n262 9.3005
R23409 vdd.n2433 vdd.n2432 9.3005
R23410 vdd.n2435 vdd.n2434 9.3005
R23411 vdd.n259 vdd.n258 9.3005
R23412 vdd.n2443 vdd.n2442 9.3005
R23413 vdd.n2445 vdd.n2444 9.3005
R23414 vdd.n255 vdd.n254 9.3005
R23415 vdd.n2454 vdd.n2453 9.3005
R23416 vdd.n2455 vdd.n253 9.3005
R23417 vdd.n2457 vdd.n2456 9.3005
R23418 vdd.n251 vdd.n250 9.3005
R23419 vdd.n2465 vdd.n2464 9.3005
R23420 vdd.n2467 vdd.n2466 9.3005
R23421 vdd.n246 vdd.n245 9.3005
R23422 vdd.n2474 vdd.n2473 9.3005
R23423 vdd.n2476 vdd.n2475 9.3005
R23424 vdd.n242 vdd.n241 9.3005
R23425 vdd.n2348 vdd.n2347 9.3005
R23426 vdd.n2345 vdd.n2344 9.3005
R23427 vdd.n1811 vdd.n1810 9.03579
R23428 vdd.n1114 vdd.n1112 8.65932
R23429 vdd.n1231 vdd.n1230 8.28285
R23430 vdd.n2327 vdd.n2326 7.70883
R23431 vdd.n2326 vdd.n2325 7.70883
R23432 vdd.n1301 vdd.n1300 7.70883
R23433 vdd.n1300 vdd.n617 7.70883
R23434 vdd.n2323 vdd.n294 7.70883
R23435 vdd.n2324 vdd.n2323 7.70883
R23436 vdd.n1509 vdd.n1508 7.70883
R23437 vdd.n1510 vdd.n1509 7.70883
R23438 vdd.n1162 vdd.n1161 7.70883
R23439 vdd.n2483 vdd.n2482 7.70883
R23440 vdd.n2484 vdd.n2483 7.70883
R23441 vdd.n357 vdd.n307 7.15344
R23442 vdd.n2813 vdd.n2812 6.85235
R23443 vdd.t278 vdd.n2813 6.85235
R23444 vdd.n2808 vdd.n2807 6.85235
R23445 vdd.n2807 vdd.t191 6.85235
R23446 vdd.n2566 vdd.n2565 6.85235
R23447 vdd.t164 vdd.n2566 6.85235
R23448 vdd.n2568 vdd.n2567 6.85235
R23449 vdd.n2567 vdd.t164 6.85235
R23450 vdd.n2806 vdd.n2805 6.85235
R23451 vdd.t191 vdd.n2806 6.85235
R23452 vdd.n2815 vdd.n2814 6.85235
R23453 vdd.n2814 vdd.t278 6.85235
R23454 vdd.n2563 vdd.n2562 6.77697
R23455 vdd.n2764 vdd.n2685 6.77697
R23456 vdd.n1657 vdd.n526 6.77697
R23457 vdd.n2344 vdd.n2343 6.64659
R23458 vdd.n1507 vdd.n1506 6.4005
R23459 vdd.n2411 vdd.n266 6.02403
R23460 vdd.n2204 vdd.n2203 4.5005
R23461 vdd.n2197 vdd.n2183 4.5005
R23462 vdd.n2207 vdd.n2192 4.5005
R23463 vdd.n2207 vdd.n2188 4.5005
R23464 vdd.n2207 vdd.n2195 4.5005
R23465 vdd.n2207 vdd.n2187 4.5005
R23466 vdd.n2207 vdd.n2197 4.5005
R23467 vdd.n1642 vdd.n1641 4.5005
R23468 vdd.n1661 vdd.n1660 4.5005
R23469 vdd.n1642 vdd.n515 4.5005
R23470 vdd.n1601 vdd.n515 4.5005
R23471 vdd.n1606 vdd.n515 4.5005
R23472 vdd.n1608 vdd.n515 4.5005
R23473 vdd.n1610 vdd.n515 4.5005
R23474 vdd.n1612 vdd.n515 4.5005
R23475 vdd.n1614 vdd.n515 4.5005
R23476 vdd.n1605 vdd.n515 4.5005
R23477 vdd.n1618 vdd.n515 4.5005
R23478 vdd.n518 vdd.n515 4.5005
R23479 vdd.n1661 vdd.n515 4.5005
R23480 vdd.n1886 vdd.n341 4.5005
R23481 vdd.n1886 vdd.n364 4.5005
R23482 vdd.n367 vdd.n364 4.5005
R23483 vdd.n1893 vdd.n367 4.5005
R23484 vdd.n1890 vdd.n367 4.5005
R23485 vdd.n1888 vdd.n367 4.5005
R23486 vdd.n1875 vdd.n367 4.5005
R23487 vdd.n1878 vdd.n367 4.5005
R23488 vdd.n1880 vdd.n367 4.5005
R23489 vdd.n1877 vdd.n367 4.5005
R23490 vdd.n1884 vdd.n367 4.5005
R23491 vdd.n367 vdd.n341 4.5005
R23492 vdd.n2342 vdd.n2341 4.5005
R23493 vdd.n1492 vdd.n1295 4.5005
R23494 vdd.n1502 vdd.n1295 4.5005
R23495 vdd.n2339 vdd.n2338 4.5005
R23496 vdd.n2649 vdd.n141 4.20505
R23497 vdd.n155 vdd.n141 4.20505
R23498 vdd.n149 vdd.n141 4.20505
R23499 vdd.n1511 vdd.n580 4.20505
R23500 vdd.n2322 vdd.n310 4.20505
R23501 vdd.n1112 vdd.n618 4.20505
R23502 vdd.t80 vdd.n618 4.20505
R23503 vdd.n1810 vdd.n308 4.20505
R23504 vdd.t215 vdd.n308 4.20505
R23505 vdd.n2027 vdd.n238 4.20505
R23506 vdd.t96 vdd.n238 4.20505
R23507 vdd.n1230 vdd.n619 4.20505
R23508 vdd.t80 vdd.n619 4.20505
R23509 vdd.n1335 vdd.n309 4.20505
R23510 vdd.t215 vdd.n309 4.20505
R23511 vdd.n266 vdd.n239 4.20505
R23512 vdd.t96 vdd.n239 4.20505
R23513 vdd.n2346 vdd.n2345 4.14168
R23514 vdd.n355 vdd.n344 3.76521
R23515 vdd.n2205 vdd.n2204 3.47482
R23516 vdd.n2207 vdd.n2186 3.46142
R23517 vdd.n2186 vdd.n2182 3.46142
R23518 vdd.n2206 vdd.n2183 3.4105
R23519 vdd.n2208 vdd.n2183 3.4105
R23520 vdd.n2183 vdd.n2178 3.4105
R23521 vdd.n2185 vdd.n2183 3.4105
R23522 vdd.n2206 vdd.n2182 3.4105
R23523 vdd.n2208 vdd.n2182 3.4105
R23524 vdd.n2182 vdd.n2178 3.4105
R23525 vdd.n2185 vdd.n2182 3.4105
R23526 vdd.n2200 vdd.n2182 3.4105
R23527 vdd.n2207 vdd.n2200 3.4105
R23528 vdd.n2207 vdd.n2185 3.4105
R23529 vdd.n2207 vdd.n2178 3.4105
R23530 vdd.n2208 vdd.n2207 3.4105
R23531 vdd.n2207 vdd.n2206 3.4105
R23532 vdd.n778 vdd.n768 3.4105
R23533 vdd.n772 vdd.n768 3.4105
R23534 vdd.n778 vdd.n777 3.4105
R23535 vdd.n2816 vdd.n2815 3.38874
R23536 vdd.n1632 vdd.n525 3.38874
R23537 vdd.n1488 vdd.n1302 3.01226
R23538 vdd.n2190 vdd.n2189 2.26334
R23539 vdd.n2480 vdd.n2479 2.25519
R23540 vdd.n2203 vdd.n2201 2.25201
R23541 vdd.n1167 vdd.n1166 2.2505
R23542 vdd.n1169 vdd.n1168 2.2505
R23543 vdd.n684 vdd.n683 2.2505
R23544 vdd.n1175 vdd.n1174 2.2505
R23545 vdd.n1178 vdd.n1177 2.2505
R23546 vdd.n679 vdd.n678 2.2505
R23547 vdd.n1184 vdd.n1183 2.2505
R23548 vdd.n1187 vdd.n1186 2.2505
R23549 vdd.n1188 vdd.n673 2.2505
R23550 vdd.n1195 vdd.n1194 2.2505
R23551 vdd.n1198 vdd.n1197 2.2505
R23552 vdd.n669 vdd.n668 2.2505
R23553 vdd.n1204 vdd.n1203 2.2505
R23554 vdd.n1207 vdd.n1206 2.2505
R23555 vdd.n664 vdd.n663 2.2505
R23556 vdd.n1213 vdd.n1212 2.2505
R23557 vdd.n1216 vdd.n1215 2.2505
R23558 vdd.n1217 vdd.n658 2.2505
R23559 vdd.n1224 vdd.n1223 2.2505
R23560 vdd.n1227 vdd.n1226 2.2505
R23561 vdd.n654 vdd.n653 2.2505
R23562 vdd.n1234 vdd.n1233 2.2505
R23563 vdd.n1237 vdd.n1236 2.2505
R23564 vdd.n649 vdd.n648 2.2505
R23565 vdd.n1243 vdd.n1242 2.2505
R23566 vdd.n1246 vdd.n1245 2.2505
R23567 vdd.n1247 vdd.n643 2.2505
R23568 vdd.n1254 vdd.n1253 2.2505
R23569 vdd.n1257 vdd.n1256 2.2505
R23570 vdd.n639 vdd.n638 2.2505
R23571 vdd.n1263 vdd.n1262 2.2505
R23572 vdd.n1266 vdd.n1265 2.2505
R23573 vdd.n1264 vdd.n634 2.2505
R23574 vdd.n1273 vdd.n1272 2.2505
R23575 vdd.n1274 vdd.n631 2.2505
R23576 vdd.n1276 vdd.n1275 2.2505
R23577 vdd.n1283 vdd.n1282 2.2505
R23578 vdd.n1286 vdd.n1285 2.2505
R23579 vdd.n1284 vdd.n624 2.2505
R23580 vdd.n1293 vdd.n1292 2.2505
R23581 vdd.n1294 vdd.n622 2.2505
R23582 vdd.n1504 vdd.n1503 2.2505
R23583 vdd.n1491 vdd.n1490 2.2505
R23584 vdd.n1299 vdd.n1298 2.2505
R23585 vdd.n1484 vdd.n1483 2.2505
R23586 vdd.n1481 vdd.n1480 2.2505
R23587 vdd.n1307 vdd.n1306 2.2505
R23588 vdd.n1475 vdd.n1474 2.2505
R23589 vdd.n1472 vdd.n1471 2.2505
R23590 vdd.n1313 vdd.n1312 2.2505
R23591 vdd.n1466 vdd.n1465 2.2505
R23592 vdd.n1463 vdd.n1462 2.2505
R23593 vdd.n1318 vdd.n1317 2.2505
R23594 vdd.n1456 vdd.n1455 2.2505
R23595 vdd.n1453 vdd.n1452 2.2505
R23596 vdd.n1323 vdd.n1322 2.2505
R23597 vdd.n1447 vdd.n1446 2.2505
R23598 vdd.n1444 vdd.n1443 2.2505
R23599 vdd.n1329 vdd.n1328 2.2505
R23600 vdd.n1438 vdd.n1437 2.2505
R23601 vdd.n1435 vdd.n1434 2.2505
R23602 vdd.n1334 vdd.n1333 2.2505
R23603 vdd.n1340 vdd.n1336 2.2505
R23604 vdd.n1425 vdd.n1424 2.2505
R23605 vdd.n1423 vdd.n1422 2.2505
R23606 vdd.n1343 vdd.n1342 2.2505
R23607 vdd.n1417 vdd.n1416 2.2505
R23608 vdd.n1415 vdd.n1414 2.2505
R23609 vdd.n1349 vdd.n1348 2.2505
R23610 vdd.n1409 vdd.n1408 2.2505
R23611 vdd.n1407 vdd.n1406 2.2505
R23612 vdd.n1357 vdd.n1354 2.2505
R23613 vdd.n1400 vdd.n1399 2.2505
R23614 vdd.n1398 vdd.n1397 2.2505
R23615 vdd.n1362 vdd.n1361 2.2505
R23616 vdd.n1392 vdd.n1391 2.2505
R23617 vdd.n1390 vdd.n1389 2.2505
R23618 vdd.n1368 vdd.n1367 2.2505
R23619 vdd.n1384 vdd.n1383 2.2505
R23620 vdd.n1382 vdd.n1381 2.2505
R23621 vdd.n1376 vdd.n1374 2.2505
R23622 vdd.n305 vdd.n304 2.2505
R23623 vdd.n2333 vdd.n2332 2.2505
R23624 vdd.n293 vdd.n292 2.2505
R23625 vdd.n2350 vdd.n2349 2.2505
R23626 vdd.n2354 vdd.n2353 2.2505
R23627 vdd.n2355 vdd.n288 2.2505
R23628 vdd.n2362 vdd.n2361 2.2505
R23629 vdd.n2366 vdd.n2365 2.2505
R23630 vdd.n285 vdd.n284 2.2505
R23631 vdd.n2372 vdd.n2371 2.2505
R23632 vdd.n2376 vdd.n2375 2.2505
R23633 vdd.n281 vdd.n280 2.2505
R23634 vdd.n2382 vdd.n2381 2.2505
R23635 vdd.n2386 vdd.n2385 2.2505
R23636 vdd.n2387 vdd.n276 2.2505
R23637 vdd.n2394 vdd.n2393 2.2505
R23638 vdd.n2398 vdd.n2397 2.2505
R23639 vdd.n273 vdd.n272 2.2505
R23640 vdd.n2404 vdd.n2403 2.2505
R23641 vdd.n2408 vdd.n2407 2.2505
R23642 vdd.n269 vdd.n268 2.2505
R23643 vdd.n2415 vdd.n2414 2.2505
R23644 vdd.n2419 vdd.n2418 2.2505
R23645 vdd.n2420 vdd.n264 2.2505
R23646 vdd.n2427 vdd.n2426 2.2505
R23647 vdd.n2431 vdd.n2430 2.2505
R23648 vdd.n261 vdd.n260 2.2505
R23649 vdd.n2437 vdd.n2436 2.2505
R23650 vdd.n2441 vdd.n2440 2.2505
R23651 vdd.n257 vdd.n256 2.2505
R23652 vdd.n2447 vdd.n2446 2.2505
R23653 vdd.n2451 vdd.n2450 2.2505
R23654 vdd.n2452 vdd.n252 2.2505
R23655 vdd.n2459 vdd.n2458 2.2505
R23656 vdd.n2463 vdd.n2462 2.2505
R23657 vdd.n249 vdd.n248 2.2505
R23658 vdd.n2469 vdd.n2468 2.2505
R23659 vdd.n2472 vdd.n2471 2.2505
R23660 vdd.n244 vdd.n243 2.2505
R23661 vdd.n2478 vdd.n2477 2.2505
R23662 vdd.n871 vdd.n870 2.2505
R23663 vdd.n845 vdd.n843 2.2505
R23664 vdd.n865 vdd.n864 2.2505
R23665 vdd.n863 vdd.n862 2.2505
R23666 vdd.n853 vdd.n849 2.2505
R23667 vdd.n855 vdd.n854 2.2505
R23668 vdd.n851 vdd.n687 2.2505
R23669 vdd.n1641 vdd.n516 2.2419
R23670 vdd.n1641 vdd.n1619 2.2419
R23671 vdd.n1641 vdd.n1604 2.2419
R23672 vdd.n1641 vdd.n1603 2.2419
R23673 vdd.n1641 vdd.n1602 2.2419
R23674 vdd.n1660 vdd.n523 2.2419
R23675 vdd.n1660 vdd.n522 2.2419
R23676 vdd.n1660 vdd.n520 2.2419
R23677 vdd.n1660 vdd.n519 2.2419
R23678 vdd.n1886 vdd.n1885 2.2419
R23679 vdd.n1886 vdd.n1876 2.2419
R23680 vdd.n1887 vdd.n1886 2.2419
R23681 vdd.n1886 vdd.n368 2.2419
R23682 vdd.n1895 vdd.n1894 2.2419
R23683 vdd.n1895 vdd.n362 2.2419
R23684 vdd.n1895 vdd.n361 2.2419
R23685 vdd.n1895 vdd.n360 2.2419
R23686 vdd.n1660 vdd.n521 2.24179
R23687 vdd.n1895 vdd.n363 2.24179
R23688 vdd.n2194 vdd.n2183 2.24131
R23689 vdd.n2191 vdd.n2183 2.24131
R23690 vdd.n2196 vdd.n2182 2.24131
R23691 vdd.n2193 vdd.n2182 2.24131
R23692 vdd.n2190 vdd.n2182 2.24131
R23693 vdd.n2342 vdd.n302 2.23548
R23694 vdd.n2342 vdd.n301 2.23548
R23695 vdd.n2342 vdd.n300 2.23548
R23696 vdd.n2342 vdd.n299 2.23548
R23697 vdd.n2342 vdd.n298 2.23548
R23698 vdd.n1494 vdd.n1295 2.23548
R23699 vdd.n1496 vdd.n1295 2.23548
R23700 vdd.n1498 vdd.n1295 2.23548
R23701 vdd.n1296 vdd.n1295 2.23548
R23702 vdd.n1501 vdd.n1500 2.23548
R23703 vdd.n1500 vdd.n1499 2.23548
R23704 vdd.n1500 vdd.n1497 2.23548
R23705 vdd.n1500 vdd.n1495 2.23548
R23706 vdd.n1500 vdd.n1493 2.23548
R23707 vdd.n2340 vdd.n2339 2.23548
R23708 vdd.n2339 vdd.n2334 2.23548
R23709 vdd.n2339 vdd.n2335 2.23548
R23710 vdd.n2339 vdd.n2336 2.23548
R23711 vdd.n2339 vdd.n2337 2.23548
R23712 vdd.n1513 vdd.n1512 2.10277
R23713 vdd.n1512 vdd.n1511 2.10277
R23714 vdd.n319 vdd.n311 2.10277
R23715 vdd.n2322 vdd.n311 2.10277
R23716 vdd.n604 vdd.n312 2.10277
R23717 vdd.n1511 vdd.n312 2.10277
R23718 vdd.n2321 vdd.n2320 2.10277
R23719 vdd.n2322 vdd.n2321 2.10277
R23720 vdd.n2027 vdd.n2019 1.88285
R23721 vdd.n2205 vdd.n2201 1.72167
R23722 vdd.n2198 vdd.n2183 1.70434
R23723 vdd.n775 vdd.n766 1.70257
R23724 vdd.n776 vdd.n772 1.70069
R23725 vdd.n771 vdd.n769 1.70069
R23726 vdd.n775 vdd.n774 1.50297
R23727 vdd.n460 vdd.n453 1.5005
R23728 vdd.n946 vdd.n945 1.5005
R23729 vdd.n947 vdd.n692 1.5005
R23730 vdd.n704 vdd.n699 1.5005
R23731 vdd.n1150 vdd.n1149 1.5005
R23732 vdd.n1146 vdd.n951 1.5005
R23733 vdd.n1145 vdd.n952 1.5005
R23734 vdd.n1144 vdd.n953 1.5005
R23735 vdd.n1141 vdd.n957 1.5005
R23736 vdd.n1140 vdd.n958 1.5005
R23737 vdd.n1139 vdd.n959 1.5005
R23738 vdd.n1136 vdd.n963 1.5005
R23739 vdd.n1135 vdd.n964 1.5005
R23740 vdd.n1134 vdd.n965 1.5005
R23741 vdd.n1131 vdd.n969 1.5005
R23742 vdd.n1130 vdd.n970 1.5005
R23743 vdd.n1129 vdd.n971 1.5005
R23744 vdd.n1126 vdd.n975 1.5005
R23745 vdd.n1125 vdd.n976 1.5005
R23746 vdd.n1124 vdd.n977 1.5005
R23747 vdd.n1121 vdd.n981 1.5005
R23748 vdd.n1120 vdd.n982 1.5005
R23749 vdd.n1119 vdd.n1117 1.5005
R23750 vdd.n986 vdd.n598 1.5005
R23751 vdd.n1527 vdd.n1524 1.5005
R23752 vdd.n603 vdd.n594 1.5005
R23753 vdd.n1531 vdd.n596 1.5005
R23754 vdd.n1533 vdd.n1532 1.5005
R23755 vdd.n1541 vdd.n1540 1.5005
R23756 vdd.n590 vdd.n583 1.5005
R23757 vdd.n1548 vdd.n1547 1.5005
R23758 vdd.n1544 vdd.n579 1.5005
R23759 vdd.n1558 vdd.n566 1.5005
R23760 vdd.n1572 vdd.n1571 1.5005
R23761 vdd.n1576 vdd.n1575 1.5005
R23762 vdd.n559 vdd.n553 1.5005
R23763 vdd.n1585 vdd.n1584 1.5005
R23764 vdd.n1589 vdd.n1588 1.5005
R23765 vdd.n546 vdd.n540 1.5005
R23766 vdd.n1598 vdd.n1597 1.5005
R23767 vdd.n1647 vdd.n1646 1.5005
R23768 vdd.n538 vdd.n527 1.5005
R23769 vdd.n1636 vdd.n512 1.5005
R23770 vdd.n1671 vdd.n1670 1.5005
R23771 vdd.n513 vdd.n508 1.5005
R23772 vdd.n1666 vdd.n505 1.5005
R23773 vdd.n1681 vdd.n495 1.5005
R23774 vdd.n1690 vdd.n1689 1.5005
R23775 vdd.n1694 vdd.n1693 1.5005
R23776 vdd.n488 vdd.n482 1.5005
R23777 vdd.n1703 vdd.n1702 1.5005
R23778 vdd.n1707 vdd.n1706 1.5005
R23779 vdd.n475 vdd.n462 1.5005
R23780 vdd.n1726 vdd.n1723 1.5005
R23781 vdd.n467 vdd.n458 1.5005
R23782 vdd.n1792 vdd.n1791 1.5005
R23783 vdd.n2489 vdd.n6 1.5005
R23784 vdd.n2965 vdd.n8 1.5005
R23785 vdd.n2964 vdd.n9 1.5005
R23786 vdd.n2963 vdd.n10 1.5005
R23787 vdd.n2553 vdd.n11 1.5005
R23788 vdd.n2959 vdd.n13 1.5005
R23789 vdd.n2958 vdd.n14 1.5005
R23790 vdd.n2957 vdd.n15 1.5005
R23791 vdd.n2514 vdd.n16 1.5005
R23792 vdd.n2953 vdd.n18 1.5005
R23793 vdd.n2952 vdd.n19 1.5005
R23794 vdd.n2951 vdd.n20 1.5005
R23795 vdd.n2524 vdd.n21 1.5005
R23796 vdd.n2947 vdd.n23 1.5005
R23797 vdd.n2946 vdd.n24 1.5005
R23798 vdd.n2945 vdd.n25 1.5005
R23799 vdd.n221 vdd.n26 1.5005
R23800 vdd.n2941 vdd.n28 1.5005
R23801 vdd.n2940 vdd.n29 1.5005
R23802 vdd.n2939 vdd.n30 1.5005
R23803 vdd.n209 vdd.n31 1.5005
R23804 vdd.n2935 vdd.n33 1.5005
R23805 vdd.n2934 vdd.n34 1.5005
R23806 vdd.n2933 vdd.n35 1.5005
R23807 vdd.n201 vdd.n36 1.5005
R23808 vdd.n2929 vdd.n38 1.5005
R23809 vdd.n2928 vdd.n39 1.5005
R23810 vdd.n2927 vdd.n40 1.5005
R23811 vdd.n186 vdd.n41 1.5005
R23812 vdd.n2923 vdd.n43 1.5005
R23813 vdd.n2922 vdd.n44 1.5005
R23814 vdd.n2921 vdd.n45 1.5005
R23815 vdd.n173 vdd.n46 1.5005
R23816 vdd.n2917 vdd.n48 1.5005
R23817 vdd.n2916 vdd.n49 1.5005
R23818 vdd.n2915 vdd.n50 1.5005
R23819 vdd.n154 vdd.n51 1.5005
R23820 vdd.n2911 vdd.n53 1.5005
R23821 vdd.n2910 vdd.n54 1.5005
R23822 vdd.n2909 vdd.n55 1.5005
R23823 vdd.n2658 vdd.n56 1.5005
R23824 vdd.n2905 vdd.n58 1.5005
R23825 vdd.n2904 vdd.n59 1.5005
R23826 vdd.n2903 vdd.n60 1.5005
R23827 vdd.n2670 vdd.n61 1.5005
R23828 vdd.n2899 vdd.n63 1.5005
R23829 vdd.n2898 vdd.n64 1.5005
R23830 vdd.n2897 vdd.n65 1.5005
R23831 vdd.n2679 vdd.n66 1.5005
R23832 vdd.n2893 vdd.n68 1.5005
R23833 vdd.n2892 vdd.n69 1.5005
R23834 vdd.n2891 vdd.n70 1.5005
R23835 vdd.n2692 vdd.n71 1.5005
R23836 vdd.n2887 vdd.n73 1.5005
R23837 vdd.n2886 vdd.n74 1.5005
R23838 vdd.n2885 vdd.n75 1.5005
R23839 vdd.n2707 vdd.n76 1.5005
R23840 vdd.n2881 vdd.n78 1.5005
R23841 vdd.n2880 vdd.n79 1.5005
R23842 vdd.n2879 vdd.n80 1.5005
R23843 vdd.n2719 vdd.n81 1.5005
R23844 vdd.n2875 vdd.n83 1.5005
R23845 vdd.n2874 vdd.n84 1.5005
R23846 vdd.n2873 vdd.n85 1.5005
R23847 vdd.n128 vdd.n86 1.5005
R23848 vdd.n2869 vdd.n88 1.5005
R23849 vdd.n2868 vdd.n89 1.5005
R23850 vdd.n2867 vdd.n90 1.5005
R23851 vdd.n113 vdd.n91 1.5005
R23852 vdd.n2863 vdd.n93 1.5005
R23853 vdd.n2862 vdd.n94 1.5005
R23854 vdd.n2861 vdd.n95 1.5005
R23855 vdd.n107 vdd.n96 1.5005
R23856 vdd.n2857 vdd.n2856 1.5005
R23857 vdd.n2249 vdd.n2159 1.5005
R23858 vdd.n2248 vdd.n2160 1.5005
R23859 vdd.n2247 vdd.n2161 1.5005
R23860 vdd.n2164 vdd.n2162 1.5005
R23861 vdd.n2243 vdd.n2165 1.5005
R23862 vdd.n2242 vdd.n2166 1.5005
R23863 vdd.n2241 vdd.n2167 1.5005
R23864 vdd.n2170 vdd.n2168 1.5005
R23865 vdd.n2237 vdd.n2171 1.5005
R23866 vdd.n2236 vdd.n2172 1.5005
R23867 vdd.n2235 vdd.n2173 1.5005
R23868 vdd.n2216 vdd.n2174 1.5005
R23869 vdd.n2218 vdd.n2217 1.5005
R23870 vdd.n2219 vdd.n2215 1.5005
R23871 vdd.n2227 vdd.n2220 1.5005
R23872 vdd.n2226 vdd.n2222 1.5005
R23873 vdd.n2221 vdd.n2 1.5005
R23874 vdd.n2971 vdd.n3 1.5005
R23875 vdd.n2970 vdd.n4 1.5005
R23876 vdd.n2969 vdd.n5 1.5005
R23877 vdd.n1905 vdd.n1904 1.5005
R23878 vdd.n345 vdd.n339 1.5005
R23879 vdd.n1909 vdd.n315 1.5005
R23880 vdd.n1910 vdd.n318 1.5005
R23881 vdd.n1912 vdd.n325 1.5005
R23882 vdd.n334 vdd.n329 1.5005
R23883 vdd.n2307 vdd.n2306 1.5005
R23884 vdd.n2303 vdd.n1916 1.5005
R23885 vdd.n2302 vdd.n1917 1.5005
R23886 vdd.n2300 vdd.n1919 1.5005
R23887 vdd.n2047 vdd.n1920 1.5005
R23888 vdd.n2296 vdd.n1922 1.5005
R23889 vdd.n2294 vdd.n1924 1.5005
R23890 vdd.n2293 vdd.n1925 1.5005
R23891 vdd.n2037 vdd.n1926 1.5005
R23892 vdd.n2289 vdd.n1930 1.5005
R23893 vdd.n2288 vdd.n1931 1.5005
R23894 vdd.n2287 vdd.n1932 1.5005
R23895 vdd.n2284 vdd.n1936 1.5005
R23896 vdd.n2283 vdd.n1937 1.5005
R23897 vdd.n2282 vdd.n1938 1.5005
R23898 vdd.n2279 vdd.n1942 1.5005
R23899 vdd.n2278 vdd.n1943 1.5005
R23900 vdd.n2277 vdd.n1944 1.5005
R23901 vdd.n2274 vdd.n1948 1.5005
R23902 vdd.n2273 vdd.n1949 1.5005
R23903 vdd.n2272 vdd.n1950 1.5005
R23904 vdd.n2269 vdd.n1954 1.5005
R23905 vdd.n2268 vdd.n1955 1.5005
R23906 vdd.n2267 vdd.n1956 1.5005
R23907 vdd.n2264 vdd.n1960 1.5005
R23908 vdd.n2263 vdd.n1961 1.5005
R23909 vdd.n2262 vdd.n1962 1.5005
R23910 vdd.n2259 vdd.n1966 1.5005
R23911 vdd.n2258 vdd.n1967 1.5005
R23912 vdd.n2257 vdd.n1968 1.5005
R23913 vdd.n2254 vdd.n1972 1.5005
R23914 vdd.n2253 vdd.n1973 1.5005
R23915 vdd.n2252 vdd.n1974 1.5005
R23916 vdd.n1787 vdd.n450 1.5005
R23917 vdd.n1786 vdd.n447 1.5005
R23918 vdd.n1784 vdd.n444 1.5005
R23919 vdd.n1731 vdd.n441 1.5005
R23920 vdd.n1780 vdd.n438 1.5005
R23921 vdd.n1778 vdd.n435 1.5005
R23922 vdd.n1777 vdd.n428 1.5005
R23923 vdd.n1734 vdd.n431 1.5005
R23924 vdd.n1773 vdd.n422 1.5005
R23925 vdd.n1772 vdd.n419 1.5005
R23926 vdd.n1771 vdd.n416 1.5005
R23927 vdd.n1768 vdd.n413 1.5005
R23928 vdd.n1767 vdd.n410 1.5005
R23929 vdd.n1766 vdd.n407 1.5005
R23930 vdd.n1763 vdd.n400 1.5005
R23931 vdd.n1762 vdd.n405 1.5005
R23932 vdd.n1761 vdd.n394 1.5005
R23933 vdd.n1758 vdd.n391 1.5005
R23934 vdd.n1757 vdd.n388 1.5005
R23935 vdd.n1756 vdd.n385 1.5005
R23936 vdd.n1753 vdd.n382 1.5005
R23937 vdd.n1752 vdd.n378 1.5005
R23938 vdd.n1751 vdd.n371 1.5005
R23939 vdd.n1870 vdd.n1869 1.5005
R23940 vdd.n1871 vdd.n358 1.5005
R23941 vdd.n765 vdd.n757 1.5005
R23942 vdd.n782 vdd.n781 1.5005
R23943 vdd.n803 vdd.n721 1.5005
R23944 vdd.n928 vdd.n722 1.5005
R23945 vdd.n796 vdd.n719 1.5005
R23946 vdd.n934 vdd.n933 1.5005
R23947 vdd.n715 vdd.n708 1.5005
R23948 vdd.n768 vdd.n754 1.5005
R23949 vdd.n777 vdd.n770 1.5005
R23950 vdd.n2212 vdd.n2211 1.49045
R23951 vdd.n2199 vdd.n2176 1.15283
R23952 vdd.n2210 vdd.n2177 1.15283
R23953 vdd.n2231 vdd.n2230 1.15283
R23954 vdd.n2224 vdd.n2223 1.15283
R23955 vdd.n2210 vdd.n2209 1.13717
R23956 vdd.n2184 vdd.n2176 1.13717
R23957 vdd.n779 vdd.n765 1.13717
R23958 vdd.n781 vdd.n780 1.13717
R23959 vdd.n721 vdd.n720 1.13717
R23960 vdd.n929 vdd.n928 1.13717
R23961 vdd.n930 vdd.n719 1.13717
R23962 vdd.n933 vdd.n932 1.13717
R23963 vdd.n931 vdd.n708 1.13717
R23964 vdd.n946 vdd.n707 1.13717
R23965 vdd.n948 vdd.n947 1.13717
R23966 vdd.n949 vdd.n704 1.13717
R23967 vdd.n1149 vdd.n1148 1.13717
R23968 vdd.n1147 vdd.n1146 1.13717
R23969 vdd.n1145 vdd.n950 1.13717
R23970 vdd.n1144 vdd.n1143 1.13717
R23971 vdd.n1142 vdd.n1141 1.13717
R23972 vdd.n1140 vdd.n956 1.13717
R23973 vdd.n1139 vdd.n1138 1.13717
R23974 vdd.n1137 vdd.n1136 1.13717
R23975 vdd.n1135 vdd.n962 1.13717
R23976 vdd.n1134 vdd.n1133 1.13717
R23977 vdd.n1132 vdd.n1131 1.13717
R23978 vdd.n1130 vdd.n968 1.13717
R23979 vdd.n1129 vdd.n1128 1.13717
R23980 vdd.n1127 vdd.n1126 1.13717
R23981 vdd.n1125 vdd.n974 1.13717
R23982 vdd.n1124 vdd.n1123 1.13717
R23983 vdd.n1122 vdd.n1121 1.13717
R23984 vdd.n1120 vdd.n980 1.13717
R23985 vdd.n1119 vdd.n1118 1.13717
R23986 vdd.n598 vdd.n597 1.13717
R23987 vdd.n1528 vdd.n1527 1.13717
R23988 vdd.n1529 vdd.n594 1.13717
R23989 vdd.n1531 vdd.n1530 1.13717
R23990 vdd.n1532 vdd.n586 1.13717
R23991 vdd.n1542 vdd.n1541 1.13717
R23992 vdd.n1543 vdd.n583 1.13717
R23993 vdd.n1547 vdd.n1546 1.13717
R23994 vdd.n1545 vdd.n1544 1.13717
R23995 vdd.n566 vdd.n565 1.13717
R23996 vdd.n1573 vdd.n1572 1.13717
R23997 vdd.n1575 vdd.n1574 1.13717
R23998 vdd.n553 vdd.n552 1.13717
R23999 vdd.n1586 vdd.n1585 1.13717
R24000 vdd.n1588 vdd.n1587 1.13717
R24001 vdd.n540 vdd.n539 1.13717
R24002 vdd.n1599 vdd.n1598 1.13717
R24003 vdd.n1646 vdd.n1645 1.13717
R24004 vdd.n1644 vdd.n538 1.13717
R24005 vdd.n1643 vdd.n1642 1.13717
R24006 vdd.n1601 vdd.n1600 1.13717
R24007 vdd.n1607 vdd.n1606 1.13717
R24008 vdd.n1609 vdd.n1608 1.13717
R24009 vdd.n1611 vdd.n1610 1.13717
R24010 vdd.n1613 vdd.n1612 1.13717
R24011 vdd.n1615 vdd.n1614 1.13717
R24012 vdd.n1616 vdd.n1605 1.13717
R24013 vdd.n1618 vdd.n1617 1.13717
R24014 vdd.n518 vdd.n514 1.13717
R24015 vdd.n1662 vdd.n1661 1.13717
R24016 vdd.n1663 vdd.n512 1.13717
R24017 vdd.n1670 vdd.n1669 1.13717
R24018 vdd.n1668 vdd.n513 1.13717
R24019 vdd.n1667 vdd.n1666 1.13717
R24020 vdd.n495 vdd.n494 1.13717
R24021 vdd.n1691 vdd.n1690 1.13717
R24022 vdd.n1693 vdd.n1692 1.13717
R24023 vdd.n482 vdd.n481 1.13717
R24024 vdd.n1704 vdd.n1703 1.13717
R24025 vdd.n1706 vdd.n1705 1.13717
R24026 vdd.n462 vdd.n461 1.13717
R24027 vdd.n1727 vdd.n1726 1.13717
R24028 vdd.n1728 vdd.n458 1.13717
R24029 vdd.n1791 vdd.n1790 1.13717
R24030 vdd.n1789 vdd.n460 1.13717
R24031 vdd.n1788 vdd.n1787 1.13717
R24032 vdd.n1786 vdd.n1729 1.13717
R24033 vdd.n1784 vdd.n1783 1.13717
R24034 vdd.n1782 vdd.n1731 1.13717
R24035 vdd.n1781 vdd.n1780 1.13717
R24036 vdd.n1778 vdd.n1732 1.13717
R24037 vdd.n1777 vdd.n1776 1.13717
R24038 vdd.n1775 vdd.n1734 1.13717
R24039 vdd.n1774 vdd.n1773 1.13717
R24040 vdd.n1772 vdd.n1735 1.13717
R24041 vdd.n1771 vdd.n1770 1.13717
R24042 vdd.n1769 vdd.n1768 1.13717
R24043 vdd.n1767 vdd.n1740 1.13717
R24044 vdd.n1766 vdd.n1765 1.13717
R24045 vdd.n1764 vdd.n1763 1.13717
R24046 vdd.n1762 vdd.n1743 1.13717
R24047 vdd.n1761 vdd.n1760 1.13717
R24048 vdd.n1759 vdd.n1758 1.13717
R24049 vdd.n1757 vdd.n1746 1.13717
R24050 vdd.n1756 vdd.n1755 1.13717
R24051 vdd.n1754 vdd.n1753 1.13717
R24052 vdd.n1752 vdd.n1749 1.13717
R24053 vdd.n1751 vdd.n1750 1.13717
R24054 vdd.n1870 vdd.n369 1.13717
R24055 vdd.n1872 vdd.n1871 1.13717
R24056 vdd.n1873 vdd.n364 1.13717
R24057 vdd.n1893 vdd.n1892 1.13717
R24058 vdd.n1891 vdd.n1890 1.13717
R24059 vdd.n1889 vdd.n1888 1.13717
R24060 vdd.n1875 vdd.n1874 1.13717
R24061 vdd.n1879 vdd.n1878 1.13717
R24062 vdd.n1881 vdd.n1880 1.13717
R24063 vdd.n1882 vdd.n1877 1.13717
R24064 vdd.n1884 vdd.n1883 1.13717
R24065 vdd.n341 vdd.n340 1.13717
R24066 vdd.n1906 vdd.n1905 1.13717
R24067 vdd.n1907 vdd.n339 1.13717
R24068 vdd.n1909 vdd.n1908 1.13717
R24069 vdd.n1910 vdd.n337 1.13717
R24070 vdd.n1913 vdd.n1912 1.13717
R24071 vdd.n1914 vdd.n334 1.13717
R24072 vdd.n2306 vdd.n2305 1.13717
R24073 vdd.n2304 vdd.n2303 1.13717
R24074 vdd.n2302 vdd.n1915 1.13717
R24075 vdd.n2300 vdd.n2299 1.13717
R24076 vdd.n2298 vdd.n1920 1.13717
R24077 vdd.n2297 vdd.n2296 1.13717
R24078 vdd.n2294 vdd.n1921 1.13717
R24079 vdd.n2293 vdd.n2292 1.13717
R24080 vdd.n2291 vdd.n1926 1.13717
R24081 vdd.n2290 vdd.n2289 1.13717
R24082 vdd.n2288 vdd.n1927 1.13717
R24083 vdd.n2287 vdd.n2286 1.13717
R24084 vdd.n2285 vdd.n2284 1.13717
R24085 vdd.n2283 vdd.n1935 1.13717
R24086 vdd.n2282 vdd.n2281 1.13717
R24087 vdd.n2280 vdd.n2279 1.13717
R24088 vdd.n2278 vdd.n1941 1.13717
R24089 vdd.n2277 vdd.n2276 1.13717
R24090 vdd.n2275 vdd.n2274 1.13717
R24091 vdd.n2273 vdd.n1947 1.13717
R24092 vdd.n2272 vdd.n2271 1.13717
R24093 vdd.n2270 vdd.n2269 1.13717
R24094 vdd.n2268 vdd.n1953 1.13717
R24095 vdd.n2267 vdd.n2266 1.13717
R24096 vdd.n2265 vdd.n2264 1.13717
R24097 vdd.n2263 vdd.n1959 1.13717
R24098 vdd.n2262 vdd.n2261 1.13717
R24099 vdd.n2260 vdd.n2259 1.13717
R24100 vdd.n2258 vdd.n1965 1.13717
R24101 vdd.n2257 vdd.n2256 1.13717
R24102 vdd.n2255 vdd.n2254 1.13717
R24103 vdd.n2253 vdd.n1971 1.13717
R24104 vdd.n2252 vdd.n2251 1.13717
R24105 vdd.n2250 vdd.n2249 1.13717
R24106 vdd.n2248 vdd.n1976 1.13717
R24107 vdd.n2247 vdd.n2246 1.13717
R24108 vdd.n2245 vdd.n2162 1.13717
R24109 vdd.n2244 vdd.n2243 1.13717
R24110 vdd.n2242 vdd.n2163 1.13717
R24111 vdd.n2241 vdd.n2240 1.13717
R24112 vdd.n2239 vdd.n2168 1.13717
R24113 vdd.n2238 vdd.n2237 1.13717
R24114 vdd.n2236 vdd.n2169 1.13717
R24115 vdd.n2235 vdd.n2234 1.13717
R24116 vdd.n2233 vdd.n2174 1.13717
R24117 vdd.n2217 vdd.n2175 1.13717
R24118 vdd.n2215 vdd.n2213 1.13717
R24119 vdd.n2228 vdd.n2227 1.13717
R24120 vdd.n2230 vdd.n2229 1.13717
R24121 vdd.n2223 vdd.n2214 1.13717
R24122 vdd.n2226 vdd.n2225 1.13717
R24123 vdd.n2 vdd.n0 1.13717
R24124 vdd.n2972 vdd.n2971 1.13717
R24125 vdd.n2970 vdd.n1 1.13717
R24126 vdd.n2969 vdd.n2968 1.13717
R24127 vdd.n2967 vdd.n6 1.13717
R24128 vdd.n2966 vdd.n2965 1.13717
R24129 vdd.n2964 vdd.n7 1.13717
R24130 vdd.n2963 vdd.n2962 1.13717
R24131 vdd.n2961 vdd.n11 1.13717
R24132 vdd.n2960 vdd.n2959 1.13717
R24133 vdd.n2958 vdd.n12 1.13717
R24134 vdd.n2957 vdd.n2956 1.13717
R24135 vdd.n2955 vdd.n16 1.13717
R24136 vdd.n2954 vdd.n2953 1.13717
R24137 vdd.n2952 vdd.n17 1.13717
R24138 vdd.n2951 vdd.n2950 1.13717
R24139 vdd.n2949 vdd.n21 1.13717
R24140 vdd.n2948 vdd.n2947 1.13717
R24141 vdd.n2946 vdd.n22 1.13717
R24142 vdd.n2945 vdd.n2944 1.13717
R24143 vdd.n2943 vdd.n26 1.13717
R24144 vdd.n2942 vdd.n2941 1.13717
R24145 vdd.n2940 vdd.n27 1.13717
R24146 vdd.n2939 vdd.n2938 1.13717
R24147 vdd.n2937 vdd.n31 1.13717
R24148 vdd.n2936 vdd.n2935 1.13717
R24149 vdd.n2934 vdd.n32 1.13717
R24150 vdd.n2933 vdd.n2932 1.13717
R24151 vdd.n2931 vdd.n36 1.13717
R24152 vdd.n2930 vdd.n2929 1.13717
R24153 vdd.n2928 vdd.n37 1.13717
R24154 vdd.n2927 vdd.n2926 1.13717
R24155 vdd.n2925 vdd.n41 1.13717
R24156 vdd.n2924 vdd.n2923 1.13717
R24157 vdd.n2922 vdd.n42 1.13717
R24158 vdd.n2921 vdd.n2920 1.13717
R24159 vdd.n2919 vdd.n46 1.13717
R24160 vdd.n2918 vdd.n2917 1.13717
R24161 vdd.n2916 vdd.n47 1.13717
R24162 vdd.n2915 vdd.n2914 1.13717
R24163 vdd.n2913 vdd.n51 1.13717
R24164 vdd.n2912 vdd.n2911 1.13717
R24165 vdd.n2910 vdd.n52 1.13717
R24166 vdd.n2909 vdd.n2908 1.13717
R24167 vdd.n2907 vdd.n56 1.13717
R24168 vdd.n2906 vdd.n2905 1.13717
R24169 vdd.n2904 vdd.n57 1.13717
R24170 vdd.n2903 vdd.n2902 1.13717
R24171 vdd.n2901 vdd.n61 1.13717
R24172 vdd.n2900 vdd.n2899 1.13717
R24173 vdd.n2898 vdd.n62 1.13717
R24174 vdd.n2897 vdd.n2896 1.13717
R24175 vdd.n2895 vdd.n66 1.13717
R24176 vdd.n2894 vdd.n2893 1.13717
R24177 vdd.n2892 vdd.n67 1.13717
R24178 vdd.n2891 vdd.n2890 1.13717
R24179 vdd.n2889 vdd.n71 1.13717
R24180 vdd.n2888 vdd.n2887 1.13717
R24181 vdd.n2886 vdd.n72 1.13717
R24182 vdd.n2885 vdd.n2884 1.13717
R24183 vdd.n2883 vdd.n76 1.13717
R24184 vdd.n2882 vdd.n2881 1.13717
R24185 vdd.n2880 vdd.n77 1.13717
R24186 vdd.n2879 vdd.n2878 1.13717
R24187 vdd.n2877 vdd.n81 1.13717
R24188 vdd.n2876 vdd.n2875 1.13717
R24189 vdd.n2874 vdd.n82 1.13717
R24190 vdd.n2873 vdd.n2872 1.13717
R24191 vdd.n2871 vdd.n86 1.13717
R24192 vdd.n2870 vdd.n2869 1.13717
R24193 vdd.n2868 vdd.n87 1.13717
R24194 vdd.n2867 vdd.n2866 1.13717
R24195 vdd.n2865 vdd.n91 1.13717
R24196 vdd.n2864 vdd.n2863 1.13717
R24197 vdd.n2862 vdd.n92 1.13717
R24198 vdd.n2861 vdd.n2860 1.13717
R24199 vdd.n2859 vdd.n96 1.13717
R24200 vdd.n1428 vdd.n1335 1.12991
R24201 vdd.n2330 vdd.n2329 0.753441
R24202 vdd.n926 vdd.n925 0.643357
R24203 vdd.n725 vdd.n723 0.643357
R24204 vdd.n734 vdd.n732 0.643357
R24205 vdd.n916 vdd.n915 0.643357
R24206 vdd.n914 vdd.n913 0.643357
R24207 vdd.n736 vdd.n735 0.643357
R24208 vdd.n748 vdd.n746 0.643357
R24209 vdd.n904 vdd.n903 0.643357
R24210 vdd.n902 vdd.n901 0.643357
R24211 vdd.n823 vdd.n822 0.643357
R24212 vdd.n824 vdd.n819 0.643357
R24213 vdd.n889 vdd.n888 0.643357
R24214 vdd.n891 vdd.n890 0.643357
R24215 vdd.n826 vdd.n825 0.643357
R24216 vdd.n836 vdd.n834 0.643357
R24217 vdd.n879 vdd.n878 0.643357
R24218 vdd.n877 vdd.n876 0.643357
R24219 vdd.n838 vdd.n837 0.643357
R24220 vdd.n728 vdd.n726 0.563
R24221 vdd.n922 vdd.n921 0.563
R24222 vdd.n920 vdd.n919 0.563
R24223 vdd.n730 vdd.n729 0.563
R24224 vdd.n740 vdd.n738 0.563
R24225 vdd.n910 vdd.n909 0.563
R24226 vdd.n908 vdd.n907 0.563
R24227 vdd.n743 vdd.n741 0.563
R24228 vdd.n753 vdd.n752 0.563
R24229 vdd.n897 vdd.n896 0.563
R24230 vdd.n895 vdd.n894 0.563
R24231 vdd.n830 vdd.n828 0.563
R24232 vdd.n818 vdd.n817 0.563
R24233 vdd.n885 vdd.n884 0.563
R24234 vdd.n883 vdd.n882 0.563
R24235 vdd.n832 vdd.n831 0.563
R24236 vdd.n842 vdd.n840 0.563
R24237 vdd.n873 vdd.n872 0.563
R24238 vdd.n2181 vdd.n2179 0.45282
R24239 vdd.n2181 vdd.n2180 0.447611
R24240 vdd.n1659 vdd.n524 0.254416
R24241 vdd.n2343 vdd.n297 0.250952
R24242 vdd.n2858 vdd.n97 0.230231
R24243 vdd.n2859 vdd.n2858 0.136149
R24244 vdd.n2204 vdd.n2202 0.111491
R24245 vdd.n2182 vdd.n2181 0.106269
R24246 vdd.n2858 vdd.n2857 0.0908604
R24247 vdd.n2232 vdd 0.081944
R24248 vdd.n1501 vdd.n1296 0.063569
R24249 vdd.n1499 vdd.n1498 0.063569
R24250 vdd.n1497 vdd.n1496 0.063569
R24251 vdd.n1495 vdd.n1494 0.063569
R24252 vdd.n2340 vdd.n298 0.063569
R24253 vdd.n2334 vdd.n299 0.063569
R24254 vdd.n2335 vdd.n300 0.063569
R24255 vdd.n2336 vdd.n301 0.063569
R24256 vdd.n2337 vdd.n302 0.063569
R24257 vdd.n2337 vdd.n301 0.063569
R24258 vdd.n2336 vdd.n300 0.063569
R24259 vdd.n2335 vdd.n299 0.063569
R24260 vdd.n2334 vdd.n298 0.063569
R24261 vdd.n1494 vdd.n1493 0.063569
R24262 vdd.n1496 vdd.n1495 0.063569
R24263 vdd.n1498 vdd.n1497 0.063569
R24264 vdd.n1499 vdd.n1296 0.063569
R24265 vdd.n1168 vdd.n1167 0.063
R24266 vdd.n1168 vdd.n683 0.063
R24267 vdd.n1175 vdd.n683 0.063
R24268 vdd.n1177 vdd.n678 0.063
R24269 vdd.n1184 vdd.n678 0.063
R24270 vdd.n1186 vdd.n673 0.063
R24271 vdd.n1195 vdd.n673 0.063
R24272 vdd.n1197 vdd.n668 0.063
R24273 vdd.n1204 vdd.n668 0.063
R24274 vdd.n1206 vdd.n663 0.063
R24275 vdd.n1213 vdd.n663 0.063
R24276 vdd.n1215 vdd.n658 0.063
R24277 vdd.n1224 vdd.n658 0.063
R24278 vdd.n1226 vdd.n653 0.063
R24279 vdd.n1234 vdd.n653 0.063
R24280 vdd.n1236 vdd.n648 0.063
R24281 vdd.n1243 vdd.n648 0.063
R24282 vdd.n1245 vdd.n643 0.063
R24283 vdd.n1254 vdd.n643 0.063
R24284 vdd.n1256 vdd.n638 0.063
R24285 vdd.n1263 vdd.n638 0.063
R24286 vdd.n1265 vdd.n1263 0.063
R24287 vdd.n1265 vdd.n1264 0.063
R24288 vdd.n1274 vdd.n1273 0.063
R24289 vdd.n1275 vdd.n1274 0.063
R24290 vdd.n1285 vdd.n1283 0.063
R24291 vdd.n1285 vdd.n1284 0.063
R24292 vdd.n1294 vdd.n1293 0.063
R24293 vdd.n1503 vdd.n1294 0.063
R24294 vdd.n1503 vdd.n1502 0.063
R24295 vdd.n1492 vdd.n1491 0.063
R24296 vdd.n1491 vdd.n1298 0.063
R24297 vdd.n1483 vdd.n1298 0.063
R24298 vdd.n1481 vdd.n1306 0.063
R24299 vdd.n1474 vdd.n1306 0.063
R24300 vdd.n1472 vdd.n1312 0.063
R24301 vdd.n1465 vdd.n1312 0.063
R24302 vdd.n1463 vdd.n1317 0.063
R24303 vdd.n1455 vdd.n1317 0.063
R24304 vdd.n1453 vdd.n1322 0.063
R24305 vdd.n1446 vdd.n1322 0.063
R24306 vdd.n1444 vdd.n1328 0.063
R24307 vdd.n1437 vdd.n1328 0.063
R24308 vdd.n1435 vdd.n1333 0.063
R24309 vdd.n1340 vdd.n1333 0.063
R24310 vdd.n1424 vdd.n1423 0.063
R24311 vdd.n1423 vdd.n1342 0.063
R24312 vdd.n1416 vdd.n1415 0.063
R24313 vdd.n1415 vdd.n1348 0.063
R24314 vdd.n1408 vdd.n1407 0.063
R24315 vdd.n1407 vdd.n1354 0.063
R24316 vdd.n1399 vdd.n1398 0.063
R24317 vdd.n1398 vdd.n1361 0.063
R24318 vdd.n1391 vdd.n1390 0.063
R24319 vdd.n1390 vdd.n1367 0.063
R24320 vdd.n1383 vdd.n1382 0.063
R24321 vdd.n1382 vdd.n1374 0.063
R24322 vdd.n2333 vdd.n304 0.063
R24323 vdd.n2341 vdd.n2333 0.063
R24324 vdd.n2338 vdd.n292 0.063
R24325 vdd.n2350 vdd.n292 0.063
R24326 vdd.n2353 vdd.n2350 0.063
R24327 vdd.n2362 vdd.n288 0.063
R24328 vdd.n2365 vdd.n2362 0.063
R24329 vdd.n2372 vdd.n284 0.063
R24330 vdd.n2375 vdd.n2372 0.063
R24331 vdd.n2382 vdd.n280 0.063
R24332 vdd.n2385 vdd.n2382 0.063
R24333 vdd.n2394 vdd.n276 0.063
R24334 vdd.n2397 vdd.n2394 0.063
R24335 vdd.n2404 vdd.n272 0.063
R24336 vdd.n2407 vdd.n2404 0.063
R24337 vdd.n2415 vdd.n268 0.063
R24338 vdd.n2418 vdd.n2415 0.063
R24339 vdd.n2427 vdd.n264 0.063
R24340 vdd.n2430 vdd.n2427 0.063
R24341 vdd.n2437 vdd.n260 0.063
R24342 vdd.n2440 vdd.n2437 0.063
R24343 vdd.n2447 vdd.n256 0.063
R24344 vdd.n2450 vdd.n2447 0.063
R24345 vdd.n2459 vdd.n252 0.063
R24346 vdd.n2462 vdd.n2459 0.063
R24347 vdd.n2469 vdd.n248 0.063
R24348 vdd.n2471 vdd.n243 0.063
R24349 vdd.n2478 vdd.n243 0.063
R24350 vdd.n1483 vdd.n1482 0.0622188
R24351 vdd.n767 vdd.n728 0.0615656
R24352 vdd.n2461 vdd.n248 0.0614375
R24353 vdd.n2470 vdd.n2469 0.0614375
R24354 vdd.n1256 vdd.n1255 0.059875
R24355 vdd.n1264 vdd.n633 0.059875
R24356 vdd.n1474 vdd.n1473 0.0590938
R24357 vdd.n2449 vdd.n252 0.0583125
R24358 vdd.n2479 vdd.n2478 0.0583125
R24359 vdd.n2971 vdd.n2 0.0582617
R24360 vdd.n2221 vdd.n3 0.0582617
R24361 vdd.n1193 vdd.n674 0.05675
R24362 vdd.n1222 vdd.n659 0.05675
R24363 vdd.n1252 vdd.n644 0.05675
R24364 vdd.n1281 vdd.n629 0.05675
R24365 vdd.n1486 vdd.n1485 0.05675
R24366 vdd.n1458 vdd.n1457 0.05675
R24367 vdd.n1430 vdd.n1429 0.05675
R24368 vdd.n1405 vdd.n1355 0.05675
R24369 vdd.n1380 vdd.n1377 0.05675
R24370 vdd.n2360 vdd.n289 0.05675
R24371 vdd.n2392 vdd.n277 0.05675
R24372 vdd.n2425 vdd.n265 0.05675
R24373 vdd.n2457 vdd.n253 0.05675
R24374 vdd.n1245 vdd.n1244 0.05675
R24375 vdd.n1275 vdd.n628 0.05675
R24376 vdd.n1166 vdd.n686 0.0559687
R24377 vdd.n1194 vdd.n671 0.0559687
R24378 vdd.n1223 vdd.n656 0.0559687
R24379 vdd.n1253 vdd.n641 0.0559687
R24380 vdd.n1282 vdd.n626 0.0559687
R24381 vdd.n1484 vdd.n1304 0.0559687
R24382 vdd.n1456 vdd.n1320 0.0559687
R24383 vdd.n1426 vdd.n1336 0.0559687
R24384 vdd.n1401 vdd.n1357 0.0559687
R24385 vdd.n1376 vdd.n1375 0.0559687
R24386 vdd.n2361 vdd.n287 0.0559687
R24387 vdd.n2393 vdd.n275 0.0559687
R24388 vdd.n2426 vdd.n263 0.0559687
R24389 vdd.n2458 vdd.n251 0.0559687
R24390 vdd.n1465 vdd.n1464 0.0559687
R24391 vdd.n2439 vdd.n256 0.0551875
R24392 vdd.n1236 vdd.n1235 0.053625
R24393 vdd.n1284 vdd.n623 0.053625
R24394 vdd.n1455 vdd.n1454 0.0528437
R24395 vdd.n1167 vdd.n687 0.0522857
R24396 vdd.n2429 vdd.n260 0.0520625
R24397 vdd.n1189 vdd.n1188 0.0512812
R24398 vdd.n1218 vdd.n1217 0.0512812
R24399 vdd.n1248 vdd.n1247 0.0512812
R24400 vdd.n1277 vdd.n1276 0.0512812
R24401 vdd.n1489 vdd.n1299 0.0512812
R24402 vdd.n1461 vdd.n1318 0.0512812
R24403 vdd.n1433 vdd.n1334 0.0512812
R24404 vdd.n1406 vdd.n1351 0.0512812
R24405 vdd.n1381 vdd.n1370 0.0512812
R24406 vdd.n2356 vdd.n2355 0.0512812
R24407 vdd.n2388 vdd.n2387 0.0512812
R24408 vdd.n2421 vdd.n2420 0.0512812
R24409 vdd.n2453 vdd.n2452 0.0512812
R24410 vdd.n1226 vdd.n1225 0.0505
R24411 vdd.n1170 vdd.n1169 0.0497188
R24412 vdd.n1199 vdd.n1198 0.0497188
R24413 vdd.n1228 vdd.n1227 0.0497188
R24414 vdd.n1258 vdd.n1257 0.0497188
R24415 vdd.n1287 vdd.n1286 0.0497188
R24416 vdd.n1480 vdd.n1479 0.0497188
R24417 vdd.n1452 vdd.n1451 0.0497188
R24418 vdd.n1425 vdd.n1338 0.0497188
R24419 vdd.n1400 vdd.n1358 0.0497188
R24420 vdd.n2331 vdd.n305 0.0497188
R24421 vdd.n2367 vdd.n2366 0.0497188
R24422 vdd.n2399 vdd.n2398 0.0497188
R24423 vdd.n2432 vdd.n2431 0.0497188
R24424 vdd.n2464 vdd.n2463 0.0497188
R24425 vdd.n1446 vdd.n1445 0.0497188
R24426 vdd.n2417 vdd.n264 0.0489375
R24427 vdd.n1165 vdd.n688 0.0475982
R24428 vdd.n1215 vdd.n1214 0.047375
R24429 vdd.n1437 vdd.n1436 0.0465938
R24430 vdd.n872 vdd.n871 0.0461565
R24431 vdd.n2406 vdd.n268 0.0458125
R24432 vdd.n871 vdd.n843 0.0451429
R24433 vdd.n864 vdd.n843 0.0451429
R24434 vdd.n864 vdd.n863 0.0451429
R24435 vdd.n854 vdd.n853 0.0451429
R24436 vdd.n854 vdd.n687 0.0451429
R24437 vdd.n1187 vdd.n676 0.0450312
R24438 vdd.n1216 vdd.n661 0.0450312
R24439 vdd.n1246 vdd.n646 0.0450312
R24440 vdd.n1271 vdd.n631 0.0450312
R24441 vdd.n1462 vdd.n1315 0.0450312
R24442 vdd.n1434 vdd.n1331 0.0450312
R24443 vdd.n1410 vdd.n1409 0.0450312
R24444 vdd.n1385 vdd.n1384 0.0450312
R24445 vdd.n2354 vdd.n291 0.0450312
R24446 vdd.n2386 vdd.n279 0.0450312
R24447 vdd.n2419 vdd.n267 0.0450312
R24448 vdd.n2451 vdd.n255 0.0450312
R24449 vdd.n2480 vdd.n242 0.0450312
R24450 vdd.n1206 vdd.n1205 0.04425
R24451 vdd.n1173 vdd.n684 0.0434688
R24452 vdd.n1202 vdd.n669 0.0434688
R24453 vdd.n1232 vdd.n654 0.0434688
R24454 vdd.n1261 vdd.n639 0.0434688
R24455 vdd.n1290 vdd.n624 0.0434688
R24456 vdd.n1476 vdd.n1307 0.0434688
R24457 vdd.n1448 vdd.n1323 0.0434688
R24458 vdd.n1422 vdd.n1421 0.0434688
R24459 vdd.n1397 vdd.n1396 0.0434688
R24460 vdd.n2332 vdd.n296 0.0434688
R24461 vdd.n2370 vdd.n285 0.0434688
R24462 vdd.n2402 vdd.n273 0.0434688
R24463 vdd.n2435 vdd.n261 0.0434688
R24464 vdd.n2467 vdd.n249 0.0434688
R24465 vdd.n1341 vdd.n1340 0.0434688
R24466 vdd.n2396 vdd.n272 0.0426875
R24467 vdd.n1197 vdd.n1196 0.041125
R24468 vdd.n1347 vdd.n1342 0.0403437
R24469 vdd.n2384 vdd.n276 0.0395625
R24470 vdd.n2203 vdd.n2197 0.0394423
R24471 vdd.n853 vdd.n848 0.0390045
R24472 vdd.n1183 vdd.n1182 0.0387813
R24473 vdd.n1212 vdd.n1211 0.0387813
R24474 vdd.n1242 vdd.n1241 0.0387813
R24475 vdd.n1272 vdd.n1270 0.0387813
R24476 vdd.n1467 vdd.n1466 0.0387813
R24477 vdd.n1439 vdd.n1438 0.0387813
R24478 vdd.n1413 vdd.n1349 0.0387813
R24479 vdd.n1388 vdd.n1368 0.0387813
R24480 vdd.n2349 vdd.n2348 0.0387813
R24481 vdd.n2381 vdd.n2380 0.0387813
R24482 vdd.n2414 vdd.n2413 0.0387813
R24483 vdd.n2446 vdd.n2445 0.0387813
R24484 vdd.n2477 vdd.n2476 0.0387813
R24485 vdd.n1373 vdd.n304 0.0387813
R24486 vdd.n1186 vdd.n1185 0.038
R24487 vdd.n813 vdd.n755 0.0379794
R24488 vdd.n1136 vdd.n1135 0.0375036
R24489 vdd.n1125 vdd.n1124 0.0375036
R24490 vdd.n1531 vdd.n594 0.0375036
R24491 vdd.n1572 vdd.n566 0.0375036
R24492 vdd.n1670 vdd.n512 0.0375036
R24493 vdd.n1703 vdd.n482 0.0375036
R24494 vdd.n1787 vdd.n460 0.0375036
R24495 vdd.n1777 vdd.n1734 0.0375036
R24496 vdd.n1753 vdd.n1752 0.0375036
R24497 vdd.n1905 vdd.n341 0.0375036
R24498 vdd.n2293 vdd.n1926 0.0375036
R24499 vdd.n2269 vdd.n2268 0.0375036
R24500 vdd.n2258 vdd.n2257 0.0375036
R24501 vdd.n2247 vdd.n2162 0.0375036
R24502 vdd.n2236 vdd.n2235 0.0375036
R24503 vdd.n2963 vdd.n11 0.0375036
R24504 vdd.n2952 vdd.n2951 0.0375036
R24505 vdd.n2941 vdd.n2940 0.0375036
R24506 vdd.n2929 vdd.n36 0.0375036
R24507 vdd.n2921 vdd.n46 0.0375036
R24508 vdd.n2910 vdd.n2909 0.0375036
R24509 vdd.n2899 vdd.n2898 0.0375036
R24510 vdd.n2887 vdd.n71 0.0375036
R24511 vdd.n2879 vdd.n81 0.0375036
R24512 vdd.n2868 vdd.n2867 0.0375036
R24513 vdd.n2164 vdd.n2161 0.0375036
R24514 vdd.n2173 vdd.n2172 0.0375036
R24515 vdd.n1174 vdd.n681 0.0372187
R24516 vdd.n1203 vdd.n666 0.0372187
R24517 vdd.n1233 vdd.n651 0.0372187
R24518 vdd.n1262 vdd.n636 0.0372187
R24519 vdd.n1292 vdd.n1291 0.0372187
R24520 vdd.n1475 vdd.n1310 0.0372187
R24521 vdd.n1447 vdd.n1326 0.0372187
R24522 vdd.n1418 vdd.n1343 0.0372187
R24523 vdd.n1393 vdd.n1362 0.0372187
R24524 vdd.n2371 vdd.n283 0.0372187
R24525 vdd.n2403 vdd.n271 0.0372187
R24526 vdd.n2436 vdd.n259 0.0372187
R24527 vdd.n2468 vdd.n246 0.0372187
R24528 vdd.n1353 vdd.n1348 0.0372187
R24529 vdd.n947 vdd.n946 0.0370523
R24530 vdd.n947 vdd.n704 0.0370523
R24531 vdd.n1149 vdd.n704 0.0370523
R24532 vdd.n1146 vdd.n1145 0.0370523
R24533 vdd.n1145 vdd.n1144 0.0370523
R24534 vdd.n1141 vdd.n1140 0.0370523
R24535 vdd.n1140 vdd.n1139 0.0370523
R24536 vdd.n1135 vdd.n1134 0.0370523
R24537 vdd.n1131 vdd.n1130 0.0370523
R24538 vdd.n1130 vdd.n1129 0.0370523
R24539 vdd.n1126 vdd.n1125 0.0370523
R24540 vdd.n1121 vdd.n1120 0.0370523
R24541 vdd.n1120 vdd.n1119 0.0370523
R24542 vdd.n1119 vdd.n598 0.0370523
R24543 vdd.n1527 vdd.n598 0.0370523
R24544 vdd.n1532 vdd.n1531 0.0370523
R24545 vdd.n1541 vdd.n583 0.0370523
R24546 vdd.n1547 vdd.n583 0.0370523
R24547 vdd.n1544 vdd.n566 0.0370523
R24548 vdd.n1575 vdd.n553 0.0370523
R24549 vdd.n1585 vdd.n553 0.0370523
R24550 vdd.n1588 vdd.n540 0.0370523
R24551 vdd.n1598 vdd.n540 0.0370523
R24552 vdd.n1646 vdd.n538 0.0370523
R24553 vdd.n1642 vdd.n538 0.0370523
R24554 vdd.n1661 vdd.n512 0.0370523
R24555 vdd.n1670 vdd.n513 0.0370523
R24556 vdd.n1666 vdd.n495 0.0370523
R24557 vdd.n1690 vdd.n495 0.0370523
R24558 vdd.n1693 vdd.n482 0.0370523
R24559 vdd.n1706 vdd.n462 0.0370523
R24560 vdd.n1726 vdd.n462 0.0370523
R24561 vdd.n1791 vdd.n458 0.0370523
R24562 vdd.n1791 vdd.n460 0.0370523
R24563 vdd.n1787 vdd.n1786 0.0370523
R24564 vdd.n1784 vdd.n1731 0.0370523
R24565 vdd.n1780 vdd.n1731 0.0370523
R24566 vdd.n1778 vdd.n1777 0.0370523
R24567 vdd.n1773 vdd.n1772 0.0370523
R24568 vdd.n1772 vdd.n1771 0.0370523
R24569 vdd.n1768 vdd.n1767 0.0370523
R24570 vdd.n1767 vdd.n1766 0.0370523
R24571 vdd.n1763 vdd.n1762 0.0370523
R24572 vdd.n1762 vdd.n1761 0.0370523
R24573 vdd.n1758 vdd.n1757 0.0370523
R24574 vdd.n1757 vdd.n1756 0.0370523
R24575 vdd.n1752 vdd.n1751 0.0370523
R24576 vdd.n1871 vdd.n1870 0.0370523
R24577 vdd.n1871 vdd.n364 0.0370523
R24578 vdd.n1905 vdd.n339 0.0370523
R24579 vdd.n1909 vdd.n339 0.0370523
R24580 vdd.n1910 vdd.n1909 0.0370523
R24581 vdd.n1912 vdd.n334 0.0370523
R24582 vdd.n2306 vdd.n334 0.0370523
R24583 vdd.n2303 vdd.n2302 0.0370523
R24584 vdd.n2300 vdd.n1920 0.0370523
R24585 vdd.n2296 vdd.n1920 0.0370523
R24586 vdd.n2294 vdd.n2293 0.0370523
R24587 vdd.n2289 vdd.n2288 0.0370523
R24588 vdd.n2288 vdd.n2287 0.0370523
R24589 vdd.n2284 vdd.n2283 0.0370523
R24590 vdd.n2283 vdd.n2282 0.0370523
R24591 vdd.n2279 vdd.n2278 0.0370523
R24592 vdd.n2278 vdd.n2277 0.0370523
R24593 vdd.n2274 vdd.n2273 0.0370523
R24594 vdd.n2273 vdd.n2272 0.0370523
R24595 vdd.n2268 vdd.n2267 0.0370523
R24596 vdd.n2264 vdd.n2263 0.0370523
R24597 vdd.n2263 vdd.n2262 0.0370523
R24598 vdd.n2259 vdd.n2258 0.0370523
R24599 vdd.n2254 vdd.n2253 0.0370523
R24600 vdd.n2253 vdd.n2252 0.0370523
R24601 vdd.n2249 vdd.n2248 0.0370523
R24602 vdd.n2248 vdd.n2247 0.0370523
R24603 vdd.n2243 vdd.n2162 0.0370523
R24604 vdd.n2243 vdd.n2242 0.0370523
R24605 vdd.n2242 vdd.n2241 0.0370523
R24606 vdd.n2241 vdd.n2168 0.0370523
R24607 vdd.n2237 vdd.n2168 0.0370523
R24608 vdd.n2237 vdd.n2236 0.0370523
R24609 vdd.n2235 vdd.n2174 0.0370523
R24610 vdd.n2217 vdd.n2174 0.0370523
R24611 vdd.n2217 vdd.n2215 0.0370523
R24612 vdd.n2227 vdd.n2215 0.0370523
R24613 vdd.n2227 vdd.n2226 0.0370523
R24614 vdd.n2226 vdd.n2 0.0370523
R24615 vdd.n2971 vdd.n2970 0.0370523
R24616 vdd.n2970 vdd.n2969 0.0370523
R24617 vdd.n2969 vdd.n6 0.0370523
R24618 vdd.n2965 vdd.n6 0.0370523
R24619 vdd.n2965 vdd.n2964 0.0370523
R24620 vdd.n2964 vdd.n2963 0.0370523
R24621 vdd.n2959 vdd.n11 0.0370523
R24622 vdd.n2959 vdd.n2958 0.0370523
R24623 vdd.n2958 vdd.n2957 0.0370523
R24624 vdd.n2957 vdd.n16 0.0370523
R24625 vdd.n2953 vdd.n16 0.0370523
R24626 vdd.n2953 vdd.n2952 0.0370523
R24627 vdd.n2951 vdd.n21 0.0370523
R24628 vdd.n2947 vdd.n21 0.0370523
R24629 vdd.n2947 vdd.n2946 0.0370523
R24630 vdd.n2946 vdd.n2945 0.0370523
R24631 vdd.n2945 vdd.n26 0.0370523
R24632 vdd.n2941 vdd.n26 0.0370523
R24633 vdd.n2940 vdd.n2939 0.0370523
R24634 vdd.n2939 vdd.n31 0.0370523
R24635 vdd.n2935 vdd.n31 0.0370523
R24636 vdd.n2935 vdd.n2934 0.0370523
R24637 vdd.n2934 vdd.n2933 0.0370523
R24638 vdd.n2933 vdd.n36 0.0370523
R24639 vdd.n2929 vdd.n2928 0.0370523
R24640 vdd.n2928 vdd.n2927 0.0370523
R24641 vdd.n2927 vdd.n41 0.0370523
R24642 vdd.n2923 vdd.n41 0.0370523
R24643 vdd.n2923 vdd.n2922 0.0370523
R24644 vdd.n2922 vdd.n2921 0.0370523
R24645 vdd.n2917 vdd.n46 0.0370523
R24646 vdd.n2917 vdd.n2916 0.0370523
R24647 vdd.n2916 vdd.n2915 0.0370523
R24648 vdd.n2915 vdd.n51 0.0370523
R24649 vdd.n2911 vdd.n51 0.0370523
R24650 vdd.n2911 vdd.n2910 0.0370523
R24651 vdd.n2909 vdd.n56 0.0370523
R24652 vdd.n2905 vdd.n56 0.0370523
R24653 vdd.n2905 vdd.n2904 0.0370523
R24654 vdd.n2904 vdd.n2903 0.0370523
R24655 vdd.n2903 vdd.n61 0.0370523
R24656 vdd.n2899 vdd.n61 0.0370523
R24657 vdd.n2898 vdd.n2897 0.0370523
R24658 vdd.n2897 vdd.n66 0.0370523
R24659 vdd.n2893 vdd.n66 0.0370523
R24660 vdd.n2893 vdd.n2892 0.0370523
R24661 vdd.n2892 vdd.n2891 0.0370523
R24662 vdd.n2891 vdd.n71 0.0370523
R24663 vdd.n2887 vdd.n2886 0.0370523
R24664 vdd.n2886 vdd.n2885 0.0370523
R24665 vdd.n2885 vdd.n76 0.0370523
R24666 vdd.n2881 vdd.n76 0.0370523
R24667 vdd.n2881 vdd.n2880 0.0370523
R24668 vdd.n2880 vdd.n2879 0.0370523
R24669 vdd.n2875 vdd.n81 0.0370523
R24670 vdd.n2875 vdd.n2874 0.0370523
R24671 vdd.n2874 vdd.n2873 0.0370523
R24672 vdd.n2873 vdd.n86 0.0370523
R24673 vdd.n2869 vdd.n86 0.0370523
R24674 vdd.n2869 vdd.n2868 0.0370523
R24675 vdd.n2867 vdd.n91 0.0370523
R24676 vdd.n2863 vdd.n91 0.0370523
R24677 vdd.n2863 vdd.n2862 0.0370523
R24678 vdd.n2862 vdd.n2861 0.0370523
R24679 vdd.n2861 vdd.n96 0.0370523
R24680 vdd.n2857 vdd.n96 0.0370523
R24681 vdd.n2160 vdd.n2159 0.0370523
R24682 vdd.n2161 vdd.n2160 0.0370523
R24683 vdd.n2165 vdd.n2164 0.0370523
R24684 vdd.n2166 vdd.n2165 0.0370523
R24685 vdd.n2167 vdd.n2166 0.0370523
R24686 vdd.n2170 vdd.n2167 0.0370523
R24687 vdd.n2171 vdd.n2170 0.0370523
R24688 vdd.n2172 vdd.n2171 0.0370523
R24689 vdd.n2216 vdd.n2173 0.0370523
R24690 vdd.n2218 vdd.n2216 0.0370523
R24691 vdd.n2219 vdd.n2218 0.0370523
R24692 vdd.n2220 vdd.n2219 0.0370523
R24693 vdd.n2222 vdd.n2220 0.0370523
R24694 vdd.n2222 vdd.n2221 0.0370523
R24695 vdd.n4 vdd.n3 0.0370523
R24696 vdd.n5 vdd.n4 0.0370523
R24697 vdd.n852 vdd.n851 0.0367723
R24698 vdd.n2302 vdd.n2301 0.0366011
R24699 vdd.n2374 vdd.n280 0.0364375
R24700 vdd.n1383 vdd.n1372 0.0356562
R24701 vdd.n1177 vdd.n1176 0.034875
R24702 vdd.n2303 vdd.n336 0.0343448
R24703 vdd.n2249 vdd.n1975 0.0343448
R24704 vdd.n1360 vdd.n1354 0.0340938
R24705 vdd.n1121 vdd.n979 0.0338935
R24706 vdd.n1527 vdd.n1526 0.0338935
R24707 vdd.n1725 vdd.n458 0.0338935
R24708 vdd.n1786 vdd.n1785 0.0334422
R24709 vdd.n2296 vdd.n2295 0.0334422
R24710 vdd.n2353 vdd.n2352 0.0333125
R24711 vdd.n2364 vdd.n284 0.0333125
R24712 vdd.n2489 vdd.n5 0.0332117
R24713 vdd.n1179 vdd.n679 0.0325312
R24714 vdd.n1208 vdd.n664 0.0325312
R24715 vdd.n1238 vdd.n649 0.0325312
R24716 vdd.n1267 vdd.n634 0.0325312
R24717 vdd.n1505 vdd.n1504 0.0325312
R24718 vdd.n1470 vdd.n1313 0.0325312
R24719 vdd.n1442 vdd.n1329 0.0325312
R24720 vdd.n1414 vdd.n1345 0.0325312
R24721 vdd.n1389 vdd.n1364 0.0325312
R24722 vdd.n2344 vdd.n293 0.0325312
R24723 vdd.n2377 vdd.n281 0.0325312
R24724 vdd.n2409 vdd.n269 0.0325312
R24725 vdd.n2442 vdd.n257 0.0325312
R24726 vdd.n2473 vdd.n244 0.0325312
R24727 vdd.n1391 vdd.n1366 0.0325312
R24728 vdd.n856 vdd.n855 0.032308
R24729 vdd.n1502 vdd.n1501 0.0320345
R24730 vdd.n2341 vdd.n2340 0.0320345
R24731 vdd.n2338 vdd.n302 0.0320345
R24732 vdd.n1493 vdd.n1492 0.0320345
R24733 vdd.n870 vdd.n869 0.031192
R24734 vdd.n2254 vdd.n1970 0.0311859
R24735 vdd.n841 vdd.n815 0.0311837
R24736 vdd.n1179 vdd.n1178 0.0309688
R24737 vdd.n1208 vdd.n1207 0.0309688
R24738 vdd.n1238 vdd.n1237 0.0309688
R24739 vdd.n1267 vdd.n1266 0.0309688
R24740 vdd.n1505 vdd.n622 0.0309688
R24741 vdd.n1471 vdd.n1470 0.0309688
R24742 vdd.n1443 vdd.n1442 0.0309688
R24743 vdd.n1417 vdd.n1345 0.0309688
R24744 vdd.n1392 vdd.n1364 0.0309688
R24745 vdd.n2377 vdd.n2376 0.0309688
R24746 vdd.n2409 vdd.n2408 0.0309688
R24747 vdd.n2442 vdd.n2441 0.0309688
R24748 vdd.n2473 vdd.n2472 0.0309688
R24749 vdd.n1366 vdd.n1361 0.0309688
R24750 vdd.n1706 vdd.n480 0.0307347
R24751 vdd.n1912 vdd.n1911 0.0307347
R24752 vdd.n2202 vdd.n2182 0.0305117
R24753 vdd.n1126 vdd.n973 0.0302834
R24754 vdd.n1532 vdd.n588 0.0302834
R24755 vdd.n1780 vdd.n1779 0.0302834
R24756 vdd.n2352 vdd.n288 0.0301875
R24757 vdd.n2365 vdd.n2364 0.0301875
R24758 vdd.n1929 vdd.n1926 0.0298321
R24759 vdd.n1399 vdd.n1360 0.0294063
R24760 vdd.n2202 vdd.n2201 0.0292978
R24761 vdd.n1176 vdd.n1175 0.028625
R24762 vdd.n859 vdd.n849 0.0278438
R24763 vdd.n1372 vdd.n1367 0.0278438
R24764 vdd.n1792 vdd.n453 0.0276448
R24765 vdd.n1870 vdd.n370 0.0275758
R24766 vdd.n2259 vdd.n1964 0.0275758
R24767 vdd.n1131 vdd.n967 0.0271245
R24768 vdd.n1547 vdd.n585 0.0271245
R24769 vdd.n1693 vdd.n493 0.0271245
R24770 vdd.n2375 vdd.n2374 0.0270625
R24771 vdd.n866 vdd.n845 0.0267277
R24772 vdd.n1737 vdd.n1734 0.0266733
R24773 vdd.n2287 vdd.n1934 0.0266733
R24774 vdd.n1796 vdd.n453 0.0265125
R24775 vdd.n1178 vdd.n681 0.0262812
R24776 vdd.n1207 vdd.n666 0.0262812
R24777 vdd.n1237 vdd.n651 0.0262812
R24778 vdd.n1266 vdd.n636 0.0262812
R24779 vdd.n1291 vdd.n622 0.0262812
R24780 vdd.n1471 vdd.n1310 0.0262812
R24781 vdd.n1443 vdd.n1326 0.0262812
R24782 vdd.n1418 vdd.n1417 0.0262812
R24783 vdd.n1393 vdd.n1392 0.0262812
R24784 vdd.n2376 vdd.n283 0.0262812
R24785 vdd.n2408 vdd.n271 0.0262812
R24786 vdd.n2441 vdd.n259 0.0262812
R24787 vdd.n2472 vdd.n246 0.0262812
R24788 vdd.n1408 vdd.n1353 0.0262812
R24789 vdd.n1185 vdd.n1184 0.0255
R24790 vdd.n2561 vdd.n2493 0.0250902
R24791 vdd.n2588 vdd.n218 0.0250902
R24792 vdd.n2610 vdd.n192 0.0250902
R24793 vdd.n2635 vdd.n167 0.0250902
R24794 vdd.n2797 vdd.n2796 0.0250902
R24795 vdd.n2742 vdd.n2741 0.0250902
R24796 vdd.n2854 vdd.n98 0.0250902
R24797 vdd.n2315 vdd.n2314 0.0250232
R24798 vdd.n2074 vdd.n2044 0.0250232
R24799 vdd.n2099 vdd.n2022 0.0250232
R24800 vdd.n2125 vdd.n2003 0.0250232
R24801 vdd.n2150 vdd.n1983 0.0250232
R24802 vdd.n1822 vdd.n425 0.0250232
R24803 vdd.n1847 vdd.n397 0.0250232
R24804 vdd.n1899 vdd.n353 0.0250232
R24805 vdd.n2584 vdd.n28 0.0247486
R24806 vdd.n2613 vdd.n38 0.0247486
R24807 vdd.n1182 vdd.n679 0.0247187
R24808 vdd.n1211 vdd.n664 0.0247187
R24809 vdd.n1241 vdd.n649 0.0247187
R24810 vdd.n1270 vdd.n634 0.0247187
R24811 vdd.n1467 vdd.n1313 0.0247187
R24812 vdd.n1439 vdd.n1329 0.0247187
R24813 vdd.n1414 vdd.n1413 0.0247187
R24814 vdd.n1389 vdd.n1388 0.0247187
R24815 vdd.n2348 vdd.n293 0.0247187
R24816 vdd.n2380 vdd.n281 0.0247187
R24817 vdd.n2413 vdd.n269 0.0247187
R24818 vdd.n2445 vdd.n257 0.0247187
R24819 vdd.n2476 vdd.n244 0.0247187
R24820 vdd.n1374 vdd.n1373 0.0247187
R24821 vdd.n2311 vdd.n325 0.0246826
R24822 vdd.n1869 vdd.n1868 0.0246826
R24823 vdd.n2264 vdd.n1958 0.024417
R24824 vdd.n2538 vdd.n18 0.0244071
R24825 vdd.n2638 vdd.n48 0.0244071
R24826 vdd.n2850 vdd.n107 0.0244071
R24827 vdd.n2077 vdd.n1924 0.024342
R24828 vdd.n1843 vdd.n405 0.024342
R24829 vdd.n946 vdd.n708 0.0243024
R24830 vdd.n1157 vdd.n694 0.0242936
R24831 vdd.n1070 vdd.n1021 0.0242936
R24832 vdd.n1097 vdd.n1003 0.0242936
R24833 vdd.n1519 vdd.n610 0.0242936
R24834 vdd.n596 vdd.n595 0.0242936
R24835 vdd.n568 vdd.n561 0.0242936
R24836 vdd.n1685 vdd.n496 0.0242936
R24837 vdd.n1718 vdd.n456 0.0242936
R24838 vdd.n2490 vdd.n8 0.0240656
R24839 vdd.n2793 vdd.n58 0.0240656
R24840 vdd.n2820 vdd.n128 0.0240656
R24841 vdd.n2102 vdd.n1938 0.0240014
R24842 vdd.n2146 vdd.n1968 0.0240014
R24843 vdd.n1818 vdd.n431 0.0240014
R24844 vdd.n1666 vdd.n1665 0.0239657
R24845 vdd.n1753 vdd.n1748 0.0239657
R24846 vdd.n1094 vdd.n976 0.0239584
R24847 vdd.n1576 vdd.n557 0.0239584
R24848 vdd.n2385 vdd.n2384 0.0239375
R24849 vdd.n2763 vdd.n68 0.023724
R24850 vdd.n1067 vdd.n959 0.0236233
R24851 vdd.n1136 vdd.n961 0.0235144
R24852 vdd.n1572 vdd.n564 0.0235144
R24853 vdd.n1771 vdd.n1739 0.0235144
R24854 vdd.n2282 vdd.n1940 0.0235144
R24855 vdd.n2771 vdd.n2679 0.0233825
R24856 vdd.n2738 vdd.n78 0.0233825
R24857 vdd.n862 vdd.n847 0.0233795
R24858 vdd.n2121 vdd.n1954 0.0233202
R24859 vdd.n2128 vdd.n1955 0.0233202
R24860 vdd.n1799 vdd.n450 0.0233202
R24861 vdd.n943 vdd.n692 0.0232882
R24862 vdd.n467 vdd.n464 0.0232882
R24863 vdd.n1416 vdd.n1347 0.0231563
R24864 vdd.n2557 vdd.n9 0.023041
R24865 vdd.n2829 vdd.n88 0.023041
R24866 vdd.n2095 vdd.n1937 0.0229796
R24867 vdd.n2153 vdd.n1972 0.0229796
R24868 vdd.n1825 vdd.n422 0.0229796
R24869 vdd.n1682 vdd.n1681 0.0229531
R24870 vdd.n1689 vdd.n490 0.0229531
R24871 vdd.n2530 vdd.n19 0.0226995
R24872 vdd.n2631 vdd.n173 0.0226995
R24873 vdd.n2070 vdd.n1922 0.022639
R24874 vdd.n1850 vdd.n394 0.022639
R24875 vdd.n701 vdd.n699 0.022618
R24876 vdd.n1196 vdd.n1195 0.022375
R24877 vdd.n2318 vdd.n318 0.0222984
R24878 vdd.n1019 vdd.n963 0.0222828
R24879 vdd.n1651 vdd.n527 0.0222828
R24880 vdd.n865 vdd.n847 0.0222634
R24881 vdd.n2606 vdd.n201 0.0220164
R24882 vdd.n1571 vdd.n567 0.0219477
R24883 vdd.n2616 vdd.n39 0.0216749
R24884 vdd.n2308 vdd.n329 0.0216172
R24885 vdd.n1865 vdd.n371 0.0216172
R24886 vdd.n1000 vdd.n977 0.0216126
R24887 vdd.n2541 vdd.n2514 0.0213333
R24888 vdd.n603 vdd.n600 0.0212775
R24889 vdd.n1534 vdd.n1533 0.0212775
R24890 vdd.n2080 vdd.n1925 0.0212766
R24891 vdd.n1840 vdd.n400 0.0212766
R24892 vdd.n2800 vdd.n2656 0.0209918
R24893 vdd.n2790 vdd.n59 0.0209918
R24894 vdd.n2817 vdd.n85 0.0209918
R24895 vdd.n1091 vdd.n975 0.0209424
R24896 vdd.n559 vdd.n554 0.0209424
R24897 vdd.n2397 vdd.n2396 0.0208125
R24898 vdd.n1149 vdd.n706 0.0208069
R24899 vdd.n1646 vdd.n537 0.0208069
R24900 vdd.n1758 vdd.n1745 0.0208069
R24901 vdd.n2269 vdd.n1952 0.0208069
R24902 vdd.n2760 vdd.n69 0.0206503
R24903 vdd.n2748 vdd.n75 0.0206503
R24904 vdd.n1064 vdd.n958 0.0206072
R24905 vdd.n2105 vdd.n1942 0.0205954
R24906 vdd.n2143 vdd.n1967 0.0205954
R24907 vdd.n1815 vdd.n428 0.0205954
R24908 vdd.n2192 vdd.n2190 0.0203873
R24909 vdd.n2192 vdd.n2191 0.0203873
R24910 vdd.n2195 vdd.n2193 0.0203873
R24911 vdd.n2195 vdd.n2194 0.0203873
R24912 vdd.n2197 vdd.n2196 0.0203873
R24913 vdd.n2194 vdd.n2187 0.0203873
R24914 vdd.n2191 vdd.n2188 0.0203873
R24915 vdd.n2196 vdd.n2187 0.0203873
R24916 vdd.n2193 vdd.n2188 0.0203873
R24917 vdd.n1141 vdd.n955 0.0203556
R24918 vdd.n1585 vdd.n551 0.0203556
R24919 vdd.n1766 vdd.n1742 0.0203556
R24920 vdd.n2774 vdd.n65 0.0203087
R24921 vdd.n2735 vdd.n79 0.0203087
R24922 vdd.n1723 vdd.n463 0.0202721
R24923 vdd.n2117 vdd.n1950 0.0202548
R24924 vdd.n2131 vdd.n1956 0.0202548
R24925 vdd.n1802 vdd.n447 0.0202548
R24926 vdd.n781 vdd.n765 0.0201221
R24927 vdd.n781 vdd.n721 0.0201221
R24928 vdd.n928 vdd.n721 0.0201221
R24929 vdd.n933 vdd.n719 0.0201221
R24930 vdd.n933 vdd.n708 0.0201221
R24931 vdd.n1174 vdd.n1173 0.0200312
R24932 vdd.n1203 vdd.n1202 0.0200312
R24933 vdd.n1233 vdd.n1232 0.0200312
R24934 vdd.n1262 vdd.n1261 0.0200312
R24935 vdd.n1292 vdd.n1290 0.0200312
R24936 vdd.n1476 vdd.n1475 0.0200312
R24937 vdd.n1448 vdd.n1447 0.0200312
R24938 vdd.n1421 vdd.n1343 0.0200312
R24939 vdd.n1396 vdd.n1362 0.0200312
R24940 vdd.n2371 vdd.n2370 0.0200312
R24941 vdd.n2403 vdd.n2402 0.0200312
R24942 vdd.n2436 vdd.n2435 0.0200312
R24943 vdd.n2468 vdd.n2467 0.0200312
R24944 vdd.n1424 vdd.n1341 0.0200312
R24945 vdd.n2803 vdd.n55 0.0199672
R24946 vdd.n2832 vdd.n89 0.0199672
R24947 vdd.n1678 vdd.n505 0.019937
R24948 vdd.n1694 vdd.n486 0.019937
R24949 vdd.n2092 vdd.n1936 0.0199142
R24950 vdd.n2156 vdd.n1973 0.0199142
R24951 vdd.n1828 vdd.n419 0.0199142
R24952 vdd.n2277 vdd.n1946 0.0199043
R24953 vdd.n2580 vdd.n221 0.0196257
R24954 vdd.n1150 vdd.n703 0.0196019
R24955 vdd.n2067 vdd.n2047 0.0195736
R24956 vdd.n1853 vdd.n391 0.0195736
R24957 vdd.n1612 vdd.n521 0.019426
R24958 vdd.n1890 vdd.n363 0.019426
R24959 vdd.n1610 vdd.n521 0.019426
R24960 vdd.n1888 vdd.n363 0.019426
R24961 vdd.n2502 vdd.n10 0.0192842
R24962 vdd.n2525 vdd.n20 0.0192842
R24963 vdd.n2628 vdd.n45 0.0192842
R24964 vdd.n1648 vdd.n1647 0.0192668
R24965 vdd.n1655 vdd.n529 0.0192668
R24966 vdd.n1205 vdd.n1204 0.01925
R24967 vdd.n348 vdd.n315 0.019233
R24968 vdd.n1601 vdd.n523 0.0192022
R24969 vdd.n1602 vdd.n1601 0.0192022
R24970 vdd.n1608 vdd.n522 0.0192022
R24971 vdd.n1608 vdd.n1603 0.0192022
R24972 vdd.n1612 vdd.n1604 0.0192022
R24973 vdd.n1605 vdd.n520 0.0192022
R24974 vdd.n1619 vdd.n1605 0.0192022
R24975 vdd.n519 vdd.n518 0.0192022
R24976 vdd.n518 vdd.n516 0.0192022
R24977 vdd.n1894 vdd.n364 0.0192022
R24978 vdd.n1893 vdd.n368 0.0192022
R24979 vdd.n1888 vdd.n1887 0.0192022
R24980 vdd.n1875 vdd.n362 0.0192022
R24981 vdd.n1878 vdd.n1876 0.0192022
R24982 vdd.n1880 vdd.n361 0.0192022
R24983 vdd.n1885 vdd.n1877 0.0192022
R24984 vdd.n1884 vdd.n360 0.0192022
R24985 vdd.n1661 vdd.n516 0.0192022
R24986 vdd.n1619 vdd.n1618 0.0192022
R24987 vdd.n1614 vdd.n1604 0.0192022
R24988 vdd.n1610 vdd.n1603 0.0192022
R24989 vdd.n1606 vdd.n1602 0.0192022
R24990 vdd.n1642 vdd.n523 0.0192022
R24991 vdd.n1606 vdd.n522 0.0192022
R24992 vdd.n1614 vdd.n520 0.0192022
R24993 vdd.n1618 vdd.n519 0.0192022
R24994 vdd.n1885 vdd.n1884 0.0192022
R24995 vdd.n1880 vdd.n1876 0.0192022
R24996 vdd.n1887 vdd.n1875 0.0192022
R24997 vdd.n1890 vdd.n368 0.0192022
R24998 vdd.n1894 vdd.n1893 0.0192022
R24999 vdd.n1878 vdd.n362 0.0192022
R25000 vdd.n1877 vdd.n361 0.0192022
R25001 vdd.n360 vdd.n341 0.0192022
R25002 vdd.n810 vdd.n759 0.0189511
R25003 vdd.n2594 vdd.n30 0.0189426
R25004 vdd.n2603 vdd.n35 0.0189426
R25005 vdd.n2745 vdd.n2705 0.0189426
R25006 vdd.n1017 vdd.n964 0.0189316
R25007 vdd.n866 vdd.n865 0.0189152
R25008 vdd.n774 vdd.n773 0.0186219
R25009 vdd.n2576 vdd.n25 0.0186011
R25010 vdd.n2619 vdd.n40 0.0186011
R25011 vdd.n1110 vdd.n981 0.0185965
R25012 vdd.n1558 vdd.n1557 0.0185965
R25013 vdd.n2307 vdd.n333 0.0185518
R25014 vdd.n1862 vdd.n378 0.0185518
R25015 vdd.n1183 vdd.n676 0.0184687
R25016 vdd.n1212 vdd.n661 0.0184687
R25017 vdd.n1242 vdd.n646 0.0184687
R25018 vdd.n1272 vdd.n1271 0.0184687
R25019 vdd.n1466 vdd.n1315 0.0184687
R25020 vdd.n1438 vdd.n1331 0.0184687
R25021 vdd.n1410 vdd.n1349 0.0184687
R25022 vdd.n1385 vdd.n1368 0.0184687
R25023 vdd.n2349 vdd.n291 0.0184687
R25024 vdd.n2381 vdd.n279 0.0184687
R25025 vdd.n2414 vdd.n267 0.0184687
R25026 vdd.n2446 vdd.n255 0.0184687
R25027 vdd.n2477 vdd.n242 0.0184687
R25028 vdd.n926 vdd.n723 0.0182936
R25029 vdd.n734 vdd.n723 0.0182936
R25030 vdd.n915 vdd.n734 0.0182936
R25031 vdd.n915 vdd.n914 0.0182936
R25032 vdd.n914 vdd.n735 0.0182936
R25033 vdd.n748 vdd.n735 0.0182936
R25034 vdd.n903 vdd.n748 0.0182936
R25035 vdd.n903 vdd.n902 0.0182936
R25036 vdd.n824 vdd.n823 0.0182936
R25037 vdd.n890 vdd.n824 0.0182936
R25038 vdd.n890 vdd.n889 0.0182936
R25039 vdd.n889 vdd.n825 0.0182936
R25040 vdd.n836 vdd.n825 0.0182936
R25041 vdd.n878 vdd.n836 0.0182936
R25042 vdd.n878 vdd.n877 0.0182936
R25043 vdd.n877 vdd.n837 0.0182936
R25044 vdd.n1524 vdd.n599 0.0182614
R25045 vdd.n1540 vdd.n1539 0.0182614
R25046 vdd.n2641 vdd.n162 0.0182596
R25047 vdd.n2644 vdd.n50 0.0182596
R25048 vdd.n2841 vdd.n94 0.0182596
R25049 vdd.n1088 vdd.n971 0.0179263
R25050 vdd.n1584 vdd.n548 0.0179263
R25051 vdd.n2785 vdd.n60 0.017918
R25052 vdd.n2845 vdd.n95 0.017918
R25053 vdd.n784 vdd.n782 0.0179116
R25054 vdd.n2083 vdd.n2037 0.0178706
R25055 vdd.n1837 vdd.n407 0.0178706
R25056 vdd.n770 vdd.n762 0.0177982
R25057 vdd.n2407 vdd.n2406 0.0176875
R25058 vdd.n1763 vdd.n1742 0.017648
R25059 vdd.n2274 vdd.n1946 0.017648
R25060 vdd.n1061 vdd.n957 0.0175912
R25061 vdd.n2757 vdd.n70 0.0175765
R25062 vdd.n2751 vdd.n74 0.0175765
R25063 vdd.n2108 vdd.n1943 0.01753
R25064 vdd.n2140 vdd.n1966 0.01753
R25065 vdd.n1812 vdd.n435 0.01753
R25066 vdd.n945 vdd.n709 0.0173375
R25067 vdd.n1713 vdd.n475 0.017256
R25068 vdd.n2730 vdd.n80 0.017235
R25069 vdd.n1146 vdd.n706 0.0171968
R25070 vdd.n1144 vdd.n955 0.0171968
R25071 vdd.n1588 vdd.n551 0.0171968
R25072 vdd.n1598 vdd.n537 0.0171968
R25073 vdd.n2114 vdd.n1949 0.0171894
R25074 vdd.n2134 vdd.n1960 0.0171894
R25075 vdd.n1805 vdd.n444 0.0171894
R25076 vdd.n1633 vdd.n529 0.0169209
R25077 vdd.n1675 vdd.n508 0.0169209
R25078 vdd.n488 vdd.n483 0.0169209
R25079 vdd.n1436 vdd.n1435 0.0169062
R25080 vdd.n2768 vdd.n2767 0.0168934
R25081 vdd.n921 vdd.n728 0.0168934
R25082 vdd.n921 vdd.n920 0.0168934
R25083 vdd.n920 vdd.n729 0.0168934
R25084 vdd.n740 vdd.n729 0.0168934
R25085 vdd.n909 vdd.n740 0.0168934
R25086 vdd.n909 vdd.n908 0.0168934
R25087 vdd.n908 vdd.n741 0.0168934
R25088 vdd.n752 vdd.n741 0.0168934
R25089 vdd.n896 vdd.n895 0.0168934
R25090 vdd.n895 vdd.n817 0.0168934
R25091 vdd.n830 vdd.n817 0.0168934
R25092 vdd.n884 vdd.n830 0.0168934
R25093 vdd.n884 vdd.n883 0.0168934
R25094 vdd.n883 vdd.n831 0.0168934
R25095 vdd.n842 vdd.n831 0.0168934
R25096 vdd.n872 vdd.n842 0.0168934
R25097 vdd.n2089 vdd.n1932 0.0168488
R25098 vdd.n2158 vdd.n1974 0.0168488
R25099 vdd.n1831 vdd.n416 0.0168488
R25100 vdd.n358 vdd.n342 0.0168488
R25101 vdd.n1761 vdd.n1745 0.0167455
R25102 vdd.n2272 vdd.n1952 0.0167455
R25103 vdd.n2553 vdd.n2552 0.0165519
R25104 vdd.n2651 vdd.n54 0.0165519
R25105 vdd.n2064 vdd.n1919 0.0165082
R25106 vdd.n1856 vdd.n388 0.0165082
R25107 vdd.n1050 vdd.n951 0.0162507
R25108 vdd.n2591 vdd.n215 0.0162104
R25109 vdd.n2625 vdd.n44 0.0162104
R25110 vdd.n1903 vdd.n345 0.0161676
R25111 vdd.n1214 vdd.n1213 0.016125
R25112 vdd.n2189 vdd.n2183 0.0161007
R25113 vdd.n2207 vdd.n2189 0.0161007
R25114 vdd.n1015 vdd.n965 0.0159155
R25115 vdd.n1597 vdd.n1596 0.0159155
R25116 vdd.n2597 vdd.n209 0.0158689
R25117 vdd.n2600 vdd.n34 0.0158689
R25118 vdd.n745 vdd.n744 0.0158146
R25119 vdd.n742 vdd.n739 0.0157389
R25120 vdd.n912 vdd.n736 0.0156076
R25121 vdd.n1113 vdd.n982 0.0155804
R25122 vdd.n1552 vdd.n579 0.0155804
R25123 vdd.n803 vdd.n802 0.0155728
R25124 vdd.n861 vdd.n859 0.015567
R25125 vdd.n911 vdd.n910 0.0155329
R25126 vdd.n2573 vdd.n24 0.0155273
R25127 vdd.n814 vdd.n813 0.015327
R25128 vdd.n987 vdd.n986 0.0152453
R25129 vdd.n590 vdd.n581 0.0152453
R25130 vdd.n875 vdd.n838 0.0151937
R25131 vdd.n2549 vdd.n14 0.0151858
R25132 vdd.n2647 vdd.n154 0.0151858
R25133 vdd.n2838 vdd.n93 0.0151858
R25134 vdd.n2061 vdd.n1916 0.0151458
R25135 vdd.n1859 vdd.n382 0.0151458
R25136 vdd.n874 vdd.n873 0.0151211
R25137 vdd.n1085 vdd.n970 0.0149102
R25138 vdd.n1589 vdd.n544 0.0149102
R25139 vdd.n2782 vdd.n2670 0.0148443
R25140 vdd.n2727 vdd.n83 0.0148443
R25141 vdd.n2823 vdd.n125 0.0148443
R25142 vdd.n2855 vdd.n97 0.0148443
R25143 vdd.n2086 vdd.n1930 0.0148052
R25144 vdd.n1834 vdd.n410 0.0148052
R25145 vdd.n905 vdd.n746 0.0147798
R25146 vdd.n907 vdd.n906 0.0147092
R25147 vdd.n1058 vdd.n953 0.0145751
R25148 vdd.n2418 vdd.n2417 0.0145625
R25149 vdd.n2754 vdd.n2692 0.0145027
R25150 vdd.n2279 vdd.n1940 0.0144892
R25151 vdd.n2111 vdd.n1944 0.0144646
R25152 vdd.n2137 vdd.n1962 0.0144646
R25153 vdd.n1808 vdd.n438 0.0144646
R25154 vdd.n869 vdd.n845 0.0144509
R25155 vdd.n930 vdd.n929 0.0144134
R25156 vdd.n1148 vdd.n1147 0.0144134
R25157 vdd.n1137 vdd.n962 0.0144134
R25158 vdd.n1123 vdd.n974 0.0144134
R25159 vdd.n1530 vdd.n1529 0.0144134
R25160 vdd.n1573 vdd.n565 0.0144134
R25161 vdd.n1645 vdd.n1599 0.0144134
R25162 vdd.n1613 vdd.n1611 0.0144134
R25163 vdd.n1669 vdd.n1663 0.0144134
R25164 vdd.n1704 vdd.n481 0.0144134
R25165 vdd.n1789 vdd.n1788 0.0144134
R25166 vdd.n1776 vdd.n1775 0.0144134
R25167 vdd.n1765 vdd.n1764 0.0144134
R25168 vdd.n1754 vdd.n1749 0.0144134
R25169 vdd.n1891 vdd.n1889 0.0144134
R25170 vdd.n1906 vdd.n340 0.0144134
R25171 vdd.n2305 vdd.n2304 0.0144134
R25172 vdd.n2292 vdd.n2291 0.0144134
R25173 vdd.n2281 vdd.n2280 0.0144134
R25174 vdd.n2270 vdd.n1953 0.0144134
R25175 vdd.n2256 vdd.n1965 0.0144134
R25176 vdd.n2246 vdd.n2245 0.0144134
R25177 vdd.n2234 vdd.n2169 0.0144134
R25178 vdd.n2962 vdd.n2961 0.0144134
R25179 vdd.n2950 vdd.n17 0.0144134
R25180 vdd.n2942 vdd.n27 0.0144134
R25181 vdd.n2931 vdd.n2930 0.0144134
R25182 vdd.n2920 vdd.n2919 0.0144134
R25183 vdd.n2908 vdd.n52 0.0144134
R25184 vdd.n2900 vdd.n62 0.0144134
R25185 vdd.n2889 vdd.n2888 0.0144134
R25186 vdd.n2878 vdd.n2877 0.0144134
R25187 vdd.n2866 vdd.n87 0.0144134
R25188 vdd.n913 vdd.n733 0.0143659
R25189 vdd.n738 vdd.n737 0.0142974
R25190 vdd.n772 vdd.n771 0.0142437
R25191 vdd.n779 vdd.n778 0.0142437
R25192 vdd.n780 vdd.n779 0.0142437
R25193 vdd.n780 vdd.n720 0.0142437
R25194 vdd.n929 vdd.n720 0.0142437
R25195 vdd.n932 vdd.n930 0.0142437
R25196 vdd.n932 vdd.n931 0.0142437
R25197 vdd.n931 vdd.n707 0.0142437
R25198 vdd.n948 vdd.n707 0.0142437
R25199 vdd.n949 vdd.n948 0.0142437
R25200 vdd.n1148 vdd.n949 0.0142437
R25201 vdd.n1147 vdd.n950 0.0142437
R25202 vdd.n1143 vdd.n950 0.0142437
R25203 vdd.n1143 vdd.n1142 0.0142437
R25204 vdd.n1142 vdd.n956 0.0142437
R25205 vdd.n1138 vdd.n956 0.0142437
R25206 vdd.n1138 vdd.n1137 0.0142437
R25207 vdd.n1133 vdd.n962 0.0142437
R25208 vdd.n1133 vdd.n1132 0.0142437
R25209 vdd.n1132 vdd.n968 0.0142437
R25210 vdd.n1128 vdd.n968 0.0142437
R25211 vdd.n1128 vdd.n1127 0.0142437
R25212 vdd.n1127 vdd.n974 0.0142437
R25213 vdd.n1123 vdd.n1122 0.0142437
R25214 vdd.n1122 vdd.n980 0.0142437
R25215 vdd.n1118 vdd.n980 0.0142437
R25216 vdd.n1118 vdd.n597 0.0142437
R25217 vdd.n1528 vdd.n597 0.0142437
R25218 vdd.n1529 vdd.n1528 0.0142437
R25219 vdd.n1530 vdd.n586 0.0142437
R25220 vdd.n1542 vdd.n586 0.0142437
R25221 vdd.n1543 vdd.n1542 0.0142437
R25222 vdd.n1546 vdd.n1543 0.0142437
R25223 vdd.n1546 vdd.n1545 0.0142437
R25224 vdd.n1545 vdd.n565 0.0142437
R25225 vdd.n1574 vdd.n1573 0.0142437
R25226 vdd.n1574 vdd.n552 0.0142437
R25227 vdd.n1586 vdd.n552 0.0142437
R25228 vdd.n1587 vdd.n1586 0.0142437
R25229 vdd.n1587 vdd.n539 0.0142437
R25230 vdd.n1599 vdd.n539 0.0142437
R25231 vdd.n1645 vdd.n1644 0.0142437
R25232 vdd.n1644 vdd.n1643 0.0142437
R25233 vdd.n1643 vdd.n1600 0.0142437
R25234 vdd.n1607 vdd.n1600 0.0142437
R25235 vdd.n1609 vdd.n1607 0.0142437
R25236 vdd.n1611 vdd.n1609 0.0142437
R25237 vdd.n1615 vdd.n1613 0.0142437
R25238 vdd.n1616 vdd.n1615 0.0142437
R25239 vdd.n1617 vdd.n1616 0.0142437
R25240 vdd.n1617 vdd.n514 0.0142437
R25241 vdd.n1662 vdd.n514 0.0142437
R25242 vdd.n1663 vdd.n1662 0.0142437
R25243 vdd.n1669 vdd.n1668 0.0142437
R25244 vdd.n1668 vdd.n1667 0.0142437
R25245 vdd.n1667 vdd.n494 0.0142437
R25246 vdd.n1691 vdd.n494 0.0142437
R25247 vdd.n1692 vdd.n1691 0.0142437
R25248 vdd.n1692 vdd.n481 0.0142437
R25249 vdd.n1705 vdd.n1704 0.0142437
R25250 vdd.n1705 vdd.n461 0.0142437
R25251 vdd.n1727 vdd.n461 0.0142437
R25252 vdd.n1728 vdd.n1727 0.0142437
R25253 vdd.n1790 vdd.n1728 0.0142437
R25254 vdd.n1790 vdd.n1789 0.0142437
R25255 vdd.n1788 vdd.n1729 0.0142437
R25256 vdd.n1783 vdd.n1729 0.0142437
R25257 vdd.n1783 vdd.n1782 0.0142437
R25258 vdd.n1782 vdd.n1781 0.0142437
R25259 vdd.n1781 vdd.n1732 0.0142437
R25260 vdd.n1776 vdd.n1732 0.0142437
R25261 vdd.n1775 vdd.n1774 0.0142437
R25262 vdd.n1774 vdd.n1735 0.0142437
R25263 vdd.n1770 vdd.n1735 0.0142437
R25264 vdd.n1770 vdd.n1769 0.0142437
R25265 vdd.n1769 vdd.n1740 0.0142437
R25266 vdd.n1765 vdd.n1740 0.0142437
R25267 vdd.n1764 vdd.n1743 0.0142437
R25268 vdd.n1760 vdd.n1743 0.0142437
R25269 vdd.n1760 vdd.n1759 0.0142437
R25270 vdd.n1759 vdd.n1746 0.0142437
R25271 vdd.n1755 vdd.n1746 0.0142437
R25272 vdd.n1755 vdd.n1754 0.0142437
R25273 vdd.n1750 vdd.n1749 0.0142437
R25274 vdd.n1750 vdd.n369 0.0142437
R25275 vdd.n1872 vdd.n369 0.0142437
R25276 vdd.n1873 vdd.n1872 0.0142437
R25277 vdd.n1892 vdd.n1873 0.0142437
R25278 vdd.n1892 vdd.n1891 0.0142437
R25279 vdd.n1889 vdd.n1874 0.0142437
R25280 vdd.n1879 vdd.n1874 0.0142437
R25281 vdd.n1881 vdd.n1879 0.0142437
R25282 vdd.n1882 vdd.n1881 0.0142437
R25283 vdd.n1883 vdd.n1882 0.0142437
R25284 vdd.n1883 vdd.n340 0.0142437
R25285 vdd.n1907 vdd.n1906 0.0142437
R25286 vdd.n1908 vdd.n1907 0.0142437
R25287 vdd.n1908 vdd.n337 0.0142437
R25288 vdd.n1913 vdd.n337 0.0142437
R25289 vdd.n1914 vdd.n1913 0.0142437
R25290 vdd.n2305 vdd.n1914 0.0142437
R25291 vdd.n2304 vdd.n1915 0.0142437
R25292 vdd.n2299 vdd.n1915 0.0142437
R25293 vdd.n2299 vdd.n2298 0.0142437
R25294 vdd.n2298 vdd.n2297 0.0142437
R25295 vdd.n2297 vdd.n1921 0.0142437
R25296 vdd.n2292 vdd.n1921 0.0142437
R25297 vdd.n2291 vdd.n2290 0.0142437
R25298 vdd.n2290 vdd.n1927 0.0142437
R25299 vdd.n2286 vdd.n1927 0.0142437
R25300 vdd.n2286 vdd.n2285 0.0142437
R25301 vdd.n2285 vdd.n1935 0.0142437
R25302 vdd.n2281 vdd.n1935 0.0142437
R25303 vdd.n2280 vdd.n1941 0.0142437
R25304 vdd.n2276 vdd.n1941 0.0142437
R25305 vdd.n2276 vdd.n2275 0.0142437
R25306 vdd.n2275 vdd.n1947 0.0142437
R25307 vdd.n2271 vdd.n1947 0.0142437
R25308 vdd.n2271 vdd.n2270 0.0142437
R25309 vdd.n2266 vdd.n1953 0.0142437
R25310 vdd.n2266 vdd.n2265 0.0142437
R25311 vdd.n2265 vdd.n1959 0.0142437
R25312 vdd.n2261 vdd.n1959 0.0142437
R25313 vdd.n2261 vdd.n2260 0.0142437
R25314 vdd.n2260 vdd.n1965 0.0142437
R25315 vdd.n2256 vdd.n2255 0.0142437
R25316 vdd.n2255 vdd.n1971 0.0142437
R25317 vdd.n2251 vdd.n1971 0.0142437
R25318 vdd.n2251 vdd.n2250 0.0142437
R25319 vdd.n2250 vdd.n1976 0.0142437
R25320 vdd.n2246 vdd.n1976 0.0142437
R25321 vdd.n2245 vdd.n2244 0.0142437
R25322 vdd.n2244 vdd.n2163 0.0142437
R25323 vdd.n2240 vdd.n2163 0.0142437
R25324 vdd.n2240 vdd.n2239 0.0142437
R25325 vdd.n2239 vdd.n2238 0.0142437
R25326 vdd.n2238 vdd.n2169 0.0142437
R25327 vdd.n2234 vdd.n2233 0.0142437
R25328 vdd.n2972 vdd.n1 0.0142437
R25329 vdd.n2968 vdd.n1 0.0142437
R25330 vdd.n2968 vdd.n2967 0.0142437
R25331 vdd.n2967 vdd.n2966 0.0142437
R25332 vdd.n2966 vdd.n7 0.0142437
R25333 vdd.n2962 vdd.n7 0.0142437
R25334 vdd.n2961 vdd.n2960 0.0142437
R25335 vdd.n2960 vdd.n12 0.0142437
R25336 vdd.n2956 vdd.n12 0.0142437
R25337 vdd.n2956 vdd.n2955 0.0142437
R25338 vdd.n2955 vdd.n2954 0.0142437
R25339 vdd.n2954 vdd.n17 0.0142437
R25340 vdd.n2950 vdd.n2949 0.0142437
R25341 vdd.n2949 vdd.n2948 0.0142437
R25342 vdd.n2948 vdd.n22 0.0142437
R25343 vdd.n2944 vdd.n22 0.0142437
R25344 vdd.n2944 vdd.n2943 0.0142437
R25345 vdd.n2943 vdd.n2942 0.0142437
R25346 vdd.n2938 vdd.n27 0.0142437
R25347 vdd.n2938 vdd.n2937 0.0142437
R25348 vdd.n2937 vdd.n2936 0.0142437
R25349 vdd.n2936 vdd.n32 0.0142437
R25350 vdd.n2932 vdd.n32 0.0142437
R25351 vdd.n2932 vdd.n2931 0.0142437
R25352 vdd.n2930 vdd.n37 0.0142437
R25353 vdd.n2926 vdd.n37 0.0142437
R25354 vdd.n2926 vdd.n2925 0.0142437
R25355 vdd.n2925 vdd.n2924 0.0142437
R25356 vdd.n2924 vdd.n42 0.0142437
R25357 vdd.n2920 vdd.n42 0.0142437
R25358 vdd.n2919 vdd.n2918 0.0142437
R25359 vdd.n2918 vdd.n47 0.0142437
R25360 vdd.n2914 vdd.n47 0.0142437
R25361 vdd.n2914 vdd.n2913 0.0142437
R25362 vdd.n2913 vdd.n2912 0.0142437
R25363 vdd.n2912 vdd.n52 0.0142437
R25364 vdd.n2908 vdd.n2907 0.0142437
R25365 vdd.n2907 vdd.n2906 0.0142437
R25366 vdd.n2906 vdd.n57 0.0142437
R25367 vdd.n2902 vdd.n57 0.0142437
R25368 vdd.n2902 vdd.n2901 0.0142437
R25369 vdd.n2901 vdd.n2900 0.0142437
R25370 vdd.n2896 vdd.n62 0.0142437
R25371 vdd.n2896 vdd.n2895 0.0142437
R25372 vdd.n2895 vdd.n2894 0.0142437
R25373 vdd.n2894 vdd.n67 0.0142437
R25374 vdd.n2890 vdd.n67 0.0142437
R25375 vdd.n2890 vdd.n2889 0.0142437
R25376 vdd.n2888 vdd.n72 0.0142437
R25377 vdd.n2884 vdd.n72 0.0142437
R25378 vdd.n2884 vdd.n2883 0.0142437
R25379 vdd.n2883 vdd.n2882 0.0142437
R25380 vdd.n2882 vdd.n77 0.0142437
R25381 vdd.n2878 vdd.n77 0.0142437
R25382 vdd.n2877 vdd.n2876 0.0142437
R25383 vdd.n2876 vdd.n82 0.0142437
R25384 vdd.n2872 vdd.n82 0.0142437
R25385 vdd.n2872 vdd.n2871 0.0142437
R25386 vdd.n2871 vdd.n2870 0.0142437
R25387 vdd.n2870 vdd.n87 0.0142437
R25388 vdd.n2866 vdd.n2865 0.0142437
R25389 vdd.n2865 vdd.n2864 0.0142437
R25390 vdd.n2864 vdd.n92 0.0142437
R25391 vdd.n2860 vdd.n92 0.0142437
R25392 vdd.n2860 vdd.n2859 0.0142437
R25393 vdd.n1636 vdd.n510 0.0142399
R25394 vdd.n1708 vdd.n1707 0.0142399
R25395 vdd.n2111 vdd.n1948 0.014124
R25396 vdd.n2137 vdd.n1961 0.014124
R25397 vdd.n1808 vdd.n441 0.014124
R25398 vdd.n1139 vdd.n961 0.0140379
R25399 vdd.n1575 vdd.n564 0.0140379
R25400 vdd.n1768 vdd.n1739 0.0140379
R25401 vdd.n876 vdd.n835 0.013952
R25402 vdd.n1672 vdd.n1671 0.0139048
R25403 vdd.n840 vdd.n839 0.0138855
R25404 vdd.n2782 vdd.n63 0.0138197
R25405 vdd.n2727 vdd.n2719 0.0138197
R25406 vdd.n2086 vdd.n1931 0.0137834
R25407 vdd.n1834 vdd.n413 0.0137834
R25408 vdd.n1170 vdd.n684 0.0137813
R25409 vdd.n1199 vdd.n669 0.0137813
R25410 vdd.n1228 vdd.n654 0.0137813
R25411 vdd.n1258 vdd.n639 0.0137813
R25412 vdd.n1287 vdd.n624 0.0137813
R25413 vdd.n1479 vdd.n1307 0.0137813
R25414 vdd.n1451 vdd.n1323 0.0137813
R25415 vdd.n1422 vdd.n1338 0.0137813
R25416 vdd.n1397 vdd.n1358 0.0137813
R25417 vdd.n2332 vdd.n2331 0.0137813
R25418 vdd.n2367 vdd.n285 0.0137813
R25419 vdd.n2399 vdd.n273 0.0137813
R25420 vdd.n2432 vdd.n261 0.0137813
R25421 vdd.n2464 vdd.n249 0.0137813
R25422 vdd.n1445 vdd.n1444 0.0137813
R25423 vdd.n1640 vdd.n1620 0.013753
R25424 vdd.n366 vdd.n351 0.013753
R25425 vdd.n1665 vdd.n513 0.0135866
R25426 vdd.n1756 vdd.n1748 0.0135866
R25427 vdd.n927 vdd.n719 0.0135814
R25428 vdd.n1702 vdd.n477 0.0135697
R25429 vdd.n904 vdd.n747 0.0135381
R25430 vdd.n939 vdd.n715 0.0134938
R25431 vdd.n2549 vdd.n13 0.0134781
R25432 vdd.n2535 vdd.n2534 0.0134781
R25433 vdd.n2647 vdd.n53 0.0134781
R25434 vdd.n2838 vdd.n113 0.0134781
R25435 vdd.n751 vdd.n743 0.0134736
R25436 vdd.n1660 vdd.n1659 0.0134518
R25437 vdd.n1895 vdd.n297 0.0134518
R25438 vdd.n2061 vdd.n1917 0.0134428
R25439 vdd.n1859 vdd.n385 0.0134428
R25440 vdd.n844 vdd.n815 0.0133348
R25441 vdd.n856 vdd.n849 0.0133348
R25442 vdd.n1031 vdd.n952 0.0132346
R25443 vdd.n2573 vdd.n23 0.0131366
R25444 vdd.n2622 vdd.n43 0.0131366
R25445 vdd.n117 vdd.n90 0.0131366
R25446 vdd.n2267 vdd.n1958 0.0131354
R25447 vdd.n917 vdd.n916 0.0131242
R25448 vdd.n918 vdd.n730 0.0130618
R25449 vdd.n1225 vdd.n1224 0.013
R25450 vdd.n1013 vdd.n969 0.0128995
R25451 vdd.n1593 vdd.n546 0.0128995
R25452 vdd.n2597 vdd.n33 0.0127951
R25453 vdd.n880 vdd.n879 0.0127103
R25454 vdd.n2213 vdd.n2175 0.0127019
R25455 vdd.n881 vdd.n832 0.0126499
R25456 vdd.n2159 vdd.n2158 0.0126251
R25457 vdd.n1117 vdd.n1116 0.0125643
R25458 vdd.n1549 vdd.n1548 0.0125643
R25459 vdd.n2570 vdd.n23 0.0124536
R25460 vdd.n2625 vdd.n43 0.0124536
R25461 vdd.n1904 vdd.n1903 0.012421
R25462 vdd.n1117 vdd.n984 0.0122292
R25463 vdd.n1548 vdd.n577 0.0122292
R25464 vdd.n1189 vdd.n1187 0.0122188
R25465 vdd.n1218 vdd.n1216 0.0122188
R25466 vdd.n1248 vdd.n1246 0.0122188
R25467 vdd.n1277 vdd.n631 0.0122188
R25468 vdd.n1490 vdd.n1489 0.0122188
R25469 vdd.n1462 vdd.n1461 0.0122188
R25470 vdd.n1434 vdd.n1433 0.0122188
R25471 vdd.n1409 vdd.n1351 0.0122188
R25472 vdd.n1384 vdd.n1370 0.0122188
R25473 vdd.n2356 vdd.n2354 0.0122188
R25474 vdd.n2388 vdd.n2386 0.0122188
R25475 vdd.n2421 vdd.n2419 0.0122188
R25476 vdd.n2453 vdd.n2451 0.0122188
R25477 vdd.n2552 vdd.n13 0.012112
R25478 vdd.n2545 vdd.n15 0.012112
R25479 vdd.n2534 vdd.n2533 0.012112
R25480 vdd.n2754 vdd.n2697 0.012112
R25481 vdd.n2835 vdd.n113 0.012112
R25482 vdd.n2208 vdd.n2177 0.0120994
R25483 vdd.n2229 vdd.n2228 0.0120994
R25484 vdd.n2064 vdd.n1917 0.0120804
R25485 vdd.n1856 vdd.n385 0.0120804
R25486 vdd.n1082 vdd.n969 0.0118941
R25487 vdd.n546 vdd.n541 0.0118941
R25488 vdd.n732 vdd.n731 0.0118825
R25489 vdd.n919 vdd.n727 0.0118262
R25490 vdd.n2779 vdd.n63 0.0117705
R25491 vdd.n2730 vdd.n2719 0.0117705
R25492 vdd.n2089 vdd.n1931 0.0117398
R25493 vdd.n1831 vdd.n413 0.0117398
R25494 vdd.n776 vdd.n775 0.0116225
R25495 vdd.n769 vdd.n768 0.0116225
R25496 vdd.n777 vdd.n776 0.0116225
R25497 vdd.n777 vdd.n769 0.0116225
R25498 vdd.n1055 vdd.n952 0.011559
R25499 vdd.n2199 vdd.n2185 0.0114968
R25500 vdd.n834 vdd.n833 0.0114685
R25501 vdd.n2430 vdd.n2429 0.0114375
R25502 vdd.n2524 vdd.n234 0.011429
R25503 vdd.n2651 vdd.n151 0.011429
R25504 vdd.n882 vdd.n829 0.0114143
R25505 vdd.n2114 vdd.n1948 0.0113992
R25506 vdd.n2134 vdd.n1961 0.0113992
R25507 vdd.n1805 vdd.n441 0.0113992
R25508 vdd.n2973 vdd 0.0113592
R25509 vdd.n1702 vdd.n1701 0.0112239
R25510 vdd.n935 vdd.n934 0.0111549
R25511 vdd.n2757 vdd.n2692 0.0110874
R25512 vdd.n2751 vdd.n73 0.0110874
R25513 vdd.n2108 vdd.n1944 0.0110586
R25514 vdd.n2140 vdd.n1962 0.0110586
R25515 vdd.n1812 vdd.n438 0.0110586
R25516 vdd.n822 vdd.n821 0.0110546
R25517 vdd.n897 vdd.n816 0.0110025
R25518 vdd.n1671 vdd.n507 0.0108887
R25519 vdd.n1773 vdd.n1737 0.0108791
R25520 vdd.n2284 vdd.n1934 0.0108791
R25521 vdd.n2785 vdd.n2670 0.0107459
R25522 vdd.n2723 vdd.n83 0.0107459
R25523 vdd.n2826 vdd.n125 0.0107459
R25524 vdd.n2083 vdd.n1930 0.010718
R25525 vdd.n1837 vdd.n410 0.010718
R25526 vdd.n1454 vdd.n1453 0.0106562
R25527 vdd.n924 vdd.n725 0.0106407
R25528 vdd.n796 vdd.n717 0.0106351
R25529 vdd.n923 vdd.n922 0.0105906
R25530 vdd.n1637 vdd.n1636 0.0105536
R25531 vdd.n1707 vdd.n470 0.0105536
R25532 vdd.n2343 vdd.n2342 0.0104398
R25533 vdd.n1134 vdd.n967 0.0104278
R25534 vdd.n1544 vdd.n585 0.0104278
R25535 vdd.n1690 vdd.n493 0.0104278
R25536 vdd.n2546 vdd.n14 0.0104044
R25537 vdd.n2644 vdd.n154 0.0104044
R25538 vdd.n2722 vdd.n84 0.0104044
R25539 vdd.n2841 vdd.n93 0.0104044
R25540 vdd.n1916 vdd.n333 0.0103774
R25541 vdd.n1862 vdd.n382 0.0103774
R25542 vdd.n887 vdd.n826 0.0102268
R25543 vdd.n1029 vdd.n953 0.0102185
R25544 vdd.n886 vdd.n885 0.0101788
R25545 vdd vdd.n2973 0.010141
R25546 vdd.n2576 vdd.n24 0.0100628
R25547 vdd.n2619 vdd.n186 0.0100628
R25548 vdd.n2779 vdd.n2778 0.0100628
R25549 vdd.n870 vdd.n844 0.00998661
R25550 vdd.n1751 vdd.n370 0.00997653
R25551 vdd.n2262 vdd.n1964 0.00997653
R25552 vdd.n1011 vdd.n970 0.00988338
R25553 vdd.n1590 vdd.n1589 0.00988338
R25554 vdd.n1235 vdd.n1234 0.009875
R25555 vdd.n1293 vdd.n623 0.009875
R25556 vdd.n892 vdd.n819 0.00981291
R25557 vdd.n894 vdd.n893 0.00976689
R25558 vdd.n2594 vdd.n209 0.00972131
R25559 vdd.n2603 vdd.n34 0.00972131
R25560 vdd.n986 vdd.n985 0.00954826
R25561 vdd.n591 vdd.n590 0.00954826
R25562 vdd.n925 vdd.n724 0.00939901
R25563 vdd.n927 vdd.n926 0.0093968
R25564 vdd.n902 vdd.n749 0.0093968
R25565 vdd.n823 vdd.n749 0.0093968
R25566 vdd.n848 vdd.n837 0.0093968
R25567 vdd.n2525 vdd.n2524 0.00937978
R25568 vdd.n2600 vdd.n206 0.00937978
R25569 vdd.n2628 vdd.n44 0.00937978
R25570 vdd.n348 vdd.n345 0.00935559
R25571 vdd.n755 vdd.n726 0.00935502
R25572 vdd.n1109 vdd.n982 0.00921314
R25573 vdd.n579 vdd.n570 0.00921314
R25574 vdd.n2554 vdd.n2553 0.00903825
R25575 vdd.n2803 vdd.n54 0.00903825
R25576 vdd.n2832 vdd.n90 0.00903825
R25577 vdd.n2067 vdd.n1919 0.00901499
R25578 vdd.n1853 vdd.n388 0.00901499
R25579 vdd.n888 vdd.n820 0.0089851
R25580 vdd.n828 vdd.n827 0.00894316
R25581 vdd.n2223 vdd.n2212 0.0089359
R25582 vdd.n1079 vdd.n965 0.00887802
R25583 vdd.n1597 vdd.n535 0.00887802
R25584 vdd.n855 vdd.n852 0.00887054
R25585 vdd.n798 vdd.n796 0.00881601
R25586 vdd.n186 vdd.n182 0.00869672
R25587 vdd.n2767 vdd.n2766 0.00869672
R25588 vdd.n752 vdd.n749 0.00869672
R25589 vdd.n896 vdd.n749 0.00869672
R25590 vdd.n2092 vdd.n1932 0.00867439
R25591 vdd.n2156 vdd.n1974 0.00867439
R25592 vdd.n1828 vdd.n416 0.00867439
R25593 vdd.n2209 vdd.n2178 0.00863461
R25594 vdd.n2225 vdd.n2214 0.00863461
R25595 vdd.n891 vdd.n820 0.00857119
R25596 vdd.n1052 vdd.n951 0.0085429
R25597 vdd.n827 vdd.n818 0.0085313
R25598 vdd.n2774 vdd.n64 0.00835519
R25599 vdd.n2856 vdd.n2855 0.00835519
R25600 vdd.n2117 vdd.n1949 0.00833379
R25601 vdd.n2131 vdd.n1960 0.00833379
R25602 vdd.n1802 vdd.n444 0.00833379
R25603 vdd.n2211 vdd.n2176 0.00833333
R25604 vdd.n2211 vdd.n2210 0.00833333
R25605 vdd.n2232 vdd.n2231 0.00833333
R25606 vdd.n2440 vdd.n2439 0.0083125
R25607 vdd.n934 vdd.n712 0.00829626
R25608 vdd.n793 vdd.n724 0.00815728
R25609 vdd.n900 vdd.n750 0.00815728
R25610 vdd.n861 vdd.n860 0.00815728
R25611 vdd.n2184 vdd.n2178 0.00803205
R25612 vdd.n2225 vdd.n2224 0.00803205
R25613 vdd.n2760 vdd.n70 0.00801366
R25614 vdd.n2748 vdd.n74 0.00801366
R25615 vdd.n2723 vdd.n2722 0.00801366
R25616 vdd.n2105 vdd.n1943 0.00799319
R25617 vdd.n2143 vdd.n1966 0.00799319
R25618 vdd.n1815 vdd.n435 0.00799319
R25619 vdd.n508 vdd.n504 0.00787265
R25620 vdd.n1698 vdd.n488 0.00787265
R25621 vdd.n778 vdd.n766 0.00785802
R25622 vdd.n771 vdd.n766 0.00785802
R25623 vdd vdd.n2972 0.00779603
R25624 vdd.n799 vdd.n793 0.00777651
R25625 vdd.n892 vdd.n891 0.00774338
R25626 vdd.n2206 vdd.n2205 0.00773077
R25627 vdd.n2230 vdd.n2212 0.00773077
R25628 vdd.n2289 vdd.n1929 0.00772022
R25629 vdd.n893 vdd.n818 0.00770758
R25630 vdd.n2778 vdd.n64 0.00767213
R25631 vdd.n2734 vdd.n80 0.00767213
R25632 vdd.n2817 vdd.n84 0.00767213
R25633 vdd.n2080 vdd.n2037 0.00765259
R25634 vdd.n1840 vdd.n407 0.00765259
R25635 vdd.n475 vdd.n474 0.00753753
R25636 vdd.n1169 vdd.n686 0.00753125
R25637 vdd.n1198 vdd.n671 0.00753125
R25638 vdd.n1227 vdd.n656 0.00753125
R25639 vdd.n1257 vdd.n641 0.00753125
R25640 vdd.n1286 vdd.n626 0.00753125
R25641 vdd.n1480 vdd.n1304 0.00753125
R25642 vdd.n1452 vdd.n1320 0.00753125
R25643 vdd.n1426 vdd.n1425 0.00753125
R25644 vdd.n1401 vdd.n1400 0.00753125
R25645 vdd.n1375 vdd.n305 0.00753125
R25646 vdd.n2366 vdd.n287 0.00753125
R25647 vdd.n2398 vdd.n275 0.00753125
R25648 vdd.n2431 vdd.n263 0.00753125
R25649 vdd.n2463 vdd.n251 0.00753125
R25650 vdd.n1464 vdd.n1463 0.00753125
R25651 vdd.n2541 vdd.n15 0.0073306
R25652 vdd.n2622 vdd.n182 0.0073306
R25653 vdd.n2641 vdd.n50 0.0073306
R25654 vdd.n2846 vdd.n94 0.0073306
R25655 vdd.n888 vdd.n887 0.00732947
R25656 vdd.n886 vdd.n828 0.00729572
R25657 vdd.n928 vdd.n927 0.00728295
R25658 vdd.n1129 vdd.n973 0.00726895
R25659 vdd.n1541 vdd.n588 0.00726895
R25660 vdd.n1779 vdd.n1778 0.00726895
R25661 vdd.n1027 vdd.n957 0.00720241
R25662 vdd.n367 vdd.n342 0.00712651
R25663 vdd.n2581 vdd.n25 0.00698907
R25664 vdd.n2616 vdd.n40 0.00698907
R25665 vdd.n529 vdd.n517 0.0069759
R25666 vdd.n1295 vdd.n524 0.0069759
R25667 vdd.n2308 vdd.n2307 0.00697139
R25668 vdd.n1865 vdd.n378 0.00697139
R25669 vdd.n925 vdd.n924 0.00691556
R25670 vdd.n923 vdd.n726 0.00688385
R25671 vdd.n1009 vdd.n971 0.00686729
R25672 vdd.n1584 vdd.n1583 0.00686729
R25673 vdd.n1703 vdd.n480 0.00681769
R25674 vdd.n1911 vdd.n1910 0.00681769
R25675 vdd.n1244 vdd.n1243 0.00675
R25676 vdd.n1283 vdd.n628 0.00675
R25677 vdd.n529 vdd.n515 0.0066747
R25678 vdd.n1500 vdd.n1297 0.0066747
R25679 vdd.n2339 vdd.n303 0.0066747
R25680 vdd.n2546 vdd.n2545 0.00664754
R25681 vdd.n2591 vdd.n30 0.00664754
R25682 vdd.n2606 vdd.n35 0.00664754
R25683 vdd.n863 vdd.n848 0.00663839
R25684 vdd.n1524 vdd.n1523 0.00653217
R25685 vdd.n1540 vdd.n589 0.00653217
R25686 vdd.n1896 vdd.n342 0.0065241
R25687 vdd.n821 vdd.n819 0.00650166
R25688 vdd.n894 vdd.n816 0.00647199
R25689 vdd.n1297 vdd.n1295 0.00637349
R25690 vdd.n2342 vdd.n303 0.00637349
R25691 vdd.n2257 vdd.n1970 0.00636643
R25692 vdd.n2530 vdd.n20 0.00630601
R25693 vdd.n215 vdd.n29 0.00630601
R25694 vdd.n2631 vdd.n45 0.00630601
R25695 vdd.n2318 vdd.n315 0.00629019
R25696 vdd.n787 vdd.n722 0.00621726
R25697 vdd.n1103 vdd.n981 0.00619705
R25698 vdd.n1559 vdd.n1558 0.00619705
R25699 vdd.n833 vdd.n826 0.00608775
R25700 vdd.n885 vdd.n829 0.00606013
R25701 vdd.n1188 vdd.n674 0.00596875
R25702 vdd.n1217 vdd.n659 0.00596875
R25703 vdd.n1247 vdd.n644 0.00596875
R25704 vdd.n1276 vdd.n629 0.00596875
R25705 vdd.n1486 vdd.n1299 0.00596875
R25706 vdd.n1458 vdd.n1318 0.00596875
R25707 vdd.n1430 vdd.n1334 0.00596875
R25708 vdd.n1406 vdd.n1405 0.00596875
R25709 vdd.n1381 vdd.n1380 0.00596875
R25710 vdd.n2355 vdd.n289 0.00596875
R25711 vdd.n2387 vdd.n277 0.00596875
R25712 vdd.n2420 vdd.n265 0.00596875
R25713 vdd.n2452 vdd.n253 0.00596875
R25714 vdd.n793 vdd.n722 0.00595738
R25715 vdd.n789 vdd.n715 0.00595738
R25716 vdd.n2070 vdd.n2047 0.00594959
R25717 vdd.n1850 vdd.n391 0.00594959
R25718 vdd.n1076 vdd.n964 0.00586193
R25719 vdd.n761 vdd.n757 0.00569751
R25720 vdd.n731 vdd.n725 0.00567384
R25721 vdd.n922 vdd.n727 0.00564827
R25722 vdd.n2557 vdd.n10 0.00562295
R25723 vdd.n2800 vdd.n55 0.00562295
R25724 vdd.n2829 vdd.n89 0.00562295
R25725 vdd.n1904 vdd.n342 0.00560899
R25726 vdd.n2095 vdd.n1936 0.00560899
R25727 vdd.n2153 vdd.n1973 0.00560899
R25728 vdd.n1825 vdd.n419 0.00560899
R25729 vdd.n1647 vdd.n532 0.00552681
R25730 vdd.n2570 vdd.n234 0.00528142
R25731 vdd.n2771 vdd.n65 0.00528142
R25732 vdd.n2707 vdd.n2705 0.00528142
R25733 vdd.n2738 vdd.n79 0.00528142
R25734 vdd.n2121 vdd.n1950 0.00526839
R25735 vdd.n2128 vdd.n1956 0.00526839
R25736 vdd.n1799 vdd.n447 0.00526839
R25737 vdd.n822 vdd.n750 0.00525993
R25738 vdd.n898 vdd.n897 0.00523641
R25739 vdd.n1151 vdd.n1150 0.00519169
R25740 vdd.n2450 vdd.n2449 0.0051875
R25741 vdd.n2185 vdd.n2184 0.00516987
R25742 vdd.n2224 vdd.n0 0.00516987
R25743 vdd.n2789 vdd.n60 0.00493989
R25744 vdd.n2763 vdd.n69 0.00493989
R25745 vdd.n2745 vdd.n75 0.00493989
R25746 vdd.n2102 vdd.n1942 0.00492779
R25747 vdd.n2146 vdd.n1967 0.00492779
R25748 vdd.n1818 vdd.n428 0.00492779
R25749 vdd.n505 vdd.n502 0.00485657
R25750 vdd.n1695 vdd.n1694 0.00485657
R25751 vdd.n880 vdd.n834 0.00484603
R25752 vdd.n882 vdd.n881 0.00482455
R25753 vdd.n901 vdd.n900 0.00463907
R25754 vdd.n900 vdd.n753 0.00461862
R25755 vdd.n900 vdd.n899 0.00461862
R25756 vdd.n2490 vdd.n2489 0.00459836
R25757 vdd.n2793 vdd.n59 0.00459836
R25758 vdd.n2820 vdd.n85 0.00459836
R25759 vdd.n2209 vdd.n2208 0.00456731
R25760 vdd.n2228 vdd.n2214 0.00456731
R25761 vdd.n945 vdd.n944 0.00452145
R25762 vdd.n1723 vdd.n1722 0.00452145
R25763 vdd.n917 vdd.n732 0.00443212
R25764 vdd.n919 vdd.n918 0.00441269
R25765 vdd.n851 vdd.n688 0.00440625
R25766 vdd.n1473 vdd.n1472 0.00440625
R25767 vdd.n2198 vdd.n2186 0.00431088
R25768 vdd.n2200 vdd.n2198 0.00431088
R25769 vdd.n2538 vdd.n2514 0.00425683
R25770 vdd.n2638 vdd.n49 0.00425683
R25771 vdd.n2850 vdd.n95 0.00425683
R25772 vdd.n2077 vdd.n1925 0.00424659
R25773 vdd.n1843 vdd.n400 0.00424659
R25774 vdd.n1025 vdd.n958 0.00418633
R25775 vdd.n1785 vdd.n1784 0.00411011
R25776 vdd.n2295 vdd.n2294 0.00411011
R25777 vdd.n901 vdd.n747 0.00401821
R25778 vdd.n753 vdd.n751 0.00400082
R25779 vdd.n899 vdd.n898 0.00400082
R25780 vdd.n2584 vdd.n221 0.0039153
R25781 vdd.n206 vdd.n33 0.0039153
R25782 vdd.n2613 vdd.n39 0.0039153
R25783 vdd.n2835 vdd.n117 0.0039153
R25784 vdd.n2846 vdd.n2845 0.0039153
R25785 vdd.n2311 vdd.n329 0.00390599
R25786 vdd.n1868 vdd.n371 0.00390599
R25787 vdd.n804 vdd.n803 0.00387838
R25788 vdd.n1007 vdd.n975 0.00385121
R25789 vdd.n1580 vdd.n559 0.00385121
R25790 vdd.n2973 vdd.n0 0.00366346
R25791 vdd.n1124 vdd.n979 0.00365884
R25792 vdd.n1526 vdd.n594 0.00365884
R25793 vdd.n1726 vdd.n1725 0.00365884
R25794 vdd.n2306 vdd.n336 0.00365884
R25795 vdd.n1255 vdd.n1254 0.003625
R25796 vdd.n1273 vdd.n633 0.003625
R25797 vdd.n879 vdd.n835 0.0036043
R25798 vdd.n839 vdd.n832 0.00358896
R25799 vdd.n2588 vdd.n29 0.00357377
R25800 vdd.n162 vdd.n49 0.00357377
R25801 vdd.n1520 vdd.n603 0.00351609
R25802 vdd.n1533 vdd.n593 0.00351609
R25803 vdd.n1660 vdd.n517 0.00351205
R25804 vdd.n1896 vdd.n1895 0.00351205
R25805 vdd.n814 vdd.n754 0.00338303
R25806 vdd.n2231 vdd.n2175 0.00336218
R25807 vdd.n2790 vdd.n2789 0.00323224
R25808 vdd.n2315 vdd.n318 0.0032248
R25809 vdd.n1899 vdd.n358 0.0032248
R25810 vdd.n2252 vdd.n1975 0.00320758
R25811 vdd.n916 vdd.n733 0.0031904
R25812 vdd.n1100 vdd.n977 0.00318097
R25813 vdd.n737 vdd.n730 0.0031771
R25814 vdd.n768 vdd.n767 0.00316393
R25815 vdd.n2533 vdd.n19 0.00289071
R25816 vdd.n173 vdd.n167 0.00289071
R25817 vdd.n2697 vdd.n73 0.00289071
R25818 vdd.n2856 vdd.n2854 0.00289071
R25819 vdd.n2044 vdd.n1922 0.0028842
R25820 vdd.n1847 vdd.n394 0.0028842
R25821 vdd.n1571 vdd.n1570 0.00284584
R25822 vdd.n905 vdd.n904 0.00277649
R25823 vdd.n762 vdd.n761 0.00276524
R25824 vdd.n906 vdd.n743 0.00276524
R25825 vdd.n862 vdd.n861 0.00273214
R25826 vdd.n2493 vdd.n9 0.00254918
R25827 vdd.n2581 vdd.n2580 0.00254918
R25828 vdd.n200 vdd.n192 0.00254918
R25829 vdd.n2658 vdd.n2656 0.00254918
R25830 vdd.n2797 vdd.n2658 0.00254918
R25831 vdd.n2826 vdd.n88 0.00254918
R25832 vdd.n2022 vdd.n1937 0.0025436
R25833 vdd.n2150 vdd.n1972 0.0025436
R25834 vdd.n1822 vdd.n422 0.0025436
R25835 vdd.n1073 vdd.n963 0.00251072
R25836 vdd.n1656 vdd.n527 0.00251072
R25837 vdd.n876 vdd.n875 0.00236258
R25838 vdd.n761 vdd.n754 0.00235338
R25839 vdd.n874 vdd.n840 0.00235338
R25840 vdd.n1641 vdd.n1640 0.00230723
R25841 vdd.n1886 vdd.n351 0.00230723
R25842 vdd.n2768 vdd.n2679 0.00220765
R25843 vdd.n2741 vdd.n78 0.00220765
R25844 vdd.n2003 vdd.n1954 0.002203
R25845 vdd.n2125 vdd.n1955 0.002203
R25846 vdd.n1796 vdd.n450 0.002203
R25847 vdd.n2233 vdd.n2232 0.00219675
R25848 vdd.n1154 vdd.n699 0.0021756
R25849 vdd.n1793 vdd.n1792 0.0021756
R25850 vdd.n2462 vdd.n2461 0.0020625
R25851 vdd.n2471 vdd.n2470 0.0020625
R25852 vdd.n767 vdd.n765 0.00195349
R25853 vdd.n913 vdd.n912 0.00194868
R25854 vdd.n911 vdd.n738 0.00194152
R25855 vdd.n2766 vdd.n68 0.00186612
R25856 vdd.n2742 vdd.n2707 0.00186612
R25857 vdd.n1681 vdd.n499 0.00184048
R25858 vdd.n1689 vdd.n1688 0.00184048
R25859 vdd.n2200 vdd.n2199 0.00170513
R25860 vdd.n811 vdd.n757 0.0015395
R25861 vdd.n807 vdd.n782 0.0015395
R25862 vdd.n746 vdd.n745 0.00153477
R25863 vdd.n907 vdd.n742 0.00152965
R25864 vdd.n2561 vdd.n8 0.00152459
R25865 vdd.n201 vdd.n200 0.00152459
R25866 vdd.n2796 vdd.n58 0.00152459
R25867 vdd.n2823 vdd.n128 0.00152459
R25868 vdd.n2099 vdd.n1938 0.0015218
R25869 vdd.n1983 vdd.n1968 0.0015218
R25870 vdd.n431 vdd.n425 0.0015218
R25871 vdd.n1158 vdd.n692 0.00150536
R25872 vdd.n1719 vdd.n467 0.00150536
R25873 vdd.n773 vdd.n770 0.00132372
R25874 vdd.n1166 vdd.n1165 0.00128125
R25875 vdd.n1194 vdd.n1193 0.00128125
R25876 vdd.n1223 vdd.n1222 0.00128125
R25877 vdd.n1253 vdd.n1252 0.00128125
R25878 vdd.n1282 vdd.n1281 0.00128125
R25879 vdd.n1485 vdd.n1484 0.00128125
R25880 vdd.n1457 vdd.n1456 0.00128125
R25881 vdd.n1429 vdd.n1336 0.00128125
R25882 vdd.n1357 vdd.n1355 0.00128125
R25883 vdd.n1377 vdd.n1376 0.00128125
R25884 vdd.n2361 vdd.n2360 0.00128125
R25885 vdd.n2393 vdd.n2392 0.00128125
R25886 vdd.n2426 vdd.n2425 0.00128125
R25887 vdd.n2458 vdd.n2457 0.00128125
R25888 vdd.n1482 vdd.n1481 0.00128125
R25889 vdd.n2554 vdd.n2502 0.00118306
R25890 vdd.n2535 vdd.n18 0.00118306
R25891 vdd.n2635 vdd.n48 0.00118306
R25892 vdd.n151 vdd.n53 0.00118306
R25893 vdd.n2735 vdd.n2734 0.00118306
R25894 vdd.n107 vdd.n98 0.00118306
R25895 vdd.n2074 vdd.n1924 0.0011812
R25896 vdd.n405 vdd.n397 0.0011812
R25897 vdd.n1023 vdd.n959 0.00117024
R25898 vdd.n1297 vdd.n621 0.00113542
R25899 vdd.n1659 vdd.n1658 0.00113542
R25900 vdd.n1653 vdd.n517 0.00113542
R25901 vdd.n1634 vdd.n1620 0.00113542
R25902 vdd.n1640 vdd.n1639 0.00113542
R25903 vdd.n356 vdd.n297 0.00113542
R25904 vdd.n1897 vdd.n1896 0.00113542
R25905 vdd.n366 vdd.n365 0.00113542
R25906 vdd.n1901 vdd.n351 0.00113542
R25907 vdd.n860 vdd.n838 0.00112086
R25908 vdd.n873 vdd.n841 0.00111779
R25909 vdd.n303 vdd.n295 0.00111306
R25910 vdd.n2206 vdd.n2177 0.00110256
R25911 vdd.n2229 vdd.n2213 0.00110256
R25912 vdd.n1620 vdd.n515 0.00110241
R25913 vdd.n367 vdd.n366 0.00110241
R25914 vdd.n2301 vdd.n2300 0.000951264
R25915 vdd.n218 vdd.n28 0.00084153
R25916 vdd.n2610 vdd.n38 0.00084153
R25917 vdd.n2314 vdd.n325 0.000840599
R25918 vdd.n1869 vdd.n353 0.000840599
R25919 vdd.n944 vdd.n943 0.000835121
R25920 vdd.n1158 vdd.n1157 0.000835121
R25921 vdd.n1154 vdd.n694 0.000835121
R25922 vdd.n1151 vdd.n701 0.000835121
R25923 vdd.n1052 vdd.n703 0.000835121
R25924 vdd.n1055 vdd.n1050 0.000835121
R25925 vdd.n1058 vdd.n1031 0.000835121
R25926 vdd.n1061 vdd.n1029 0.000835121
R25927 vdd.n1064 vdd.n1027 0.000835121
R25928 vdd.n1067 vdd.n1025 0.000835121
R25929 vdd.n1070 vdd.n1023 0.000835121
R25930 vdd.n1073 vdd.n1021 0.000835121
R25931 vdd.n1076 vdd.n1019 0.000835121
R25932 vdd.n1079 vdd.n1017 0.000835121
R25933 vdd.n1082 vdd.n1015 0.000835121
R25934 vdd.n1085 vdd.n1013 0.000835121
R25935 vdd.n1088 vdd.n1011 0.000835121
R25936 vdd.n1091 vdd.n1009 0.000835121
R25937 vdd.n1094 vdd.n1007 0.000835121
R25938 vdd.n1005 vdd.n976 0.000835121
R25939 vdd.n1097 vdd.n1005 0.000835121
R25940 vdd.n1100 vdd.n1003 0.000835121
R25941 vdd.n1103 vdd.n1000 0.000835121
R25942 vdd.n1110 vdd.n1109 0.000835121
R25943 vdd.n1113 vdd.n984 0.000835121
R25944 vdd.n1116 vdd.n987 0.000835121
R25945 vdd.n985 vdd.n599 0.000835121
R25946 vdd.n1523 vdd.n600 0.000835121
R25947 vdd.n1520 vdd.n1519 0.000835121
R25948 vdd.n610 vdd.n596 0.000835121
R25949 vdd.n595 vdd.n593 0.000835121
R25950 vdd.n1534 vdd.n589 0.000835121
R25951 vdd.n1539 vdd.n591 0.000835121
R25952 vdd.n1549 vdd.n581 0.000835121
R25953 vdd.n1552 vdd.n577 0.000835121
R25954 vdd.n1557 vdd.n570 0.000835121
R25955 vdd.n1559 vdd.n567 0.000835121
R25956 vdd.n1570 vdd.n568 0.000835121
R25957 vdd.n1577 vdd.n561 0.000835121
R25958 vdd.n1577 vdd.n1576 0.000835121
R25959 vdd.n1580 vdd.n557 0.000835121
R25960 vdd.n1583 vdd.n554 0.000835121
R25961 vdd.n1590 vdd.n548 0.000835121
R25962 vdd.n1593 vdd.n544 0.000835121
R25963 vdd.n1596 vdd.n541 0.000835121
R25964 vdd.n1648 vdd.n535 0.000835121
R25965 vdd.n1651 vdd.n532 0.000835121
R25966 vdd.n1656 vdd.n1655 0.000835121
R25967 vdd.n1637 vdd.n1633 0.000835121
R25968 vdd.n1672 vdd.n510 0.000835121
R25969 vdd.n1675 vdd.n507 0.000835121
R25970 vdd.n1678 vdd.n504 0.000835121
R25971 vdd.n1682 vdd.n502 0.000835121
R25972 vdd.n1685 vdd.n499 0.000835121
R25973 vdd.n1688 vdd.n496 0.000835121
R25974 vdd.n1695 vdd.n490 0.000835121
R25975 vdd.n1698 vdd.n486 0.000835121
R25976 vdd.n1701 vdd.n483 0.000835121
R25977 vdd.n1708 vdd.n477 0.000835121
R25978 vdd.n1713 vdd.n470 0.000835121
R25979 vdd.n474 vdd.n463 0.000835121
R25980 vdd.n1722 vdd.n464 0.000835121
R25981 vdd.n1719 vdd.n1718 0.000835121
R25982 vdd.n1793 vdd.n456 0.000835121
R25983 vdd.n2202 vdd.n2183 0.000791375
R25984 vdd.n811 vdd.n810 0.000759875
R25985 vdd.n807 vdd.n759 0.000759875
R25986 vdd.n804 vdd.n784 0.000759875
R25987 vdd.n802 vdd.n787 0.000759875
R25988 vdd.n799 vdd.n798 0.000759875
R25989 vdd.n935 vdd.n717 0.000759875
R25990 vdd.n939 vdd.n712 0.000759875
R25991 vdd.n789 vdd.n709 0.000759875
R25992 vdd.n744 vdd.n736 0.000706954
R25993 vdd.n910 vdd.n739 0.000705931
R25994 a_10611_n7515.n1 a_10611_n7515.t1 126.15
R25995 a_10611_n7515.n0 a_10611_n7515.t2 126.094
R25996 a_10611_n7515.n1 a_10611_n7515.t3 126.037
R25997 a_10611_n7515.n0 a_10611_n7515.t0 126.037
R25998 a_10611_n7515.n0 a_10611_n7515.t4 126.037
R25999 a_10611_n7515.t5 a_10611_n7515.n1 126.037
R26000 a_10611_n7515.t10 a_10611_n7515.n0 0.59297
R26001 a_10611_n7515.n4 a_10611_n7515.n2 0.214595
R26002 a_10611_n7515.n3 a_10611_n7515.t8 0.348901
R26003 a_10611_n7515.n4 a_10611_n7515.n3 0.686012
R26004 a_10611_n7515.t10 a_10611_n7515.n4 0.645791
R26005 a_10611_n7515.t10 a_10611_n7515.t7 0.568679
R26006 a_10611_n7515.n3 a_10611_n7515.t11 0.350693
R26007 a_10611_n7515.n2 a_10611_n7515.t9 0.357917
R26008 a_10611_n7515.n2 a_10611_n7515.t6 0.341402
R26009 a_10611_n7515.n1 a_10611_n7515.n0 0.317717
C0 vin_n vin_p 0.125714f
C1 vdd vin_p 0.022884f
C2 iref vout 15.642901f
C3 vdd vout 0.123081p
C4 iref vin_n 0.089257f
C5 vdd vin_n 0.086828f
C6 vdd iref 49.5943f
C7 vin_p vss 11.341963f
C8 vout vss 0.210875p
C9 vin_n vss 11.22703f
C10 iref vss 13.256209f
C11 vdd vss 0.147511p
C12 a_10611_n7515.t10 vss 31.115902f
C13 a_10611_n7515.n0 vss 1.10718f
C14 a_10611_n7515.n1 vss 0.338734f
C15 a_10611_n7515.n2 vss 3.97193f
C16 a_10611_n7515.n3 vss 5.32214f
C17 a_10611_n7515.n4 vss 4.22076f
C18 a_10611_n7515.t6 vss 25.5957f
C19 a_10611_n7515.t8 vss 25.6346f
C20 a_10611_n7515.t11 vss 25.6492f
C21 a_10611_n7515.t9 vss 25.6853f
C22 a_10611_n7515.t7 vss 25.656599f
C23 a_10611_n7515.t2 vss 0.017022f
C24 a_10611_n7515.t4 vss 0.01699f
C25 a_10611_n7515.t0 vss 0.01699f
C26 a_10611_n7515.t1 vss 0.017073f
C27 a_10611_n7515.t3 vss 0.01699f
C28 a_10611_n7515.t5 vss 0.01699f
C29 vdd.n0 vss 0.017558f
C30 vdd.n1 vss 0.048562f
C31 vdd.n2 vss 0.062653f
C32 vdd.n3 vss 0.062653f
C33 vdd.n4 vss 0.048562f
C34 vdd.n5 vss 0.048176f
C35 vdd.n6 vss 0.048562f
C36 vdd.n7 vss 0.048562f
C37 vdd.n8 vss 0.028519f
C38 vdd.n9 vss 0.028519f
C39 vdd.n10 vss 0.027727f
C40 vdd.n11 vss 0.048863f
C41 vdd.n12 vss 0.048562f
C42 vdd.n13 vss 0.028519f
C43 vdd.n14 vss 0.028519f
C44 vdd.n15 vss 0.021389f
C45 vdd.n16 vss 0.048562f
C46 vdd.n17 vss 0.048863f
C47 vdd.n18 vss 0.028519f
C48 vdd.n19 vss 0.028519f
C49 vdd.n20 vss 0.028519f
C50 vdd.n21 vss 0.048562f
C51 vdd.n22 vss 0.048562f
C52 vdd.n23 vss 0.028519f
C53 vdd.n24 vss 0.028519f
C54 vdd.n25 vss 0.028519f
C55 vdd.n26 vss 0.048562f
C56 vdd.n27 vss 0.048863f
C57 vdd.n28 vss 0.028519f
C58 vdd.n29 vss 0.010299f
C59 vdd.n30 vss 0.028519f
C60 vdd.n31 vss 0.048562f
C61 vdd.n32 vss 0.048562f
C62 vdd.n33 vss 0.018221f
C63 vdd.n34 vss 0.028519f
C64 vdd.n35 vss 0.028519f
C65 vdd.n36 vss 0.048863f
C66 vdd.n37 vss 0.048562f
C67 vdd.n38 vss 0.028519f
C68 vdd.n39 vss 0.028519f
C69 vdd.n40 vss 0.028519f
C70 vdd.n41 vss 0.048562f
C71 vdd.n42 vss 0.048562f
C72 vdd.n43 vss 0.028519f
C73 vdd.n44 vss 0.028519f
C74 vdd.n45 vss 0.028519f
C75 vdd.n46 vss 0.048863f
C76 vdd.n47 vss 0.048562f
C77 vdd.n48 vss 0.028519f
C78 vdd.n49 vss 0.007922f
C79 vdd.n50 vss 0.028519f
C80 vdd.n51 vss 0.048562f
C81 vdd.n52 vss 0.048863f
C82 vdd.n53 vss 0.015844f
C83 vdd.n54 vss 0.028519f
C84 vdd.n55 vss 0.028519f
C85 vdd.n56 vss 0.048562f
C86 vdd.n57 vss 0.048562f
C87 vdd.n58 vss 0.028519f
C88 vdd.n59 vss 0.028519f
C89 vdd.n60 vss 0.02535f
C90 vdd.n61 vss 0.048562f
C91 vdd.n62 vss 0.048863f
C92 vdd.n63 vss 0.028519f
C93 vdd.n64 vss 0.017428f
C94 vdd.n65 vss 0.028519f
C95 vdd.n66 vss 0.048562f
C96 vdd.n67 vss 0.048562f
C97 vdd.n68 vss 0.028519f
C98 vdd.n69 vss 0.028519f
C99 vdd.n70 vss 0.028519f
C100 vdd.n71 vss 0.048863f
C101 vdd.n72 vss 0.048562f
C102 vdd.n73 vss 0.015052f
C103 vdd.n74 vss 0.028519f
C104 vdd.n75 vss 0.028519f
C105 vdd.n76 vss 0.048562f
C106 vdd.n77 vss 0.048562f
C107 vdd.n78 vss 0.028519f
C108 vdd.n79 vss 0.028519f
C109 vdd.n80 vss 0.027727f
C110 vdd.n81 vss 0.048863f
C111 vdd.n82 vss 0.048562f
C112 vdd.n83 vss 0.028519f
C113 vdd.n84 vss 0.019805f
C114 vdd.n85 vss 0.028519f
C115 vdd.n86 vss 0.048562f
C116 vdd.n87 vss 0.048863f
C117 vdd.n88 vss 0.028519f
C118 vdd.n89 vss 0.028519f
C119 vdd.n90 vss 0.024558f
C120 vdd.n91 vss 0.048562f
C121 vdd.n92 vss 0.048562f
C122 vdd.n93 vss 0.028519f
C123 vdd.n94 vss 0.028519f
C124 vdd.n95 vss 0.024558f
C125 vdd.n96 vss 0.048562f
C126 vdd.n97 vss 0.722237f
C127 vdd.n98 vss 0.029311f
C128 vdd.n99 vss 0.006445f
C129 vdd.n100 vss 0.005299f
C130 vdd.n101 vss 0.006445f
C131 vdd.n102 vss 0.005299f
C132 vdd.n103 vss 0.005299f
C133 vdd.n104 vss 0.005299f
C134 vdd.n105 vss 0.005299f
C135 vdd.n106 vss 0.005299f
C136 vdd.n107 vss 0.028519f
C137 vdd.n108 vss 0.005299f
C138 vdd.n109 vss 0.005299f
C139 vdd.n110 vss 0.005299f
C140 vdd.n111 vss 0.005299f
C141 vdd.n112 vss 0.005299f
C142 vdd.n113 vss 0.028519f
C143 vdd.n114 vss 0.005299f
C144 vdd.n115 vss 0.005299f
C145 vdd.t286 vss 0.018831f
C146 vdd.t113 vss 0.018831f
C147 vdd.n116 vss 0.039834f
C148 vdd.n117 vss 0.133772f
C149 vdd.n118 vss 0.005299f
C150 vdd.n119 vss 0.005299f
C151 vdd.n120 vss 0.005299f
C152 vdd.n121 vss 0.005299f
C153 vdd.n122 vss 0.005299f
C154 vdd.n123 vss 0.005299f
C155 vdd.t194 vss 0.018831f
C156 vdd.t71 vss 0.018831f
C157 vdd.n124 vss 0.039834f
C158 vdd.n125 vss 0.143675f
C159 vdd.n126 vss 0.005299f
C160 vdd.n127 vss 0.004967f
C161 vdd.n128 vss 0.028519f
C162 vdd.n129 vss 0.005299f
C163 vdd.n130 vss 0.005299f
C164 vdd.n131 vss 0.005299f
C165 vdd.n132 vss 0.005299f
C166 vdd.n133 vss 0.005299f
C167 vdd.n134 vss 0.005299f
C168 vdd.n135 vss 0.09004f
C169 vdd.n136 vss 0.459657f
C170 vdd.t160 vss 0.337394f
C171 vdd.t138 vss 0.463521f
C172 vdd.t252 vss 0.337394f
C173 vdd.t248 vss 0.337394f
C174 vdd.t112 vss 0.337394f
C175 vdd.t285 vss 0.337394f
C176 vdd.t70 vss 0.337394f
C177 vdd.t193 vss 0.337394f
C178 vdd.n137 vss 0.09004f
C179 vdd.n138 vss 0.033043f
C180 vdd.n139 vss 0.09004f
C181 vdd.n140 vss 0.09004f
C182 vdd.n141 vss -0.498418f
C183 vdd.t14 vss 0.337394f
C184 vdd.t10 vss 0.337394f
C185 vdd.t126 vss 0.337394f
C186 vdd.t241 vss 0.337394f
C187 vdd.t2 vss 0.337394f
C188 vdd.t181 vss 0.416023f
C189 vdd.n142 vss 0.033043f
C190 vdd.n143 vss 0.494652f
C191 vdd.t20 vss 0.416023f
C192 vdd.t136 vss 0.337394f
C193 vdd.t130 vss 0.337394f
C194 vdd.t76 vss 0.337394f
C195 vdd.t198 vss 0.337394f
C196 vdd.t283 vss 0.337394f
C197 vdd.t68 vss 0.337394f
C198 vdd.n144 vss 0.09004f
C199 vdd.n145 vss 0.003643f
C200 vdd.n146 vss 0.005299f
C201 vdd.n147 vss 0.005299f
C202 vdd.n148 vss 0.005299f
C203 vdd.n149 vss -0.221586f
C204 vdd.t5 vss 0.018831f
C205 vdd.t192 vss 0.018831f
C206 vdd.n150 vss 0.039834f
C207 vdd.n151 vss 0.128623f
C208 vdd.n152 vss 0.004121f
C209 vdd.n153 vss 0.005299f
C210 vdd.n154 vss 0.028519f
C211 vdd.n155 vss -0.21879f
C212 vdd.n156 vss 0.003827f
C213 vdd.n157 vss 0.005299f
C214 vdd.n158 vss 0.005299f
C215 vdd.n159 vss 0.005299f
C216 vdd.n160 vss 0.005299f
C217 vdd.t224 vss 0.018831f
C218 vdd.t247 vss 0.018831f
C219 vdd.n161 vss 0.039834f
C220 vdd.n162 vss 0.139318f
C221 vdd.n163 vss 0.005299f
C222 vdd.n164 vss 0.005299f
C223 vdd.n165 vss 0.005299f
C224 vdd.n166 vss 0.005299f
C225 vdd.n167 vss 0.031292f
C226 vdd.n168 vss 0.005299f
C227 vdd.n169 vss 0.005299f
C228 vdd.t123 vss 0.018831f
C229 vdd.t9 vss 0.018831f
C230 vdd.n170 vss 0.039834f
C231 vdd.n171 vss 0.005299f
C232 vdd.n172 vss 0.005299f
C233 vdd.n173 vss 0.028519f
C234 vdd.n174 vss 0.005299f
C235 vdd.n175 vss 0.005299f
C236 vdd.n176 vss 0.005299f
C237 vdd.n177 vss 0.005299f
C238 vdd.n178 vss 0.005299f
C239 vdd.n179 vss 0.005299f
C240 vdd.n180 vss 0.005299f
C241 vdd.t184 vss 0.018831f
C242 vdd.t289 vss 0.018831f
C243 vdd.n181 vss 0.039834f
C244 vdd.n182 vss 0.132584f
C245 vdd.n183 vss 0.005299f
C246 vdd.n184 vss 0.005299f
C247 vdd.n185 vss 0.005299f
C248 vdd.n186 vss 0.020597f
C249 vdd.n187 vss 0.005299f
C250 vdd.n188 vss 0.005299f
C251 vdd.n189 vss 0.019171f
C252 vdd.n190 vss 0.005299f
C253 vdd.n191 vss 0.005299f
C254 vdd.n192 vss 0.030896f
C255 vdd.n193 vss 0.005299f
C256 vdd.n194 vss 0.003974f
C257 vdd.n195 vss 0.005299f
C258 vdd.n196 vss 0.005299f
C259 vdd.n197 vss 0.005299f
C260 vdd.n198 vss 0.005299f
C261 vdd.n199 vss 0.005299f
C262 vdd.t255 vss 0.070922f
C263 vdd.n200 vss 0.125294f
C264 vdd.n201 vss 0.026143f
C265 vdd.n202 vss 0.005299f
C266 vdd.n203 vss 0.005299f
C267 vdd.n204 vss 0.005299f
C268 vdd.t117 vss 0.018831f
C269 vdd.t19 vss 0.018831f
C270 vdd.n205 vss 0.039834f
C271 vdd.n206 vss 0.129415f
C272 vdd.n207 vss 0.005299f
C273 vdd.n208 vss 0.005299f
C274 vdd.n209 vss 0.028519f
C275 vdd.n210 vss 0.005299f
C276 vdd.n211 vss 0.005299f
C277 vdd.n212 vss 0.005299f
C278 vdd.n213 vss 0.005299f
C279 vdd.t75 vss 0.018831f
C280 vdd.t294 vss 0.018831f
C281 vdd.n214 vss 0.039834f
C282 vdd.n215 vss 0.14011f
C283 vdd.n216 vss 0.005299f
C284 vdd.n217 vss 0.005299f
C285 vdd.n218 vss 0.028915f
C286 vdd.n219 vss 0.005299f
C287 vdd.n220 vss 0.005299f
C288 vdd.n221 vss 0.026143f
C289 vdd.n222 vss 0.005299f
C290 vdd.n223 vss 0.005299f
C291 vdd.n224 vss 0.005299f
C292 vdd.n225 vss 0.005299f
C293 vdd.n226 vss 0.005299f
C294 vdd.n227 vss 0.005299f
C295 vdd.n228 vss 0.003643f
C296 vdd.n229 vss 0.005299f
C297 vdd.n230 vss 0.005299f
C298 vdd.n231 vss 0.005299f
C299 vdd.n232 vss 0.005299f
C300 vdd.t186 vss 0.018831f
C301 vdd.t165 vss 0.018831f
C302 vdd.n233 vss 0.039834f
C303 vdd.n234 vss 0.133376f
C304 vdd.n235 vss 0.005299f
C305 vdd.n236 vss 0.005299f
C306 vdd.n237 vss 0.108288f
C307 vdd.t118 vss 0.679306f
C308 vdd.n238 vss 0.181626f
C309 vdd.n239 vss 0.181626f
C310 vdd.n240 vss 0.038356f
C311 vdd.n241 vss 0.005299f
C312 vdd.n242 vss 0.013853f
C313 vdd.t119 vss 0.072462f
C314 vdd.n243 vss 0.027705f
C315 vdd.n244 vss 0.012467f
C316 vdd.n245 vss 0.005299f
C317 vdd.n246 vss 0.013853f
C318 vdd.t313 vss 0.018831f
C319 vdd.t233 vss 0.018831f
C320 vdd.n247 vss 0.041538f
C321 vdd.n248 vss 0.027359f
C322 vdd.n249 vss 0.012467f
C323 vdd.n250 vss 0.005299f
C324 vdd.n251 vss 0.013853f
C325 vdd.n252 vss 0.026666f
C326 vdd.n253 vss 0.013679f
C327 vdd.n254 vss 0.005299f
C328 vdd.n255 vss 0.013853f
C329 vdd.n256 vss 0.025974f
C330 vdd.n257 vss 0.012467f
C331 vdd.n258 vss 0.005299f
C332 vdd.n259 vss 0.013853f
C333 vdd.n260 vss 0.025281f
C334 vdd.n261 vss 0.012467f
C335 vdd.n262 vss 0.005299f
C336 vdd.n263 vss 0.013853f
C337 vdd.n264 vss 0.024588f
C338 vdd.n265 vss 0.013679f
C339 vdd.n266 vss 0.002649f
C340 vdd.n267 vss 0.013853f
C341 vdd.n268 vss 0.023896f
C342 vdd.n269 vss 0.012467f
C343 vdd.n270 vss 0.005299f
C344 vdd.n271 vss 0.013853f
C345 vdd.n272 vss 0.023203f
C346 vdd.n273 vss 0.012467f
C347 vdd.n274 vss 0.005299f
C348 vdd.n275 vss 0.013853f
C349 vdd.n276 vss 0.022511f
C350 vdd.n277 vss 0.013679f
C351 vdd.n278 vss 0.005299f
C352 vdd.n279 vss 0.013853f
C353 vdd.n280 vss 0.021818f
C354 vdd.n281 vss 0.012467f
C355 vdd.n282 vss 0.005299f
C356 vdd.n283 vss 0.013853f
C357 vdd.n284 vss 0.021125f
C358 vdd.n285 vss 0.012467f
C359 vdd.n286 vss 0.005299f
C360 vdd.n287 vss 0.013853f
C361 vdd.n288 vss 0.020433f
C362 vdd.n289 vss 0.013679f
C363 vdd.n290 vss 0.005299f
C364 vdd.n291 vss 0.013853f
C365 vdd.n292 vss 0.027705f
C366 vdd.n293 vss 0.012467f
C367 vdd.n294 vss 0.063804f
C368 vdd.n295 vss 0.055418f
C369 vdd.n296 vss 0.011197f
C370 vdd.n297 vss 2.09024f
C371 vdd.n298 vss 0.027705f
C372 vdd.n299 vss 0.027705f
C373 vdd.n300 vss 0.027705f
C374 vdd.n301 vss 0.027705f
C375 vdd.n302 vss 0.013853f
C376 vdd.n303 vss 0.071861f
C377 vdd.n304 vss 0.022337f
C378 vdd.n305 vss 0.012467f
C379 vdd.n306 vss 0.005299f
C380 vdd.n307 vss 0.034552f
C381 vdd.n308 vss 0.181626f
C382 vdd.n309 vss 0.181626f
C383 vdd.t110 vss 0.679306f
C384 vdd.n310 vss -0.21879f
C385 vdd.t232 vss 0.550915f
C386 vdd.t108 vss 0.550915f
C387 vdd.t201 vss 0.550915f
C388 vdd.t44 vss 0.550915f
C389 vdd.t56 vss 0.550915f
C390 vdd.t162 vss 0.550915f
C391 vdd.t38 vss 0.550915f
C392 vdd.t52 vss 0.550915f
C393 vdd.t100 vss 0.550915f
C394 vdd.t114 vss 0.550915f
C395 vdd.t230 vss 0.550915f
C396 vdd.t96 vss 0.550915f
C397 vdd.t90 vss 0.550915f
C398 vdd.t187 vss 0.550915f
C399 vdd.t48 vss 0.550915f
C400 vdd.t158 vss 0.550915f
C401 vdd.t30 vss 0.550915f
C402 vdd.t42 vss 0.550915f
C403 vdd.t0 vss 0.550915f
C404 vdd.t104 vss 0.550915f
C405 vdd.t98 vss 0.550915f
C406 vdd.t218 vss 0.550915f
C407 vdd.t78 vss 0.550915f
C408 vdd.t175 vss 0.413185f
C409 vdd.n311 vss 0.44733f
C410 vdd.n312 vss 0.450127f
C411 vdd.n313 vss 0.003827f
C412 vdd.n314 vss 0.005299f
C413 vdd.n315 vss 0.028595f
C414 vdd.n316 vss 0.004121f
C415 vdd.n317 vss 0.005299f
C416 vdd.n318 vss 0.028597f
C417 vdd.n319 vss 0.002649f
C418 vdd.n320 vss 0.005299f
C419 vdd.n321 vss 0.005299f
C420 vdd.n322 vss 0.005299f
C421 vdd.n323 vss 0.005299f
C422 vdd.n324 vss 0.005299f
C423 vdd.n325 vss 0.028595f
C424 vdd.n326 vss 0.005299f
C425 vdd.n327 vss 0.005299f
C426 vdd.n328 vss 0.005299f
C427 vdd.n329 vss 0.028597f
C428 vdd.n330 vss 0.005299f
C429 vdd.n331 vss 0.005299f
C430 vdd.n332 vss 0.005299f
C431 vdd.n333 vss 0.032567f
C432 vdd.n334 vss 0.048562f
C433 vdd.t295 vss 0.018831f
C434 vdd.t209 vss 0.018831f
C435 vdd.n335 vss 0.042405f
C436 vdd.n336 vss 0.238925f
C437 vdd.n337 vss 0.048562f
C438 vdd.t271 vss 0.018831f
C439 vdd.t79 vss 0.018831f
C440 vdd.n338 vss 0.042405f
C441 vdd.n339 vss 0.048562f
C442 vdd.n340 vss 0.048863f
C443 vdd.n341 vss 0.048863f
C444 vdd.n342 vss 0.100475f
C445 vdd.n343 vss 0.00673f
C446 vdd.n344 vss 0.003017f
C447 vdd.n345 vss 0.028597f
C448 vdd.n346 vss 0.003827f
C449 vdd.n347 vss 0.005299f
C450 vdd.n348 vss 0.032171f
C451 vdd.n349 vss 0.003827f
C452 vdd.n350 vss 0.00673f
C453 vdd.n351 vss 0.089826f
C454 vdd.n352 vss 0.005299f
C455 vdd.n353 vss 0.028993f
C456 vdd.n354 vss 0.006739f
C457 vdd.n355 vss 0.036071f
C458 vdd.n356 vss 0.060256f
C459 vdd.n357 vss 0.004789f
C460 vdd.n358 vss 0.022242f
C461 vdd.n359 vss 0.005299f
C462 vdd.n364 vss 0.048562f
C463 vdd.n365 vss 0.060712f
C464 vdd.n366 vss 0.08264f
C465 vdd.n367 vss 0.043116f
C466 vdd.n369 vss 0.048562f
C467 vdd.t217 vss 0.073257f
C468 vdd.n370 vss 0.245436f
C469 vdd.n371 vss 0.028597f
C470 vdd.n372 vss 0.005299f
C471 vdd.n373 vss 0.005299f
C472 vdd.n374 vss 0.0046f
C473 vdd.n375 vss 0.005299f
C474 vdd.n376 vss 0.005299f
C475 vdd.n377 vss 0.005299f
C476 vdd.n378 vss 0.028595f
C477 vdd.n379 vss 0.005299f
C478 vdd.n380 vss 0.005299f
C479 vdd.n381 vss 0.005299f
C480 vdd.n382 vss 0.028595f
C481 vdd.n383 vss 0.005299f
C482 vdd.n384 vss 0.005299f
C483 vdd.n385 vss 0.028597f
C484 vdd.n386 vss 0.005299f
C485 vdd.n387 vss 0.005299f
C486 vdd.n388 vss 0.028595f
C487 vdd.n389 vss 0.005299f
C488 vdd.n390 vss 0.005299f
C489 vdd.n391 vss 0.028597f
C490 vdd.n392 vss 0.005299f
C491 vdd.n393 vss 0.005299f
C492 vdd.n394 vss 0.028595f
C493 vdd.n395 vss 0.005299f
C494 vdd.n396 vss 0.005299f
C495 vdd.n397 vss 0.029391f
C496 vdd.n398 vss 0.005299f
C497 vdd.n399 vss 0.005299f
C498 vdd.n400 vss 0.028595f
C499 vdd.n401 vss 0.005299f
C500 vdd.n402 vss 0.005299f
C501 vdd.n403 vss 0.005299f
C502 vdd.n404 vss 0.005299f
C503 vdd.n405 vss 0.028597f
C504 vdd.n406 vss 0.005299f
C505 vdd.n407 vss 0.028595f
C506 vdd.n408 vss 0.005299f
C507 vdd.n409 vss 0.005299f
C508 vdd.n410 vss 0.028597f
C509 vdd.n411 vss 0.005299f
C510 vdd.n412 vss 0.005299f
C511 vdd.n413 vss 0.028595f
C512 vdd.n414 vss 0.005299f
C513 vdd.n415 vss 0.005299f
C514 vdd.n416 vss 0.028597f
C515 vdd.n417 vss 0.005299f
C516 vdd.n418 vss 0.005299f
C517 vdd.n419 vss 0.028595f
C518 vdd.n420 vss 0.005299f
C519 vdd.n421 vss 0.005299f
C520 vdd.n422 vss 0.028597f
C521 vdd.n423 vss 0.005299f
C522 vdd.n424 vss 0.005299f
C523 vdd.n425 vss 0.029788f
C524 vdd.n426 vss 0.005299f
C525 vdd.n427 vss 0.005299f
C526 vdd.n428 vss 0.028595f
C527 vdd.n429 vss 0.005299f
C528 vdd.n430 vss 0.005299f
C529 vdd.n431 vss 0.028595f
C530 vdd.n432 vss 0.005299f
C531 vdd.n433 vss 0.005299f
C532 vdd.n434 vss 0.005299f
C533 vdd.n435 vss 0.028597f
C534 vdd.n436 vss 0.005299f
C535 vdd.n437 vss 0.005299f
C536 vdd.n438 vss 0.028595f
C537 vdd.n439 vss 0.005299f
C538 vdd.n440 vss 0.005299f
C539 vdd.n441 vss 0.028597f
C540 vdd.n442 vss 0.005299f
C541 vdd.n443 vss 0.005299f
C542 vdd.n444 vss 0.028595f
C543 vdd.n445 vss 0.005299f
C544 vdd.n446 vss 0.005299f
C545 vdd.n447 vss 0.028597f
C546 vdd.n448 vss 0.005299f
C547 vdd.n449 vss 0.008684f
C548 vdd.n450 vss 0.028595f
C549 vdd.n451 vss 0.005299f
C550 vdd.n452 vss 0.008647f
C551 vdd.n453 vss 0.063781f
C552 vdd.n454 vss 0.008647f
C553 vdd.n455 vss 0.005299f
C554 vdd.n456 vss 0.029062f
C555 vdd.n457 vss 0.008647f
C556 vdd.n458 vss 0.046465f
C557 vdd.t251 vss 0.018831f
C558 vdd.t135 vss 0.018831f
C559 vdd.n459 vss 0.042405f
C560 vdd.n460 vss 0.263208f
C561 vdd.n461 vss 0.048562f
C562 vdd.n462 vss 0.048562f
C563 vdd.n463 vss 0.024218f
C564 vdd.n464 vss 0.027853f
C565 vdd.n465 vss 0.005299f
C566 vdd.n466 vss 0.008684f
C567 vdd.n467 vss 0.02866f
C568 vdd.n468 vss 0.005299f
C569 vdd.n469 vss 0.005299f
C570 vdd.n470 vss 0.012513f
C571 vdd.n471 vss 0.005299f
C572 vdd.n472 vss 0.005299f
C573 vdd.n473 vss 0.005299f
C574 vdd.n474 vss 0.008879f
C575 vdd.n475 vss 0.02866f
C576 vdd.n476 vss 0.005299f
C577 vdd.n477 vss 0.016145f
C578 vdd.n478 vss 0.005299f
C579 vdd.t67 vss 0.018831f
C580 vdd.t311 vss 0.018831f
C581 vdd.n479 vss 0.042405f
C582 vdd.n480 vss 0.238626f
C583 vdd.n481 vss 0.048863f
C584 vdd.n482 vss 0.048863f
C585 vdd.n483 vss 0.020182f
C586 vdd.n484 vss 0.005299f
C587 vdd.n485 vss 0.005299f
C588 vdd.n486 vss 0.023816f
C589 vdd.n487 vss 0.005299f
C590 vdd.n488 vss 0.02866f
C591 vdd.n489 vss 0.005299f
C592 vdd.n490 vss 0.027448f
C593 vdd.n491 vss 0.005299f
C594 vdd.t280 vss 0.018831f
C595 vdd.t190 vss 0.018831f
C596 vdd.n492 vss 0.042405f
C597 vdd.n493 vss 0.238626f
C598 vdd.n494 vss 0.048562f
C599 vdd.n495 vss 0.048562f
C600 vdd.n496 vss 0.029062f
C601 vdd.n497 vss 0.005299f
C602 vdd.n498 vss 0.005299f
C603 vdd.n499 vss 0.002017f
C604 vdd.n500 vss 0.005299f
C605 vdd.n501 vss 0.005299f
C606 vdd.n502 vss 0.005649f
C607 vdd.n503 vss 0.005299f
C608 vdd.n504 vss 0.009283f
C609 vdd.n505 vss 0.02866f
C610 vdd.n506 vss 0.005299f
C611 vdd.n507 vss 0.012915f
C612 vdd.n508 vss 0.02866f
C613 vdd.n509 vss 0.00673f
C614 vdd.n510 vss 0.016952f
C615 vdd.n511 vss 0.005299f
C616 vdd.n512 vss 0.048863f
C617 vdd.n513 vss 0.032974f
C618 vdd.n514 vss 0.048562f
C619 vdd.n515 vss 0.040422f
C620 vdd.n517 vss 0.05659f
C621 vdd.n518 vss 0.048562f
C622 vdd.n524 vss 2.13652f
C623 vdd.n525 vss 0.036061f
C624 vdd.n526 vss 0.034552f
C625 vdd.n527 vss 0.02866f
C626 vdd.n528 vss 0.006739f
C627 vdd.n529 vss 0.117838f
C628 vdd.n530 vss 0.006739f
C629 vdd.n531 vss 0.005299f
C630 vdd.n532 vss 0.006457f
C631 vdd.n533 vss 0.005299f
C632 vdd.n534 vss 0.005299f
C633 vdd.n535 vss 0.010493f
C634 vdd.n536 vss 0.005299f
C635 vdd.t148 vss 0.073257f
C636 vdd.n537 vss 0.245735f
C637 vdd.n538 vss 0.048562f
C638 vdd.n539 vss 0.048562f
C639 vdd.n540 vss 0.048562f
C640 vdd.n541 vss 0.014128f
C641 vdd.n542 vss 0.005299f
C642 vdd.n543 vss 0.005299f
C643 vdd.n544 vss 0.01776f
C644 vdd.n545 vss 0.005299f
C645 vdd.n546 vss 0.02866f
C646 vdd.n547 vss 0.005299f
C647 vdd.n548 vss 0.021394f
C648 vdd.n549 vss 0.005299f
C649 vdd.t93 vss 0.018831f
C650 vdd.t7 vss 0.018831f
C651 vdd.n550 vss 0.042405f
C652 vdd.n551 vss 0.238626f
C653 vdd.n552 vss 0.048562f
C654 vdd.n553 vss 0.048562f
C655 vdd.n554 vss 0.025026f
C656 vdd.n555 vss 0.005299f
C657 vdd.n556 vss 0.005299f
C658 vdd.n557 vss 0.02866f
C659 vdd.n558 vss 0.005299f
C660 vdd.n559 vss 0.02866f
C661 vdd.n560 vss 0.005299f
C662 vdd.n561 vss 0.029062f
C663 vdd.n562 vss 0.005299f
C664 vdd.t298 vss 0.018831f
C665 vdd.t212 vss 0.018831f
C666 vdd.n563 vss 0.042405f
C667 vdd.n564 vss 0.238626f
C668 vdd.n565 vss 0.048863f
C669 vdd.n566 vss 0.048863f
C670 vdd.n567 vss 0.026238f
C671 vdd.n568 vss 0.029062f
C672 vdd.n569 vss 0.005299f
C673 vdd.n570 vss 0.010898f
C674 vdd.n571 vss 0.005299f
C675 vdd.n572 vss 0.005299f
C676 vdd.n573 vss 0.005299f
C677 vdd.n574 vss 0.005299f
C678 vdd.n575 vss 0.005299f
C679 vdd.n576 vss 0.004121f
C680 vdd.n577 vss 0.01453f
C681 vdd.n578 vss 0.005299f
C682 vdd.n579 vss 0.02866f
C683 vdd.n580 vss -0.21879f
C684 vdd.n581 vss 0.018164f
C685 vdd.n582 vss 0.004121f
C686 vdd.n583 vss 0.048562f
C687 vdd.t272 vss 0.018831f
C688 vdd.t85 vss 0.018831f
C689 vdd.n584 vss 0.042405f
C690 vdd.n585 vss 0.238626f
C691 vdd.n586 vss 0.048562f
C692 vdd.t257 vss 0.018831f
C693 vdd.t144 vss 0.018831f
C694 vdd.n587 vss 0.042405f
C695 vdd.n588 vss 0.238626f
C696 vdd.n589 vss 0.007669f
C697 vdd.n590 vss 0.02866f
C698 vdd.n591 vss 0.011301f
C699 vdd.n592 vss 0.005299f
C700 vdd.n593 vss 0.004035f
C701 vdd.n594 vss 0.026679f
C702 vdd.n595 vss 0.029062f
C703 vdd.n596 vss 0.029062f
C704 vdd.n597 vss 0.048562f
C705 vdd.n598 vss 0.048562f
C706 vdd.n599 vss 0.021796f
C707 vdd.n600 vss 0.02543f
C708 vdd.n601 vss 0.005299f
C709 vdd.n602 vss 0.005299f
C710 vdd.n603 vss 0.02866f
C711 vdd.n604 vss 0.002649f
C712 vdd.n605 vss 0.003827f
C713 vdd.n606 vss 0.005299f
C714 vdd.n607 vss 0.005299f
C715 vdd.n608 vss 0.005299f
C716 vdd.n609 vss 0.005299f
C717 vdd.n610 vss 0.029062f
C718 vdd.n611 vss 0.003827f
C719 vdd.n612 vss 0.005299f
C720 vdd.n613 vss 0.005299f
C721 vdd.n614 vss 0.005299f
C722 vdd.n615 vss 0.005299f
C723 vdd.n616 vss 0.005299f
C724 vdd.t40 vss 0.373502f
C725 vdd.t228 vss 0.550915f
C726 vdd.t64 vss 0.550915f
C727 vdd.t60 vss 0.550915f
C728 vdd.t179 vss 0.550915f
C729 vdd.t46 vss 0.550915f
C730 vdd.t155 vss 0.550915f
C731 vdd.t26 vss 0.550915f
C732 vdd.t120 vss 0.550915f
C733 vdd.t239 vss 0.550915f
C734 vdd.t102 vss 0.550915f
C735 vdd.t221 vss 0.550915f
C736 vdd.t215 vss 0.550915f
C737 vdd.t58 vss 0.550915f
C738 vdd.t172 vss 0.550915f
C739 vdd.t34 vss 0.550915f
C740 vdd.t149 vss 0.550915f
C741 vdd.t16 vss 0.550915f
C742 vdd.t28 vss 0.550915f
C743 vdd.t237 vss 0.550915f
C744 vdd.t66 vss 0.550915f
C745 vdd.t86 vss 0.550915f
C746 vdd.t207 vss 0.550915f
C747 vdd.t62 vss 0.550915f
C748 vdd.t167 vss 0.679306f
C749 vdd.n617 vss 2.60984f
C750 vdd.n618 vss 0.181626f
C751 vdd.n619 vss 0.181626f
C752 vdd.n620 vss 0.004673f
C753 vdd.n621 vss 0.060349f
C754 vdd.n622 vss 0.012467f
C755 vdd.t51 vss 0.072462f
C756 vdd.n623 vss 0.220946f
C757 vdd.n624 vss 0.012467f
C758 vdd.n625 vss 0.005299f
C759 vdd.n626 vss 0.013853f
C760 vdd.t306 vss 0.018831f
C761 vdd.t244 vss 0.018831f
C762 vdd.n627 vss 0.041538f
C763 vdd.n628 vss 0.214207f
C764 vdd.n629 vss 0.013679f
C765 vdd.n630 vss 0.005299f
C766 vdd.n631 vss 0.012467f
C767 vdd.t226 vss 0.018831f
C768 vdd.t107 vss 0.018831f
C769 vdd.n632 vss 0.041538f
C770 vdd.n633 vss 0.214207f
C771 vdd.n634 vss 0.012467f
C772 vdd.n635 vss 0.005299f
C773 vdd.n636 vss 0.013853f
C774 vdd.t178 vss 0.018831f
C775 vdd.t305 vss 0.018831f
C776 vdd.n637 vss 0.041538f
C777 vdd.n638 vss 0.027705f
C778 vdd.n639 vss 0.012467f
C779 vdd.n640 vss 0.005299f
C780 vdd.n641 vss 0.013853f
C781 vdd.t154 vss 0.018831f
C782 vdd.t41 vss 0.018831f
C783 vdd.n642 vss 0.041538f
C784 vdd.n643 vss 0.027705f
C785 vdd.n644 vss 0.013679f
C786 vdd.n645 vss 0.005299f
C787 vdd.n646 vss 0.013853f
C788 vdd.t37 vss 0.018831f
C789 vdd.t261 vss 0.018831f
C790 vdd.n647 vss 0.041538f
C791 vdd.n648 vss 0.027705f
C792 vdd.n649 vss 0.012467f
C793 vdd.n650 vss 0.005299f
C794 vdd.n651 vss 0.013853f
C795 vdd.t302 vss 0.018831f
C796 vdd.t33 vss 0.018831f
C797 vdd.n652 vss 0.041538f
C798 vdd.n653 vss 0.027705f
C799 vdd.n654 vss 0.012467f
C800 vdd.n655 vss 0.005299f
C801 vdd.n656 vss 0.013853f
C802 vdd.t214 vss 0.018831f
C803 vdd.t95 vss 0.018831f
C804 vdd.n657 vss 0.041538f
C805 vdd.n658 vss 0.027705f
C806 vdd.n659 vss 0.013679f
C807 vdd.n660 vss 0.005299f
C808 vdd.n661 vss 0.013853f
C809 vdd.t89 vss 0.018831f
C810 vdd.t300 vss 0.018831f
C811 vdd.n662 vss 0.041538f
C812 vdd.n663 vss 0.027705f
C813 vdd.n664 vss 0.012467f
C814 vdd.n665 vss 0.005299f
C815 vdd.n666 vss 0.013853f
C816 vdd.t147 vss 0.018831f
C817 vdd.t274 vss 0.018831f
C818 vdd.n667 vss 0.041538f
C819 vdd.n668 vss 0.027705f
C820 vdd.n669 vss 0.012467f
C821 vdd.n670 vss 0.005299f
C822 vdd.n671 vss 0.013853f
C823 vdd.t256 vss 0.018831f
C824 vdd.t142 vss 0.018831f
C825 vdd.n672 vss 0.041538f
C826 vdd.n673 vss 0.027705f
C827 vdd.n674 vss 0.013679f
C828 vdd.n675 vss 0.005299f
C829 vdd.n676 vss 0.013853f
C830 vdd.t236 vss 0.018831f
C831 vdd.t23 vss 0.018831f
C832 vdd.n677 vss 0.041538f
C833 vdd.n678 vss 0.027705f
C834 vdd.n679 vss 0.012467f
C835 vdd.n680 vss 0.005299f
C836 vdd.n681 vss 0.013853f
C837 vdd.t206 vss 0.018831f
C838 vdd.t83 vss 0.018831f
C839 vdd.n682 vss 0.041538f
C840 vdd.n683 vss 0.027705f
C841 vdd.n684 vss 0.012467f
C842 vdd.n685 vss 0.003643f
C843 vdd.n686 vss 0.013853f
C844 vdd.n687 vss 0.039322f
C845 vdd.n688 vss 0.019507f
C846 vdd.n689 vss 0.005299f
C847 vdd.n690 vss 0.004268f
C848 vdd.n691 vss 0.005299f
C849 vdd.n692 vss 0.02866f
C850 vdd.n693 vss 0.005299f
C851 vdd.n694 vss 0.029062f
C852 vdd.n695 vss 0.005299f
C853 vdd.n696 vss 0.005299f
C854 vdd.n697 vss 0.005299f
C855 vdd.n698 vss 0.005299f
C856 vdd.n699 vss 0.02866f
C857 vdd.n700 vss 0.005299f
C858 vdd.n701 vss 0.027045f
C859 vdd.n702 vss 0.005299f
C860 vdd.n703 vss 0.023411f
C861 vdd.n704 vss 0.048562f
C862 vdd.t277 vss 0.018831f
C863 vdd.t189 vss 0.018831f
C864 vdd.n705 vss 0.042405f
C865 vdd.n706 vss 0.238925f
C866 vdd.n707 vss 0.048562f
C867 vdd.n708 vss 0.094488f
C868 vdd.n709 vss 0.032115f
C869 vdd.n710 vss 0.005299f
C870 vdd.n711 vss 0.005299f
C871 vdd.n712 vss 0.016136f
C872 vdd.n713 vss 0.005299f
C873 vdd.n714 vss 0.005299f
C874 vdd.n715 vss 0.036958f
C875 vdd.n716 vss 0.005299f
C876 vdd.n717 vss 0.02082f
C877 vdd.n718 vss 0.005299f
C878 vdd.n719 vss 0.075389f
C879 vdd.n720 vss 0.048562f
C880 vdd.n721 vss 0.090466f
C881 vdd.n722 vss 0.022383f
C882 vdd.n723 vss 0.097315f
C883 vdd.n724 vss 0.093267f
C884 vdd.n725 vss 0.048372f
C885 vdd.n726 vss 0.04861f
C886 vdd.n727 vss 0.067066f
C887 vdd.n728 vss 0.249542f
C888 vdd.n729 vss 0.105626f
C889 vdd.n730 vss 0.04861f
C890 vdd.n731 vss 0.093267f
C891 vdd.n732 vss 0.048372f
C892 vdd.n733 vss 0.093267f
C893 vdd.n734 vss 0.097315f
C894 vdd.n735 vss 0.097315f
C895 vdd.n736 vss 0.048372f
C896 vdd.n737 vss 0.067066f
C897 vdd.n738 vss 0.04861f
C898 vdd.n739 vss 0.063783f
C899 vdd.n740 vss 0.105626f
C900 vdd.n741 vss 0.105626f
C901 vdd.n742 vss 0.06641f
C902 vdd.n743 vss 0.04861f
C903 vdd.n744 vss 0.089999f
C904 vdd.n745 vss 0.092614f
C905 vdd.n746 vss 0.048372f
C906 vdd.n747 vss 0.093267f
C907 vdd.n748 vss 0.097315f
C908 vdd.n749 vss 0.101471f
C909 vdd.n750 vss 0.080194f
C910 vdd.n751 vss 0.067066f
C911 vdd.n752 vss 0.07922f
C912 vdd.n753 vss 0.024305f
C913 vdd.n754 vss 0.015108f
C914 vdd.n755 vss 0.162321f
C915 vdd.n756 vss 0.005299f
C916 vdd.n757 vss 0.012493f
C917 vdd.n758 vss 0.006771f
C918 vdd.n759 vss 0.037478f
C919 vdd.n760 vss 0.006771f
C920 vdd.n761 vss 0.023547f
C921 vdd.n762 vss 0.072341f
C922 vdd.n763 vss 0.005299f
C923 vdd.n764 vss 0.005299f
C924 vdd.n765 vss 0.048584f
C925 vdd.n767 vss 0.208662f
C926 vdd.n768 vss 0.077239f
C927 vdd.n770 vss 0.057809f
C928 vdd.n771 vss 0.048562f
C929 vdd.n772 vss 0.051261f
C930 vdd.n773 vss 0.070371f
C931 vdd.n774 vss 0.138587f
C932 vdd.n775 vss 0.117613f
C933 vdd.n777 vss 0.137314f
C934 vdd.n778 vss 0.048562f
C935 vdd.n779 vss 0.048562f
C936 vdd.n780 vss 0.048562f
C937 vdd.n781 vss 0.090466f
C938 vdd.n782 vss 0.036958f
C939 vdd.n783 vss 0.005299f
C940 vdd.n784 vss 0.035396f
C941 vdd.n785 vss 0.005299f
C942 vdd.n786 vss 0.005299f
C943 vdd.n787 vss 0.011972f
C944 vdd.n788 vss 0.005299f
C945 vdd.n789 vss 0.01145f
C946 vdd.n790 vss 0.005299f
C947 vdd.n791 vss 0.005299f
C948 vdd.n792 vss 0.005299f
C949 vdd.n793 vss 0.049692f
C950 vdd.n794 vss 0.005299f
C951 vdd.n795 vss 0.005299f
C952 vdd.n796 vss 0.036958f
C953 vdd.n797 vss 0.005299f
C954 vdd.n798 vss 0.017177f
C955 vdd.n799 vss 0.015095f
C956 vdd.n800 vss 0.005299f
C957 vdd.n801 vss 0.005299f
C958 vdd.n802 vss 0.030712f
C959 vdd.n803 vss 0.036958f
C960 vdd.n804 vss 0.007286f
C961 vdd.n805 vss 0.005299f
C962 vdd.n806 vss 0.005299f
C963 vdd.n807 vss 0.002602f
C964 vdd.n808 vss 0.005299f
C965 vdd.n809 vss 0.006771f
C966 vdd.n810 vss 0.037478f
C967 vdd.n811 vss 0.002602f
C968 vdd.n812 vss 0.006771f
C969 vdd.n813 vss 0.176792f
C970 vdd.n814 vss 0.058591f
C971 vdd.n815 vss 0.251329f
C972 vdd.n816 vss 0.067066f
C973 vdd.n817 vss 0.105626f
C974 vdd.n818 vss 0.04861f
C975 vdd.n819 vss 0.048372f
C976 vdd.n820 vss 0.093267f
C977 vdd.n821 vss 0.093267f
C978 vdd.n822 vss 0.048372f
C979 vdd.n823 vss 0.072986f
C980 vdd.n824 vss 0.097315f
C981 vdd.n825 vss 0.097315f
C982 vdd.n826 vss 0.048372f
C983 vdd.n827 vss 0.067066f
C984 vdd.n828 vss 0.04861f
C985 vdd.n829 vss 0.067066f
C986 vdd.n830 vss 0.105626f
C987 vdd.n831 vss 0.105626f
C988 vdd.n832 vss 0.04861f
C989 vdd.n833 vss 0.093267f
C990 vdd.n834 vss 0.048372f
C991 vdd.n835 vss 0.093267f
C992 vdd.n836 vss 0.097315f
C993 vdd.n837 vss 0.072986f
C994 vdd.n838 vss 0.048372f
C995 vdd.n839 vss 0.067066f
C996 vdd.n840 vss 0.04861f
C997 vdd.n841 vss 0.114364f
C998 vdd.n842 vss 0.105626f
C999 vdd.n843 vss 0.038787f
C1000 vdd.n844 vss 0.014245f
C1001 vdd.n845 vss 0.017454f
C1002 vdd.n846 vss 0.005299f
C1003 vdd.n847 vss 0.019394f
C1004 vdd.n848 vss 0.043722f
C1005 vdd.n849 vss 0.017454f
C1006 vdd.n850 vss 0.005299f
C1007 vdd.n851 vss 0.017454f
C1008 vdd.n852 vss 0.019394f
C1009 vdd.n853 vss 0.036121f
C1010 vdd.n854 vss 0.038787f
C1011 vdd.n855 vss 0.017454f
C1012 vdd.n856 vss 0.019394f
C1013 vdd.n857 vss 0.005299f
C1014 vdd.n858 vss 0.005299f
C1015 vdd.n859 vss 0.018424f
C1016 vdd.n860 vss 0.06712f
C1017 vdd.n861 vss 0.031701f
C1018 vdd.n862 vss 0.010909f
C1019 vdd.n863 vss 0.02206f
C1020 vdd.n864 vss 0.038787f
C1021 vdd.n865 vss 0.017454f
C1022 vdd.n866 vss 0.019394f
C1023 vdd.n867 vss 0.005299f
C1024 vdd.n868 vss 0.006859f
C1025 vdd.n869 vss 0.019394f
C1026 vdd.n870 vss 0.017454f
C1027 vdd.n871 vss 0.198437f
C1028 vdd.n872 vss 0.233623f
C1029 vdd.n873 vss 0.04861f
C1030 vdd.n874 vss 0.067066f
C1031 vdd.n875 vss 0.093267f
C1032 vdd.n876 vss 0.048372f
C1033 vdd.n877 vss 0.097315f
C1034 vdd.n878 vss 0.097315f
C1035 vdd.n879 vss 0.048372f
C1036 vdd.n880 vss 0.093267f
C1037 vdd.n881 vss 0.067066f
C1038 vdd.n882 vss 0.04861f
C1039 vdd.n883 vss 0.105626f
C1040 vdd.n884 vss 0.105626f
C1041 vdd.n885 vss 0.04861f
C1042 vdd.n886 vss 0.067066f
C1043 vdd.n887 vss 0.093267f
C1044 vdd.n888 vss 0.048372f
C1045 vdd.n889 vss 0.097315f
C1046 vdd.n890 vss 0.097315f
C1047 vdd.n891 vss 0.048372f
C1048 vdd.n892 vss 0.093267f
C1049 vdd.n893 vss 0.067066f
C1050 vdd.n894 vss 0.04861f
C1051 vdd.n895 vss 0.105626f
C1052 vdd.n896 vss 0.07922f
C1053 vdd.n897 vss 0.04861f
C1054 vdd.n898 vss 0.040789f
C1055 vdd.n899 vss 0.031115f
C1056 vdd.n900 vss 0.063536f
C1057 vdd.n901 vss 0.024186f
C1058 vdd.n902 vss 0.072986f
C1059 vdd.n903 vss 0.097315f
C1060 vdd.n904 vss 0.048372f
C1061 vdd.n905 vss 0.093267f
C1062 vdd.n906 vss 0.067066f
C1063 vdd.n907 vss 0.04861f
C1064 vdd.n908 vss 0.105626f
C1065 vdd.n909 vss 0.105626f
C1066 vdd.n910 vss 0.04861f
C1067 vdd.n911 vss 0.067066f
C1068 vdd.n912 vss 0.093267f
C1069 vdd.n913 vss 0.048372f
C1070 vdd.n914 vss 0.097315f
C1071 vdd.n915 vss 0.097315f
C1072 vdd.n916 vss 0.048372f
C1073 vdd.n917 vss 0.093267f
C1074 vdd.n918 vss 0.067066f
C1075 vdd.n919 vss 0.04861f
C1076 vdd.n920 vss 0.105626f
C1077 vdd.n921 vss 0.105626f
C1078 vdd.n922 vss 0.04861f
C1079 vdd.n923 vss 0.067066f
C1080 vdd.n924 vss 0.093267f
C1081 vdd.n925 vss 0.048372f
C1082 vdd.n926 vss 0.072986f
C1083 vdd.n927 vss 0.07012f
C1084 vdd.n928 vss 0.060869f
C1085 vdd.n929 vss 0.048863f
C1086 vdd.n930 vss 0.048863f
C1087 vdd.n931 vss 0.048562f
C1088 vdd.n932 vss 0.048562f
C1089 vdd.n933 vss 0.090466f
C1090 vdd.n934 vss 0.036958f
C1091 vdd.n935 vss 0.021861f
C1092 vdd.n936 vss 0.005299f
C1093 vdd.n937 vss 0.005299f
C1094 vdd.n938 vss 0.005299f
C1095 vdd.n939 vss 0.026547f
C1096 vdd.n940 vss 0.005299f
C1097 vdd.n941 vss 0.005299f
C1098 vdd.n942 vss 0.005299f
C1099 vdd.n943 vss 0.027853f
C1100 vdd.n944 vss 0.005247f
C1101 vdd.n945 vss 0.029997f
C1102 vdd.n946 vss 0.055147f
C1103 vdd.n947 vss 0.048562f
C1104 vdd.n948 vss 0.048562f
C1105 vdd.n949 vss 0.048562f
C1106 vdd.n950 vss 0.048562f
C1107 vdd.n951 vss 0.02866f
C1108 vdd.n952 vss 0.02866f
C1109 vdd.n953 vss 0.02866f
C1110 vdd.t309 vss 0.018831f
C1111 vdd.t128 vss 0.018831f
C1112 vdd.n954 vss 0.042405f
C1113 vdd.n955 vss 0.238626f
C1114 vdd.n956 vss 0.048562f
C1115 vdd.n957 vss 0.02866f
C1116 vdd.n958 vss 0.02866f
C1117 vdd.n959 vss 0.02866f
C1118 vdd.t13 vss 0.018831f
C1119 vdd.t245 vss 0.018831f
C1120 vdd.n960 vss 0.042405f
C1121 vdd.n961 vss 0.238626f
C1122 vdd.n962 vss 0.048863f
C1123 vdd.n963 vss 0.02866f
C1124 vdd.n964 vss 0.02866f
C1125 vdd.n965 vss 0.02866f
C1126 vdd.t250 vss 0.018831f
C1127 vdd.t55 vss 0.018831f
C1128 vdd.n966 vss 0.042405f
C1129 vdd.n967 vss 0.238626f
C1130 vdd.n968 vss 0.048562f
C1131 vdd.n969 vss 0.02866f
C1132 vdd.n970 vss 0.02866f
C1133 vdd.n971 vss 0.02866f
C1134 vdd.t195 vss 0.018831f
C1135 vdd.t73 vss 0.018831f
C1136 vdd.n972 vss 0.042405f
C1137 vdd.n973 vss 0.238626f
C1138 vdd.n974 vss 0.048863f
C1139 vdd.n975 vss 0.02866f
C1140 vdd.n976 vss 0.02866f
C1141 vdd.n977 vss 0.02866f
C1142 vdd.t287 vss 0.018831f
C1143 vdd.t200 vss 0.018831f
C1144 vdd.n978 vss 0.042405f
C1145 vdd.n979 vss 0.238626f
C1146 vdd.n980 vss 0.048562f
C1147 vdd.n981 vss 0.02866f
C1148 vdd.n982 vss 0.02866f
C1149 vdd.t81 vss 0.018831f
C1150 vdd.t132 vss 0.018831f
C1151 vdd.n983 vss 0.042405f
C1152 vdd.n984 vss 0.01453f
C1153 vdd.n985 vss 0.011301f
C1154 vdd.n986 vss 0.02866f
C1155 vdd.n987 vss 0.018164f
C1156 vdd.n988 vss 0.005299f
C1157 vdd.n989 vss 0.005299f
C1158 vdd.n990 vss 0.005299f
C1159 vdd.n991 vss 0.005299f
C1160 vdd.n992 vss 0.005299f
C1161 vdd.n993 vss 0.005299f
C1162 vdd.n994 vss 0.005299f
C1163 vdd.n995 vss 0.005299f
C1164 vdd.n996 vss 0.005299f
C1165 vdd.n997 vss 0.005299f
C1166 vdd.n998 vss 0.005299f
C1167 vdd.n999 vss 0.005299f
C1168 vdd.n1000 vss 0.025833f
C1169 vdd.n1001 vss 0.005299f
C1170 vdd.n1002 vss 0.005299f
C1171 vdd.n1003 vss 0.029062f
C1172 vdd.n1004 vss 0.005299f
C1173 vdd.n1005 vss 8.05e-19
C1174 vdd.n1006 vss 0.005299f
C1175 vdd.n1007 vss 0.004439f
C1176 vdd.n1008 vss 0.005299f
C1177 vdd.n1009 vss 0.008071f
C1178 vdd.n1010 vss 0.005299f
C1179 vdd.n1011 vss 0.011706f
C1180 vdd.n1012 vss 0.005299f
C1181 vdd.n1013 vss 0.015337f
C1182 vdd.n1014 vss 0.005299f
C1183 vdd.n1015 vss 0.018972f
C1184 vdd.n1016 vss 0.005299f
C1185 vdd.n1017 vss 0.022604f
C1186 vdd.n1018 vss 0.005299f
C1187 vdd.n1019 vss 0.02664f
C1188 vdd.n1020 vss 0.005299f
C1189 vdd.n1021 vss 0.029062f
C1190 vdd.n1022 vss 0.005299f
C1191 vdd.n1023 vss 0.00121f
C1192 vdd.n1024 vss 0.005299f
C1193 vdd.n1025 vss 0.004842f
C1194 vdd.n1026 vss 0.005299f
C1195 vdd.n1027 vss 0.008476f
C1196 vdd.n1028 vss 0.005299f
C1197 vdd.n1029 vss 0.012108f
C1198 vdd.n1030 vss 0.005299f
C1199 vdd.n1031 vss 0.015742f
C1200 vdd.n1032 vss 0.005299f
C1201 vdd.n1033 vss 0.005299f
C1202 vdd.n1034 vss 0.005299f
C1203 vdd.n1035 vss 0.005299f
C1204 vdd.n1036 vss 0.005299f
C1205 vdd.n1037 vss 0.005299f
C1206 vdd.n1038 vss 0.005299f
C1207 vdd.n1039 vss 0.005299f
C1208 vdd.n1040 vss 0.005299f
C1209 vdd.n1041 vss 0.005299f
C1210 vdd.n1042 vss 0.005299f
C1211 vdd.n1043 vss 0.005299f
C1212 vdd.n1044 vss 0.005299f
C1213 vdd.n1045 vss 0.005299f
C1214 vdd.n1046 vss 0.005299f
C1215 vdd.n1047 vss 0.005299f
C1216 vdd.n1048 vss 0.005299f
C1217 vdd.n1049 vss 0.005299f
C1218 vdd.n1050 vss 0.019374f
C1219 vdd.n1051 vss 0.005299f
C1220 vdd.n1052 vss 0.010091f
C1221 vdd.n1053 vss 0.005299f
C1222 vdd.n1054 vss 0.005299f
C1223 vdd.n1055 vss 0.013723f
C1224 vdd.n1056 vss 0.005299f
C1225 vdd.n1057 vss 0.005299f
C1226 vdd.n1058 vss 0.017357f
C1227 vdd.n1059 vss 0.005299f
C1228 vdd.n1060 vss 0.005299f
C1229 vdd.n1061 vss 0.020989f
C1230 vdd.n1062 vss 0.005299f
C1231 vdd.n1063 vss 0.005299f
C1232 vdd.n1064 vss 0.024623f
C1233 vdd.n1065 vss 0.005299f
C1234 vdd.n1066 vss 0.005299f
C1235 vdd.n1067 vss 0.028255f
C1236 vdd.n1068 vss 0.005299f
C1237 vdd.n1069 vss 0.005299f
C1238 vdd.n1070 vss 0.029062f
C1239 vdd.n1071 vss 0.005299f
C1240 vdd.n1072 vss 0.005299f
C1241 vdd.n1073 vss 0.002825f
C1242 vdd.n1074 vss 0.005299f
C1243 vdd.n1075 vss 0.005299f
C1244 vdd.n1076 vss 0.006861f
C1245 vdd.n1077 vss 0.005299f
C1246 vdd.n1078 vss 0.005299f
C1247 vdd.n1079 vss 0.010493f
C1248 vdd.n1080 vss 0.005299f
C1249 vdd.n1081 vss 0.005299f
C1250 vdd.n1082 vss 0.014128f
C1251 vdd.n1083 vss 0.005299f
C1252 vdd.n1084 vss 0.005299f
C1253 vdd.n1085 vss 0.01776f
C1254 vdd.n1086 vss 0.005299f
C1255 vdd.n1087 vss 0.005299f
C1256 vdd.n1088 vss 0.021394f
C1257 vdd.n1089 vss 0.005299f
C1258 vdd.n1090 vss 0.005299f
C1259 vdd.n1091 vss 0.025026f
C1260 vdd.n1092 vss 0.005299f
C1261 vdd.n1093 vss 0.005299f
C1262 vdd.n1094 vss 0.02866f
C1263 vdd.n1095 vss 0.005299f
C1264 vdd.n1096 vss 0.005299f
C1265 vdd.n1097 vss 0.029062f
C1266 vdd.n1098 vss 0.005299f
C1267 vdd.n1099 vss 0.005299f
C1268 vdd.n1100 vss 0.003632f
C1269 vdd.n1101 vss 0.005299f
C1270 vdd.n1102 vss 0.005299f
C1271 vdd.n1103 vss 0.007264f
C1272 vdd.n1104 vss 0.005299f
C1273 vdd.n1105 vss 0.005299f
C1274 vdd.n1106 vss 0.005299f
C1275 vdd.n1107 vss 0.005299f
C1276 vdd.n1108 vss 0.005299f
C1277 vdd.n1109 vss 0.010898f
C1278 vdd.n1110 vss 0.022201f
C1279 vdd.n1111 vss 0.004452f
C1280 vdd.n1112 vss 0.002649f
C1281 vdd.n1113 vss 0.018567f
C1282 vdd.n1114 vss 0.003496f
C1283 vdd.n1115 vss 0.005299f
C1284 vdd.n1116 vss 0.014935f
C1285 vdd.n1117 vss 0.02866f
C1286 vdd.n1118 vss 0.048562f
C1287 vdd.n1119 vss 0.262908f
C1288 vdd.n1120 vss 0.048562f
C1289 vdd.n1121 vss 0.046465f
C1290 vdd.n1122 vss 0.048562f
C1291 vdd.n1123 vss 0.048863f
C1292 vdd.n1124 vss 0.026679f
C1293 vdd.n1125 vss 0.048863f
C1294 vdd.n1126 vss 0.044067f
C1295 vdd.n1127 vss 0.048562f
C1296 vdd.n1128 vss 0.048562f
C1297 vdd.n1129 vss 0.028777f
C1298 vdd.n1130 vss 0.048562f
C1299 vdd.n1131 vss 0.041967f
C1300 vdd.n1132 vss 0.048562f
C1301 vdd.n1133 vss 0.048562f
C1302 vdd.n1134 vss 0.030876f
C1303 vdd.n1135 vss 0.048863f
C1304 vdd.n1136 vss 0.03987f
C1305 vdd.n1137 vss 0.048863f
C1306 vdd.n1138 vss 0.048562f
C1307 vdd.n1139 vss 0.033275f
C1308 vdd.n1140 vss 0.048562f
C1309 vdd.n1141 vss 0.037471f
C1310 vdd.n1142 vss 0.048562f
C1311 vdd.n1143 vss 0.048562f
C1312 vdd.n1144 vss 0.035372f
C1313 vdd.n1145 vss 0.048562f
C1314 vdd.n1146 vss 0.035372f
C1315 vdd.n1147 vss 0.048863f
C1316 vdd.n1148 vss 0.048863f
C1317 vdd.n1149 vss 0.03777f
C1318 vdd.n1150 vss 0.02866f
C1319 vdd.n1151 vss 0.006054f
C1320 vdd.n1152 vss 0.005299f
C1321 vdd.n1153 vss 0.005299f
C1322 vdd.n1154 vss 0.00242f
C1323 vdd.n1155 vss 0.005299f
C1324 vdd.n1156 vss 0.005299f
C1325 vdd.n1157 vss 0.029062f
C1326 vdd.n1158 vss 0.001613f
C1327 vdd.n1159 vss 0.00368f
C1328 vdd.n1160 vss 0.034552f
C1329 vdd.t153 vss 0.550915f
C1330 vdd.t24 vss 0.550915f
C1331 vdd.t36 vss 0.550915f
C1332 vdd.t32 vss 0.550915f
C1333 vdd.t80 vss 0.550915f
C1334 vdd.t94 vss 0.550915f
C1335 vdd.t213 vss 0.550915f
C1336 vdd.t72 vss 0.550915f
C1337 vdd.t88 vss 0.550915f
C1338 vdd.t54 vss 0.550915f
C1339 vdd.t146 vss 0.550915f
C1340 vdd.t141 vss 0.550915f
C1341 vdd.t12 vss 0.550915f
C1342 vdd.t22 vss 0.550915f
C1343 vdd.t235 vss 0.550915f
C1344 vdd.t82 vss 0.550915f
C1345 vdd.t205 vss 1.09797f
C1346 vdd.n1161 vss 4.32067f
C1347 vdd.n1162 vss 0.063804f
C1348 vdd.n1163 vss 0.034552f
C1349 vdd.n1164 vss 0.004305f
C1350 vdd.n1165 vss 0.012977f
C1351 vdd.n1166 vss 0.012467f
C1352 vdd.n1167 vss 0.028278f
C1353 vdd.n1168 vss 0.027705f
C1354 vdd.n1169 vss 0.012467f
C1355 vdd.n1170 vss 0.013853f
C1356 vdd.n1171 vss 0.005299f
C1357 vdd.n1172 vss 0.005299f
C1358 vdd.n1173 vss 0.013853f
C1359 vdd.n1174 vss 0.012467f
C1360 vdd.n1175 vss 0.020086f
C1361 vdd.n1176 vss 0.214207f
C1362 vdd.n1177 vss 0.021472f
C1363 vdd.n1178 vss 0.012467f
C1364 vdd.n1179 vss 0.013853f
C1365 vdd.n1180 vss 0.005299f
C1366 vdd.n1181 vss 0.005299f
C1367 vdd.n1182 vss 0.013853f
C1368 vdd.n1183 vss 0.012467f
C1369 vdd.n1184 vss 0.019394f
C1370 vdd.n1185 vss 0.214207f
C1371 vdd.n1186 vss 0.022164f
C1372 vdd.n1187 vss 0.012467f
C1373 vdd.n1188 vss 0.012467f
C1374 vdd.n1189 vss 0.013853f
C1375 vdd.n1190 vss 0.005299f
C1376 vdd.n1191 vss 0.005299f
C1377 vdd.n1192 vss 0.005299f
C1378 vdd.n1193 vss 0.012641f
C1379 vdd.n1194 vss 0.012467f
C1380 vdd.n1195 vss 0.018701f
C1381 vdd.n1196 vss 0.214207f
C1382 vdd.n1197 vss 0.022857f
C1383 vdd.n1198 vss 0.012467f
C1384 vdd.n1199 vss 0.013853f
C1385 vdd.n1200 vss 0.005299f
C1386 vdd.n1201 vss 0.005299f
C1387 vdd.n1202 vss 0.013853f
C1388 vdd.n1203 vss 0.012467f
C1389 vdd.n1204 vss 0.018008f
C1390 vdd.n1205 vss 0.214207f
C1391 vdd.n1206 vss 0.023549f
C1392 vdd.n1207 vss 0.012467f
C1393 vdd.n1208 vss 0.013853f
C1394 vdd.n1209 vss 0.005299f
C1395 vdd.n1210 vss 0.005299f
C1396 vdd.n1211 vss 0.013853f
C1397 vdd.n1212 vss 0.012467f
C1398 vdd.n1213 vss 0.017316f
C1399 vdd.n1214 vss 0.214207f
C1400 vdd.n1215 vss 0.024242f
C1401 vdd.n1216 vss 0.012467f
C1402 vdd.n1217 vss 0.012467f
C1403 vdd.n1218 vss 0.013853f
C1404 vdd.n1219 vss 0.005299f
C1405 vdd.n1220 vss 0.005299f
C1406 vdd.n1221 vss 0.005299f
C1407 vdd.n1222 vss 0.012641f
C1408 vdd.n1223 vss 0.012467f
C1409 vdd.n1224 vss 0.016623f
C1410 vdd.n1225 vss 0.214207f
C1411 vdd.n1226 vss 0.024935f
C1412 vdd.n1227 vss 0.012467f
C1413 vdd.n1228 vss 0.013853f
C1414 vdd.n1229 vss 0.004489f
C1415 vdd.n1230 vss 0.002649f
C1416 vdd.n1231 vss 0.003459f
C1417 vdd.n1232 vss 0.013853f
C1418 vdd.n1233 vss 0.012467f
C1419 vdd.n1234 vss 0.01593f
C1420 vdd.n1235 vss 0.214207f
C1421 vdd.n1236 vss 0.025627f
C1422 vdd.n1237 vss 0.012467f
C1423 vdd.n1238 vss 0.013853f
C1424 vdd.n1239 vss 0.005299f
C1425 vdd.n1240 vss 0.005299f
C1426 vdd.n1241 vss 0.013853f
C1427 vdd.n1242 vss 0.012467f
C1428 vdd.n1243 vss 0.015238f
C1429 vdd.n1244 vss 0.214207f
C1430 vdd.n1245 vss 0.02632f
C1431 vdd.n1246 vss 0.012467f
C1432 vdd.n1247 vss 0.012467f
C1433 vdd.n1248 vss 0.013853f
C1434 vdd.n1249 vss 0.005299f
C1435 vdd.n1250 vss 0.005299f
C1436 vdd.n1251 vss 0.005299f
C1437 vdd.n1252 vss 0.012641f
C1438 vdd.n1253 vss 0.012467f
C1439 vdd.n1254 vss 0.014545f
C1440 vdd.n1255 vss 0.214207f
C1441 vdd.n1256 vss 0.027013f
C1442 vdd.n1257 vss 0.012467f
C1443 vdd.n1258 vss 0.013853f
C1444 vdd.n1259 vss 0.005299f
C1445 vdd.n1260 vss 0.005299f
C1446 vdd.n1261 vss 0.013853f
C1447 vdd.n1262 vss 0.012467f
C1448 vdd.n1263 vss 0.22806f
C1449 vdd.n1264 vss 0.027013f
C1450 vdd.n1265 vss 0.027705f
C1451 vdd.n1266 vss 0.012467f
C1452 vdd.n1267 vss 0.013853f
C1453 vdd.n1268 vss 0.005299f
C1454 vdd.n1269 vss 0.005299f
C1455 vdd.n1270 vss 0.013853f
C1456 vdd.n1271 vss 0.013853f
C1457 vdd.n1272 vss 0.012467f
C1458 vdd.n1273 vss 0.014545f
C1459 vdd.n1274 vss 0.027705f
C1460 vdd.n1275 vss 0.02632f
C1461 vdd.n1276 vss 0.012467f
C1462 vdd.n1277 vss 0.013853f
C1463 vdd.n1278 vss 0.005299f
C1464 vdd.n1279 vss 0.005299f
C1465 vdd.n1280 vss 0.005299f
C1466 vdd.n1281 vss 0.012641f
C1467 vdd.n1282 vss 0.012467f
C1468 vdd.n1283 vss 0.015238f
C1469 vdd.n1284 vss 0.025627f
C1470 vdd.n1285 vss 0.027705f
C1471 vdd.n1286 vss 0.012467f
C1472 vdd.n1287 vss 0.013853f
C1473 vdd.n1288 vss 0.005299f
C1474 vdd.n1289 vss 0.005299f
C1475 vdd.n1290 vss 0.013853f
C1476 vdd.n1291 vss 0.013853f
C1477 vdd.n1292 vss 0.012467f
C1478 vdd.n1293 vss 0.01593f
C1479 vdd.n1294 vss 0.027705f
C1480 vdd.n1295 vss 0.073657f
C1481 vdd.n1296 vss 0.027705f
C1482 vdd.n1297 vss 0.071861f
C1483 vdd.n1298 vss 0.027705f
C1484 vdd.n1299 vss 0.012467f
C1485 vdd.n1300 vss 0.182361f
C1486 vdd.n1301 vss 0.063804f
C1487 vdd.n1302 vss 0.036052f
C1488 vdd.n1303 vss 0.005299f
C1489 vdd.n1304 vss 0.013853f
C1490 vdd.t168 vss 0.018831f
C1491 vdd.t296 vss 0.018831f
C1492 vdd.n1305 vss 0.041538f
C1493 vdd.n1306 vss 0.027705f
C1494 vdd.n1307 vss 0.012467f
C1495 vdd.n1308 vss 0.005299f
C1496 vdd.n1309 vss 0.005299f
C1497 vdd.n1310 vss 0.013853f
C1498 vdd.t208 vss 0.018831f
C1499 vdd.t87 vss 0.018831f
C1500 vdd.n1311 vss 0.041538f
C1501 vdd.n1312 vss 0.027705f
C1502 vdd.n1313 vss 0.012467f
C1503 vdd.n1314 vss 0.005299f
C1504 vdd.n1315 vss 0.013853f
C1505 vdd.t299 vss 0.018831f
C1506 vdd.t238 vss 0.018831f
C1507 vdd.n1316 vss 0.041538f
C1508 vdd.n1317 vss 0.027705f
C1509 vdd.n1318 vss 0.012467f
C1510 vdd.n1319 vss 0.005299f
C1511 vdd.n1320 vss 0.013853f
C1512 vdd.t29 vss 0.018831f
C1513 vdd.t259 vss 0.018831f
C1514 vdd.n1321 vss 0.041538f
C1515 vdd.n1322 vss 0.027705f
C1516 vdd.n1323 vss 0.012467f
C1517 vdd.n1324 vss 0.005299f
C1518 vdd.n1325 vss 0.005299f
C1519 vdd.n1326 vss 0.013853f
C1520 vdd.t150 vss 0.018831f
C1521 vdd.t35 vss 0.018831f
C1522 vdd.n1327 vss 0.041538f
C1523 vdd.n1328 vss 0.027705f
C1524 vdd.n1329 vss 0.012467f
C1525 vdd.n1330 vss 0.005299f
C1526 vdd.n1331 vss 0.013853f
C1527 vdd.t173 vss 0.018831f
C1528 vdd.t59 vss 0.018831f
C1529 vdd.n1332 vss 0.041538f
C1530 vdd.n1333 vss 0.027705f
C1531 vdd.n1334 vss 0.012467f
C1532 vdd.n1335 vss 0.002649f
C1533 vdd.n1336 vss 0.012467f
C1534 vdd.n1337 vss 0.005299f
C1535 vdd.n1338 vss 0.013853f
C1536 vdd.t216 vss 0.018831f
C1537 vdd.t222 vss 0.018831f
C1538 vdd.n1339 vss 0.041538f
C1539 vdd.n1340 vss 0.023376f
C1540 vdd.n1341 vss 0.214207f
C1541 vdd.n1342 vss 0.022684f
C1542 vdd.n1343 vss 0.012467f
C1543 vdd.n1344 vss 0.005299f
C1544 vdd.n1345 vss 0.013853f
C1545 vdd.t103 vss 0.018831f
C1546 vdd.t240 vss 0.018831f
C1547 vdd.n1346 vss 0.041538f
C1548 vdd.n1347 vss 0.214207f
C1549 vdd.n1348 vss 0.021991f
C1550 vdd.n1349 vss 0.012467f
C1551 vdd.n1350 vss 0.005299f
C1552 vdd.n1351 vss 0.013853f
C1553 vdd.t121 vss 0.018831f
C1554 vdd.t262 vss 0.018831f
C1555 vdd.n1352 vss 0.041538f
C1556 vdd.n1353 vss 0.214207f
C1557 vdd.n1354 vss 0.021298f
C1558 vdd.n1355 vss 0.012641f
C1559 vdd.n1356 vss 0.005299f
C1560 vdd.n1357 vss 0.012467f
C1561 vdd.n1358 vss 0.013853f
C1562 vdd.t156 vss 0.018831f
C1563 vdd.t47 vss 0.018831f
C1564 vdd.n1359 vss 0.041538f
C1565 vdd.n1360 vss 0.214207f
C1566 vdd.n1361 vss 0.020606f
C1567 vdd.n1362 vss 0.012467f
C1568 vdd.n1363 vss 0.005299f
C1569 vdd.n1364 vss 0.013853f
C1570 vdd.t180 vss 0.018831f
C1571 vdd.t61 vss 0.018831f
C1572 vdd.n1365 vss 0.041538f
C1573 vdd.n1366 vss 0.214207f
C1574 vdd.n1367 vss 0.019913f
C1575 vdd.n1368 vss 0.012467f
C1576 vdd.n1369 vss 0.005299f
C1577 vdd.n1370 vss 0.013853f
C1578 vdd.t65 vss 0.018831f
C1579 vdd.t229 vss 0.018831f
C1580 vdd.n1371 vss 0.041538f
C1581 vdd.n1372 vss 0.214207f
C1582 vdd.t111 vss 0.072462f
C1583 vdd.n1373 vss 0.220946f
C1584 vdd.n1374 vss 0.019221f
C1585 vdd.n1375 vss 0.013853f
C1586 vdd.n1376 vss 0.012467f
C1587 vdd.n1377 vss 0.012641f
C1588 vdd.n1378 vss 0.005299f
C1589 vdd.n1379 vss 0.005299f
C1590 vdd.n1380 vss 0.013679f
C1591 vdd.n1381 vss 0.012467f
C1592 vdd.n1382 vss 0.027705f
C1593 vdd.n1383 vss 0.021645f
C1594 vdd.n1384 vss 0.012467f
C1595 vdd.n1385 vss 0.013853f
C1596 vdd.n1386 vss 0.005299f
C1597 vdd.n1387 vss 0.005299f
C1598 vdd.n1388 vss 0.013853f
C1599 vdd.n1389 vss 0.012467f
C1600 vdd.n1390 vss 0.027705f
C1601 vdd.n1391 vss 0.020952f
C1602 vdd.n1392 vss 0.012467f
C1603 vdd.n1393 vss 0.013853f
C1604 vdd.n1394 vss 0.005299f
C1605 vdd.n1395 vss 0.005299f
C1606 vdd.n1396 vss 0.013853f
C1607 vdd.n1397 vss 0.012467f
C1608 vdd.n1398 vss 0.027705f
C1609 vdd.n1399 vss 0.02026f
C1610 vdd.n1400 vss 0.012467f
C1611 vdd.n1401 vss 0.013853f
C1612 vdd.n1402 vss 0.005299f
C1613 vdd.n1403 vss 0.005299f
C1614 vdd.n1404 vss 0.005299f
C1615 vdd.n1405 vss 0.013679f
C1616 vdd.n1406 vss 0.012467f
C1617 vdd.n1407 vss 0.027705f
C1618 vdd.n1408 vss 0.019567f
C1619 vdd.n1409 vss 0.012467f
C1620 vdd.n1410 vss 0.013853f
C1621 vdd.n1411 vss 0.005299f
C1622 vdd.n1412 vss 0.005299f
C1623 vdd.n1413 vss 0.013853f
C1624 vdd.n1414 vss 0.012467f
C1625 vdd.n1415 vss 0.027705f
C1626 vdd.n1416 vss 0.018874f
C1627 vdd.n1417 vss 0.012467f
C1628 vdd.n1418 vss 0.013853f
C1629 vdd.n1419 vss 0.005299f
C1630 vdd.n1420 vss 0.005299f
C1631 vdd.n1421 vss 0.013853f
C1632 vdd.n1422 vss 0.012467f
C1633 vdd.n1423 vss 0.027705f
C1634 vdd.n1424 vss 0.018182f
C1635 vdd.n1425 vss 0.012467f
C1636 vdd.n1426 vss 0.013853f
C1637 vdd.n1427 vss 0.005299f
C1638 vdd.n1428 vss 0.00276f
C1639 vdd.n1429 vss 0.012641f
C1640 vdd.n1430 vss 0.013679f
C1641 vdd.n1431 vss 0.005188f
C1642 vdd.n1432 vss 0.005299f
C1643 vdd.n1433 vss 0.013853f
C1644 vdd.n1434 vss 0.012467f
C1645 vdd.n1435 vss 0.017489f
C1646 vdd.n1436 vss 0.214207f
C1647 vdd.n1437 vss 0.024069f
C1648 vdd.n1438 vss 0.012467f
C1649 vdd.n1439 vss 0.013853f
C1650 vdd.n1440 vss 0.005299f
C1651 vdd.n1441 vss 0.005299f
C1652 vdd.n1442 vss 0.013853f
C1653 vdd.n1443 vss 0.012467f
C1654 vdd.n1444 vss 0.016796f
C1655 vdd.n1445 vss 0.214207f
C1656 vdd.n1446 vss 0.024762f
C1657 vdd.n1447 vss 0.012467f
C1658 vdd.n1448 vss 0.013853f
C1659 vdd.n1449 vss 0.005299f
C1660 vdd.n1450 vss 0.005299f
C1661 vdd.n1451 vss 0.013853f
C1662 vdd.n1452 vss 0.012467f
C1663 vdd.n1453 vss 0.016104f
C1664 vdd.n1454 vss 0.214207f
C1665 vdd.n1455 vss 0.025454f
C1666 vdd.n1456 vss 0.012467f
C1667 vdd.n1457 vss 0.012641f
C1668 vdd.n1458 vss 0.013679f
C1669 vdd.n1459 vss 0.005299f
C1670 vdd.n1460 vss 0.005299f
C1671 vdd.n1461 vss 0.013853f
C1672 vdd.n1462 vss 0.012467f
C1673 vdd.n1463 vss 0.015411f
C1674 vdd.n1464 vss 0.214207f
C1675 vdd.n1465 vss 0.026147f
C1676 vdd.n1466 vss 0.012467f
C1677 vdd.n1467 vss 0.013853f
C1678 vdd.n1468 vss 0.005299f
C1679 vdd.n1469 vss 0.005299f
C1680 vdd.n1470 vss 0.013853f
C1681 vdd.n1471 vss 0.012467f
C1682 vdd.n1472 vss 0.014718f
C1683 vdd.n1473 vss 0.214207f
C1684 vdd.n1474 vss 0.02684f
C1685 vdd.n1475 vss 0.012467f
C1686 vdd.n1476 vss 0.013853f
C1687 vdd.n1477 vss 0.005299f
C1688 vdd.n1478 vss 0.005299f
C1689 vdd.n1479 vss 0.013853f
C1690 vdd.n1480 vss 0.012467f
C1691 vdd.n1481 vss 0.014026f
C1692 vdd.n1482 vss 0.214207f
C1693 vdd.n1483 vss 0.027532f
C1694 vdd.n1484 vss 0.012467f
C1695 vdd.n1485 vss 0.012641f
C1696 vdd.n1486 vss 0.013679f
C1697 vdd.n1487 vss 0.005299f
C1698 vdd.n1488 vss 0.002944f
C1699 vdd.n1489 vss 0.013853f
C1700 vdd.n1490 vss 0.013927f
C1701 vdd.n1491 vss 0.027705f
C1702 vdd.n1492 vss 0.027705f
C1703 vdd.n1493 vss 0.013853f
C1704 vdd.n1494 vss 0.027705f
C1705 vdd.n1495 vss 0.027705f
C1706 vdd.n1496 vss 0.027705f
C1707 vdd.n1497 vss 0.027705f
C1708 vdd.n1498 vss 0.027705f
C1709 vdd.n1499 vss 0.027705f
C1710 vdd.n1500 vss 0.108689f
C1711 vdd.n1501 vss 0.013853f
C1712 vdd.n1502 vss 0.027705f
C1713 vdd.n1503 vss 0.027705f
C1714 vdd.n1504 vss 0.012899f
C1715 vdd.n1505 vss 0.013853f
C1716 vdd.n1506 vss 0.004715f
C1717 vdd.n1507 vss 0.034552f
C1718 vdd.n1508 vss 0.063804f
C1719 vdd.n1509 vss 0.182361f
C1720 vdd.n1510 vss 2.60984f
C1721 vdd.t50 vss 0.679306f
C1722 vdd.t6 vss 0.550915f
C1723 vdd.t92 vss 0.550915f
C1724 vdd.t106 vss 0.550915f
C1725 vdd.t225 vss 0.550915f
C1726 vdd.t84 vss 0.550915f
C1727 vdd.t177 vss 0.452871f
C1728 vdd.n1511 vss 0.054019f
C1729 vdd.n1512 vss 0.44733f
C1730 vdd.n1513 vss 0.002649f
C1731 vdd.n1514 vss 0.003827f
C1732 vdd.n1515 vss 0.005299f
C1733 vdd.n1516 vss 0.005299f
C1734 vdd.n1517 vss 0.005299f
C1735 vdd.n1518 vss 0.005299f
C1736 vdd.n1519 vss 0.029062f
C1737 vdd.n1520 vss 0.004035f
C1738 vdd.n1521 vss 0.005299f
C1739 vdd.n1522 vss 0.005299f
C1740 vdd.n1523 vss 0.007669f
C1741 vdd.n1524 vss 0.02866f
C1742 vdd.t140 vss 0.018831f
C1743 vdd.t25 vss 0.018831f
C1744 vdd.n1525 vss 0.042405f
C1745 vdd.n1526 vss 0.238626f
C1746 vdd.n1527 vss 0.046465f
C1747 vdd.n1528 vss 0.048562f
C1748 vdd.n1529 vss 0.048863f
C1749 vdd.n1530 vss 0.048863f
C1750 vdd.n1531 vss 0.048863f
C1751 vdd.n1532 vss 0.044067f
C1752 vdd.n1533 vss 0.02866f
C1753 vdd.n1534 vss 0.02543f
C1754 vdd.n1535 vss 0.005299f
C1755 vdd.n1536 vss 0.005299f
C1756 vdd.n1537 vss 0.005299f
C1757 vdd.n1538 vss 0.005299f
C1758 vdd.n1539 vss 0.021796f
C1759 vdd.n1540 vss 0.02866f
C1760 vdd.n1541 vss 0.028777f
C1761 vdd.n1542 vss 0.048562f
C1762 vdd.n1543 vss 0.048562f
C1763 vdd.n1544 vss 0.030876f
C1764 vdd.n1545 vss 0.048562f
C1765 vdd.n1546 vss 0.048562f
C1766 vdd.n1547 vss 0.041967f
C1767 vdd.n1548 vss 0.02866f
C1768 vdd.n1549 vss 0.014935f
C1769 vdd.n1550 vss 0.004121f
C1770 vdd.n1551 vss 0.005299f
C1771 vdd.n1552 vss 0.018567f
C1772 vdd.n1553 vss 0.005299f
C1773 vdd.n1554 vss 0.005299f
C1774 vdd.n1555 vss 0.005299f
C1775 vdd.n1556 vss 0.005299f
C1776 vdd.n1557 vss 0.022201f
C1777 vdd.n1558 vss 0.02866f
C1778 vdd.n1559 vss 0.007264f
C1779 vdd.n1560 vss 0.005299f
C1780 vdd.n1561 vss 0.004636f
C1781 vdd.n1562 vss 0.005299f
C1782 vdd.n1563 vss 0.005299f
C1783 vdd.n1564 vss 0.005299f
C1784 vdd.n1565 vss 0.005299f
C1785 vdd.n1566 vss 0.005299f
C1786 vdd.n1567 vss 0.005299f
C1787 vdd.n1568 vss 0.005299f
C1788 vdd.n1569 vss 0.005299f
C1789 vdd.n1570 vss 0.003227f
C1790 vdd.n1571 vss 0.02866f
C1791 vdd.n1572 vss 0.03987f
C1792 vdd.n1573 vss 0.048863f
C1793 vdd.n1574 vss 0.048562f
C1794 vdd.n1575 vss 0.033275f
C1795 vdd.n1576 vss 0.02866f
C1796 vdd.n1577 vss 8.05e-19
C1797 vdd.n1578 vss 0.005299f
C1798 vdd.n1579 vss 0.005299f
C1799 vdd.n1580 vss 0.004439f
C1800 vdd.n1581 vss 0.005299f
C1801 vdd.n1582 vss 0.005299f
C1802 vdd.n1583 vss 0.008071f
C1803 vdd.n1584 vss 0.02866f
C1804 vdd.n1585 vss 0.037471f
C1805 vdd.n1586 vss 0.048562f
C1806 vdd.n1587 vss 0.048562f
C1807 vdd.n1588 vss 0.035372f
C1808 vdd.n1589 vss 0.02866f
C1809 vdd.n1590 vss 0.011706f
C1810 vdd.n1591 vss 0.005299f
C1811 vdd.n1592 vss 0.005299f
C1812 vdd.n1593 vss 0.015337f
C1813 vdd.n1594 vss 0.005299f
C1814 vdd.n1595 vss 0.005299f
C1815 vdd.n1596 vss 0.018972f
C1816 vdd.n1597 vss 0.02866f
C1817 vdd.n1598 vss 0.035372f
C1818 vdd.n1599 vss 0.048863f
C1819 vdd.n1600 vss 0.048562f
C1820 vdd.n1601 vss 0.048562f
C1821 vdd.n1605 vss 0.048562f
C1822 vdd.n1606 vss 0.048562f
C1823 vdd.n1607 vss 0.048562f
C1824 vdd.n1608 vss 0.048562f
C1825 vdd.n1609 vss 0.048562f
C1826 vdd.n1610 vss 0.048863f
C1827 vdd.n1611 vss 0.048863f
C1828 vdd.n1612 vss 0.048863f
C1829 vdd.n1613 vss 0.048863f
C1830 vdd.n1614 vss 0.048562f
C1831 vdd.n1615 vss 0.048562f
C1832 vdd.n1616 vss 0.048562f
C1833 vdd.n1617 vss 0.048562f
C1834 vdd.n1618 vss 0.048562f
C1835 vdd.n1620 vss 0.08264f
C1836 vdd.n1621 vss 0.005299f
C1837 vdd.n1622 vss 0.005299f
C1838 vdd.n1623 vss 0.005299f
C1839 vdd.n1624 vss 0.005299f
C1840 vdd.n1625 vss 0.005299f
C1841 vdd.n1626 vss 0.005299f
C1842 vdd.n1627 vss 0.005299f
C1843 vdd.n1628 vss 0.005299f
C1844 vdd.n1629 vss 0.005299f
C1845 vdd.n1630 vss 0.005299f
C1846 vdd.n1631 vss 0.005299f
C1847 vdd.n1632 vss 0.00298f
C1848 vdd.n1633 vss 0.020182f
C1849 vdd.n1634 vss 0.060712f
C1850 vdd.n1635 vss 0.00673f
C1851 vdd.n1636 vss 0.02866f
C1852 vdd.n1637 vss 0.012513f
C1853 vdd.n1638 vss 0.00673f
C1854 vdd.n1639 vss 0.060712f
C1855 vdd.n1640 vss 0.089826f
C1856 vdd.n1641 vss 0.086233f
C1857 vdd.n1642 vss 0.048562f
C1858 vdd.n1643 vss 0.048562f
C1859 vdd.n1644 vss 0.048562f
C1860 vdd.n1645 vss 0.048863f
C1861 vdd.n1646 vss 0.03777f
C1862 vdd.n1647 vss 0.02866f
C1863 vdd.n1648 vss 0.023008f
C1864 vdd.n1649 vss 0.005299f
C1865 vdd.n1650 vss 0.005299f
C1866 vdd.n1651 vss 0.02664f
C1867 vdd.n1652 vss 0.005299f
C1868 vdd.n1653 vss 0.060712f
C1869 vdd.n1654 vss 0.006739f
C1870 vdd.n1655 vss 0.023008f
C1871 vdd.n1656 vss 0.002825f
C1872 vdd.n1657 vss 0.004752f
C1873 vdd.n1658 vss 0.060302f
C1874 vdd.n1659 vss 2.11895f
C1875 vdd.n1660 vss 0.095215f
C1876 vdd.n1661 vss 0.048562f
C1877 vdd.n1662 vss 0.048562f
C1878 vdd.n1663 vss 0.048863f
C1879 vdd.t265 vss 0.018831f
C1880 vdd.t63 vss 0.018831f
C1881 vdd.n1664 vss 0.042405f
C1882 vdd.n1665 vss 0.238626f
C1883 vdd.n1666 vss 0.03987f
C1884 vdd.n1667 vss 0.048562f
C1885 vdd.n1668 vss 0.048562f
C1886 vdd.n1669 vss 0.048863f
C1887 vdd.n1670 vss 0.048863f
C1888 vdd.n1671 vss 0.02866f
C1889 vdd.n1672 vss 0.01655f
C1890 vdd.n1673 vss 0.005299f
C1891 vdd.n1674 vss 0.005299f
C1892 vdd.n1675 vss 0.020182f
C1893 vdd.n1676 vss 0.005299f
C1894 vdd.n1677 vss 0.005299f
C1895 vdd.n1678 vss 0.023816f
C1896 vdd.n1679 vss 0.005299f
C1897 vdd.n1680 vss 0.005299f
C1898 vdd.n1681 vss 0.02866f
C1899 vdd.n1682 vss 0.027448f
C1900 vdd.n1683 vss 0.005299f
C1901 vdd.n1684 vss 0.005299f
C1902 vdd.n1685 vss 0.029062f
C1903 vdd.n1686 vss 0.005299f
C1904 vdd.n1687 vss 0.005299f
C1905 vdd.n1688 vss 0.002017f
C1906 vdd.n1689 vss 0.02866f
C1907 vdd.n1690 vss 0.030876f
C1908 vdd.n1691 vss 0.048562f
C1909 vdd.n1692 vss 0.048562f
C1910 vdd.n1693 vss 0.041967f
C1911 vdd.n1694 vss 0.02866f
C1912 vdd.n1695 vss 0.005649f
C1913 vdd.n1696 vss 0.005299f
C1914 vdd.n1697 vss 0.005299f
C1915 vdd.n1698 vss 0.009283f
C1916 vdd.n1699 vss 0.005299f
C1917 vdd.n1700 vss 0.005299f
C1918 vdd.n1701 vss 0.01332f
C1919 vdd.n1702 vss 0.02866f
C1920 vdd.n1703 vss 0.028779f
C1921 vdd.n1704 vss 0.048863f
C1922 vdd.n1705 vss 0.048562f
C1923 vdd.n1706 vss 0.044365f
C1924 vdd.n1707 vss 0.02866f
C1925 vdd.n1708 vss 0.016952f
C1926 vdd.n1709 vss 0.005299f
C1927 vdd.n1710 vss 0.005299f
C1928 vdd.n1711 vss 0.005299f
C1929 vdd.n1712 vss 0.005299f
C1930 vdd.n1713 vss 0.020586f
C1931 vdd.n1714 vss 0.005299f
C1932 vdd.n1715 vss 0.005299f
C1933 vdd.n1716 vss 0.005299f
C1934 vdd.n1717 vss 0.005299f
C1935 vdd.n1718 vss 0.029062f
C1936 vdd.n1719 vss 0.001613f
C1937 vdd.n1720 vss 0.005299f
C1938 vdd.n1721 vss 0.005299f
C1939 vdd.n1722 vss 0.005247f
C1940 vdd.n1723 vss 0.02866f
C1941 vdd.t129 vss 0.018831f
C1942 vdd.t17 vss 0.018831f
C1943 vdd.n1724 vss 0.042405f
C1944 vdd.n1725 vss 0.238626f
C1945 vdd.n1726 vss 0.026378f
C1946 vdd.n1727 vss 0.048562f
C1947 vdd.n1728 vss 0.048562f
C1948 vdd.n1729 vss 0.048562f
C1949 vdd.t267 vss 0.018831f
C1950 vdd.t166 vss 0.018831f
C1951 vdd.n1730 vss 0.042405f
C1952 vdd.n1731 vss 0.048562f
C1953 vdd.n1732 vss 0.048562f
C1954 vdd.t290 vss 0.018831f
C1955 vdd.t297 vss 0.018831f
C1956 vdd.n1733 vss 0.042405f
C1957 vdd.n1734 vss 0.041969f
C1958 vdd.n1735 vss 0.048562f
C1959 vdd.t210 vss 0.018831f
C1960 vdd.t314 vss 0.018831f
C1961 vdd.n1736 vss 0.042405f
C1962 vdd.n1737 vss 0.238626f
C1963 vdd.t234 vss 0.018831f
C1964 vdd.t27 vss 0.018831f
C1965 vdd.n1738 vss 0.042405f
C1966 vdd.n1739 vss 0.238626f
C1967 vdd.n1740 vss 0.048562f
C1968 vdd.t258 vss 0.018831f
C1969 vdd.t145 vss 0.018831f
C1970 vdd.n1741 vss 0.042405f
C1971 vdd.n1742 vss 0.238927f
C1972 vdd.n1743 vss 0.048562f
C1973 vdd.t273 vss 0.018831f
C1974 vdd.t171 vss 0.018831f
C1975 vdd.n1744 vss 0.042405f
C1976 vdd.n1745 vss 0.238626f
C1977 vdd.n1746 vss 0.048562f
C1978 vdd.t174 vss 0.018831f
C1979 vdd.t301 vss 0.018831f
C1980 vdd.n1747 vss 0.042405f
C1981 vdd.n1748 vss 0.238626f
C1982 vdd.n1749 vss 0.048863f
C1983 vdd.n1750 vss 0.048562f
C1984 vdd.n1751 vss 0.030575f
C1985 vdd.n1752 vss 0.048863f
C1986 vdd.n1753 vss 0.040171f
C1987 vdd.n1754 vss 0.048863f
C1988 vdd.n1755 vss 0.048562f
C1989 vdd.n1756 vss 0.032974f
C1990 vdd.n1757 vss 0.048562f
C1991 vdd.n1758 vss 0.03777f
C1992 vdd.n1759 vss 0.048562f
C1993 vdd.n1760 vss 0.048562f
C1994 vdd.n1761 vss 0.035073f
C1995 vdd.n1762 vss 0.048562f
C1996 vdd.n1763 vss 0.035673f
C1997 vdd.n1764 vss 0.048863f
C1998 vdd.n1765 vss 0.048863f
C1999 vdd.n1766 vss 0.037471f
C2000 vdd.n1767 vss 0.048562f
C2001 vdd.n1768 vss 0.033275f
C2002 vdd.n1769 vss 0.048562f
C2003 vdd.n1770 vss 0.048562f
C2004 vdd.n1771 vss 0.039569f
C2005 vdd.n1772 vss 0.048562f
C2006 vdd.n1773 vss 0.031175f
C2007 vdd.n1774 vss 0.048562f
C2008 vdd.n1775 vss 0.048863f
C2009 vdd.n1776 vss 0.048863f
C2010 vdd.n1777 vss 0.048863f
C2011 vdd.n1778 vss 0.028777f
C2012 vdd.n1779 vss 0.238626f
C2013 vdd.n1780 vss 0.044067f
C2014 vdd.n1781 vss 0.048562f
C2015 vdd.n1782 vss 0.048562f
C2016 vdd.n1783 vss 0.048562f
C2017 vdd.n1784 vss 0.026679f
C2018 vdd.n1785 vss 0.238626f
C2019 vdd.n1786 vss 0.046164f
C2020 vdd.n1787 vss 0.048863f
C2021 vdd.n1788 vss 0.048863f
C2022 vdd.n1789 vss 0.048863f
C2023 vdd.n1790 vss 0.048562f
C2024 vdd.n1791 vss 0.048562f
C2025 vdd.n1792 vss 0.034714f
C2026 vdd.n1793 vss 0.00242f
C2027 vdd.n1794 vss 0.008647f
C2028 vdd.n1795 vss 0.008647f
C2029 vdd.n1796 vss 0.03257f
C2030 vdd.n1797 vss 0.008647f
C2031 vdd.n1798 vss 0.005299f
C2032 vdd.n1799 vss 0.032171f
C2033 vdd.n1800 vss 0.005299f
C2034 vdd.n1801 vss 0.005299f
C2035 vdd.n1802 vss 0.032171f
C2036 vdd.n1803 vss 0.005299f
C2037 vdd.n1804 vss 0.005299f
C2038 vdd.n1805 vss 0.032171f
C2039 vdd.n1806 vss 0.005299f
C2040 vdd.n1807 vss 0.005299f
C2041 vdd.n1808 vss 0.032171f
C2042 vdd.n1809 vss 0.004416f
C2043 vdd.n1810 vss 0.002649f
C2044 vdd.n1811 vss 0.003532f
C2045 vdd.n1812 vss 0.032171f
C2046 vdd.n1813 vss 0.005299f
C2047 vdd.n1814 vss 0.005299f
C2048 vdd.n1815 vss 0.032171f
C2049 vdd.n1816 vss 0.005299f
C2050 vdd.n1817 vss 0.005299f
C2051 vdd.n1818 vss 0.032567f
C2052 vdd.n1819 vss 0.005299f
C2053 vdd.n1820 vss 0.005299f
C2054 vdd.n1821 vss 0.005299f
C2055 vdd.n1822 vss 0.03098f
C2056 vdd.n1823 vss 0.005299f
C2057 vdd.n1824 vss 0.005299f
C2058 vdd.n1825 vss 0.032171f
C2059 vdd.n1826 vss 0.005299f
C2060 vdd.n1827 vss 0.005299f
C2061 vdd.n1828 vss 0.032171f
C2062 vdd.n1829 vss 0.005299f
C2063 vdd.n1830 vss 0.005299f
C2064 vdd.n1831 vss 0.032171f
C2065 vdd.n1832 vss 0.005299f
C2066 vdd.n1833 vss 0.005299f
C2067 vdd.n1834 vss 0.032171f
C2068 vdd.n1835 vss 0.005299f
C2069 vdd.n1836 vss 0.005299f
C2070 vdd.n1837 vss 0.032171f
C2071 vdd.n1838 vss 0.005299f
C2072 vdd.n1839 vss 0.005299f
C2073 vdd.n1840 vss 0.032567f
C2074 vdd.n1841 vss 0.005299f
C2075 vdd.n1842 vss 0.005299f
C2076 vdd.n1843 vss 0.032171f
C2077 vdd.n1844 vss 0.005299f
C2078 vdd.n1845 vss 0.005299f
C2079 vdd.n1846 vss 0.005299f
C2080 vdd.n1847 vss 0.031376f
C2081 vdd.n1848 vss 0.005299f
C2082 vdd.n1849 vss 0.005299f
C2083 vdd.n1850 vss 0.032171f
C2084 vdd.n1851 vss 0.005299f
C2085 vdd.n1852 vss 0.005299f
C2086 vdd.n1853 vss 0.032171f
C2087 vdd.n1854 vss 0.005299f
C2088 vdd.n1855 vss 0.005299f
C2089 vdd.n1856 vss 0.032171f
C2090 vdd.n1857 vss 0.005299f
C2091 vdd.n1858 vss 0.005299f
C2092 vdd.n1859 vss 0.032171f
C2093 vdd.n1860 vss 0.005299f
C2094 vdd.n1861 vss 0.005299f
C2095 vdd.n1862 vss 0.032567f
C2096 vdd.n1863 vss 0.005299f
C2097 vdd.n1864 vss 0.005299f
C2098 vdd.n1865 vss 0.032171f
C2099 vdd.n1866 vss 0.005299f
C2100 vdd.n1867 vss 0.005299f
C2101 vdd.n1868 vss 0.032171f
C2102 vdd.n1869 vss 0.028595f
C2103 vdd.n1870 vss 0.042268f
C2104 vdd.n1871 vss 0.048562f
C2105 vdd.n1872 vss 0.048562f
C2106 vdd.n1873 vss 0.048562f
C2107 vdd.n1874 vss 0.048562f
C2108 vdd.n1875 vss 0.048562f
C2109 vdd.n1877 vss 0.048562f
C2110 vdd.n1878 vss 0.048562f
C2111 vdd.n1879 vss 0.048562f
C2112 vdd.n1880 vss 0.048562f
C2113 vdd.n1881 vss 0.048562f
C2114 vdd.n1882 vss 0.048562f
C2115 vdd.n1883 vss 0.048562f
C2116 vdd.n1884 vss 0.048562f
C2117 vdd.n1886 vss 0.075454f
C2118 vdd.n1888 vss 0.048863f
C2119 vdd.n1889 vss 0.048863f
C2120 vdd.n1890 vss 0.048863f
C2121 vdd.n1891 vss 0.048863f
C2122 vdd.n1892 vss 0.048562f
C2123 vdd.n1893 vss 0.048562f
C2124 vdd.n1895 vss 0.095215f
C2125 vdd.n1896 vss 0.053895f
C2126 vdd.n1897 vss 0.060712f
C2127 vdd.n1898 vss 0.006739f
C2128 vdd.n1899 vss 0.031774f
C2129 vdd.n1900 vss 0.006739f
C2130 vdd.n1901 vss 0.060712f
C2131 vdd.n1902 vss 0.00673f
C2132 vdd.n1903 vss 0.032171f
C2133 vdd.n1904 vss 0.019857f
C2134 vdd.n1905 vss 0.048863f
C2135 vdd.n1906 vss 0.048863f
C2136 vdd.n1907 vss 0.048562f
C2137 vdd.n1908 vss 0.048562f
C2138 vdd.n1909 vss 0.048562f
C2139 vdd.n1910 vss 0.028478f
C2140 vdd.n1911 vss 0.238626f
C2141 vdd.n1912 vss 0.044365f
C2142 vdd.n1913 vss 0.048562f
C2143 vdd.n1914 vss 0.048562f
C2144 vdd.n1915 vss 0.048562f
C2145 vdd.n1916 vss 0.028595f
C2146 vdd.n1917 vss 0.028597f
C2147 vdd.t211 vss 0.018831f
C2148 vdd.t1 vss 0.018831f
C2149 vdd.n1918 vss 0.042405f
C2150 vdd.n1919 vss 0.028595f
C2151 vdd.n1920 vss 0.048562f
C2152 vdd.n1921 vss 0.048562f
C2153 vdd.n1922 vss 0.028595f
C2154 vdd.t143 vss 0.018831f
C2155 vdd.t31 vss 0.018831f
C2156 vdd.n1923 vss 0.042405f
C2157 vdd.n1924 vss 0.028597f
C2158 vdd.n1925 vss 0.028595f
C2159 vdd.n1926 vss 0.044067f
C2160 vdd.n1927 vss 0.048562f
C2161 vdd.t260 vss 0.018831f
C2162 vdd.t151 vss 0.018831f
C2163 vdd.n1928 vss 0.042405f
C2164 vdd.n1929 vss 0.238626f
C2165 vdd.n1930 vss 0.028597f
C2166 vdd.n1931 vss 0.028595f
C2167 vdd.n1932 vss 0.028597f
C2168 vdd.t275 vss 0.018831f
C2169 vdd.t91 vss 0.018831f
C2170 vdd.n1933 vss 0.042405f
C2171 vdd.n1934 vss 0.238626f
C2172 vdd.n1935 vss 0.048562f
C2173 vdd.n1936 vss 0.028595f
C2174 vdd.n1937 vss 0.028597f
C2175 vdd.n1938 vss 0.028595f
C2176 vdd.t97 vss 0.018831f
C2177 vdd.t304 vss 0.018831f
C2178 vdd.n1939 vss 0.042405f
C2179 vdd.n1940 vss 0.238925f
C2180 vdd.n1941 vss 0.048562f
C2181 vdd.n1942 vss 0.028595f
C2182 vdd.n1943 vss 0.028597f
C2183 vdd.n1944 vss 0.028595f
C2184 vdd.t220 vss 0.018831f
C2185 vdd.t101 vss 0.018831f
C2186 vdd.n1945 vss 0.042405f
C2187 vdd.n1946 vss 0.238626f
C2188 vdd.n1947 vss 0.048562f
C2189 vdd.n1948 vss 0.028597f
C2190 vdd.n1949 vss 0.028595f
C2191 vdd.n1950 vss 0.028597f
C2192 vdd.t152 vss 0.018831f
C2193 vdd.t39 vss 0.018831f
C2194 vdd.n1951 vss 0.042405f
C2195 vdd.n1952 vss 0.238626f
C2196 vdd.n1953 vss 0.048863f
C2197 vdd.n1954 vss 0.028595f
C2198 vdd.n1955 vss 0.028595f
C2199 vdd.n1956 vss 0.028597f
C2200 vdd.t263 vss 0.018831f
C2201 vdd.t157 vss 0.018831f
C2202 vdd.n1957 vss 0.042405f
C2203 vdd.n1958 vss 0.238626f
C2204 vdd.n1959 vss 0.048562f
C2205 vdd.n1960 vss 0.028595f
C2206 vdd.n1961 vss 0.028597f
C2207 vdd.n1962 vss 0.028595f
C2208 vdd.t45 vss 0.018831f
C2209 vdd.t276 vss 0.018831f
C2210 vdd.n1963 vss 0.042405f
C2211 vdd.n1964 vss 0.238626f
C2212 vdd.n1965 vss 0.048863f
C2213 vdd.n1966 vss 0.028597f
C2214 vdd.n1967 vss 0.028595f
C2215 vdd.n1968 vss 0.028595f
C2216 vdd.t109 vss 0.018831f
C2217 vdd.t308 vss 0.018831f
C2218 vdd.n1969 vss 0.042405f
C2219 vdd.n1970 vss 0.238626f
C2220 vdd.n1971 vss 0.048562f
C2221 vdd.n1972 vss 0.028597f
C2222 vdd.n1973 vss 0.028595f
C2223 vdd.n1974 vss 0.028597f
C2224 vdd.t227 vss 0.073257f
C2225 vdd.n1975 vss 0.245436f
C2226 vdd.n1976 vss 0.048562f
C2227 vdd.n1977 vss 0.006445f
C2228 vdd.n1978 vss 0.006445f
C2229 vdd.n1979 vss 0.005299f
C2230 vdd.n1980 vss 0.005299f
C2231 vdd.n1981 vss 0.005299f
C2232 vdd.n1982 vss 0.005299f
C2233 vdd.n1983 vss 0.029788f
C2234 vdd.n1984 vss 0.005299f
C2235 vdd.n1985 vss 0.005299f
C2236 vdd.n1986 vss 0.005299f
C2237 vdd.n1987 vss 0.005299f
C2238 vdd.n1988 vss 0.005299f
C2239 vdd.n1989 vss 0.005299f
C2240 vdd.n1990 vss 0.005299f
C2241 vdd.n1991 vss 0.005299f
C2242 vdd.n1992 vss 0.005299f
C2243 vdd.n1993 vss 0.005299f
C2244 vdd.n1994 vss 0.005299f
C2245 vdd.n1995 vss 0.005299f
C2246 vdd.n1996 vss 0.005299f
C2247 vdd.n1997 vss 0.005299f
C2248 vdd.n1998 vss 0.005299f
C2249 vdd.n1999 vss 0.005299f
C2250 vdd.n2000 vss 0.005299f
C2251 vdd.n2001 vss 0.005299f
C2252 vdd.n2002 vss 0.005299f
C2253 vdd.n2003 vss 0.030582f
C2254 vdd.n2004 vss 0.005299f
C2255 vdd.n2005 vss 0.005299f
C2256 vdd.n2006 vss 0.005299f
C2257 vdd.n2007 vss 0.005299f
C2258 vdd.n2008 vss 0.005299f
C2259 vdd.n2009 vss 0.005299f
C2260 vdd.n2010 vss 0.005299f
C2261 vdd.n2011 vss 0.005299f
C2262 vdd.n2012 vss 0.005299f
C2263 vdd.n2013 vss 0.005299f
C2264 vdd.n2014 vss 0.005299f
C2265 vdd.n2015 vss 0.005299f
C2266 vdd.n2016 vss 0.005299f
C2267 vdd.n2017 vss 0.005299f
C2268 vdd.n2018 vss 0.005299f
C2269 vdd.n2019 vss 0.002833f
C2270 vdd.n2020 vss 0.005299f
C2271 vdd.n2021 vss 0.005299f
C2272 vdd.n2022 vss 0.03098f
C2273 vdd.n2023 vss 0.005299f
C2274 vdd.n2024 vss 0.005299f
C2275 vdd.n2025 vss 0.005299f
C2276 vdd.n2026 vss 0.005299f
C2277 vdd.n2027 vss 0.002649f
C2278 vdd.n2028 vss 0.005115f
C2279 vdd.n2029 vss 0.005299f
C2280 vdd.n2030 vss 0.005299f
C2281 vdd.n2031 vss 0.005299f
C2282 vdd.n2032 vss 0.005299f
C2283 vdd.n2033 vss 0.005299f
C2284 vdd.n2034 vss 0.005299f
C2285 vdd.n2035 vss 0.005299f
C2286 vdd.n2036 vss 0.005299f
C2287 vdd.n2037 vss 0.028595f
C2288 vdd.n2038 vss 0.005299f
C2289 vdd.n2039 vss 0.005299f
C2290 vdd.n2040 vss 0.005299f
C2291 vdd.n2041 vss 0.005299f
C2292 vdd.n2042 vss 0.005299f
C2293 vdd.n2043 vss 0.005299f
C2294 vdd.n2044 vss 0.031376f
C2295 vdd.n2045 vss 0.005299f
C2296 vdd.n2046 vss 0.005299f
C2297 vdd.n2047 vss 0.028597f
C2298 vdd.n2048 vss 0.005299f
C2299 vdd.n2049 vss 0.005299f
C2300 vdd.n2050 vss 0.005299f
C2301 vdd.n2051 vss 0.005299f
C2302 vdd.n2052 vss 0.005299f
C2303 vdd.n2053 vss 0.005299f
C2304 vdd.n2054 vss 0.005299f
C2305 vdd.n2055 vss 0.005299f
C2306 vdd.n2056 vss 0.005299f
C2307 vdd.n2057 vss 0.005299f
C2308 vdd.n2058 vss 0.005299f
C2309 vdd.n2059 vss 0.005299f
C2310 vdd.n2060 vss 0.005299f
C2311 vdd.n2061 vss 0.032171f
C2312 vdd.n2062 vss 0.005299f
C2313 vdd.n2063 vss 0.005299f
C2314 vdd.n2064 vss 0.032171f
C2315 vdd.n2065 vss 0.005299f
C2316 vdd.n2066 vss 0.005299f
C2317 vdd.n2067 vss 0.032171f
C2318 vdd.n2068 vss 0.005299f
C2319 vdd.n2069 vss 0.005299f
C2320 vdd.n2070 vss 0.032171f
C2321 vdd.n2071 vss 0.005299f
C2322 vdd.n2072 vss 0.005299f
C2323 vdd.n2073 vss 0.005299f
C2324 vdd.n2074 vss 0.029391f
C2325 vdd.n2075 vss 0.005299f
C2326 vdd.n2076 vss 0.005299f
C2327 vdd.n2077 vss 0.032171f
C2328 vdd.n2078 vss 0.005299f
C2329 vdd.n2079 vss 0.005299f
C2330 vdd.n2080 vss 0.032567f
C2331 vdd.n2081 vss 0.005299f
C2332 vdd.n2082 vss 0.005299f
C2333 vdd.n2083 vss 0.032171f
C2334 vdd.n2084 vss 0.005299f
C2335 vdd.n2085 vss 0.005299f
C2336 vdd.n2086 vss 0.032171f
C2337 vdd.n2087 vss 0.005299f
C2338 vdd.n2088 vss 0.005299f
C2339 vdd.n2089 vss 0.032171f
C2340 vdd.n2090 vss 0.005299f
C2341 vdd.n2091 vss 0.005299f
C2342 vdd.n2092 vss 0.032171f
C2343 vdd.n2093 vss 0.005299f
C2344 vdd.n2094 vss 0.005299f
C2345 vdd.n2095 vss 0.032171f
C2346 vdd.n2096 vss 0.005299f
C2347 vdd.n2097 vss 0.005299f
C2348 vdd.n2098 vss 0.005299f
C2349 vdd.n2099 vss 0.029788f
C2350 vdd.n2100 vss 0.005299f
C2351 vdd.n2101 vss 0.005299f
C2352 vdd.n2102 vss 0.032567f
C2353 vdd.n2103 vss 0.005299f
C2354 vdd.n2104 vss 0.005299f
C2355 vdd.n2105 vss 0.032171f
C2356 vdd.n2106 vss 0.005299f
C2357 vdd.n2107 vss 0.005299f
C2358 vdd.n2108 vss 0.032171f
C2359 vdd.n2109 vss 0.005299f
C2360 vdd.n2110 vss 0.005299f
C2361 vdd.n2111 vss 0.032171f
C2362 vdd.n2112 vss 0.005299f
C2363 vdd.n2113 vss 0.005299f
C2364 vdd.n2114 vss 0.032171f
C2365 vdd.n2115 vss 0.005299f
C2366 vdd.n2116 vss 0.005299f
C2367 vdd.n2117 vss 0.032171f
C2368 vdd.n2118 vss 0.005299f
C2369 vdd.n2119 vss 0.005299f
C2370 vdd.n2120 vss 0.005299f
C2371 vdd.n2121 vss 0.032171f
C2372 vdd.n2122 vss 0.005299f
C2373 vdd.n2123 vss 0.005299f
C2374 vdd.n2124 vss 0.005299f
C2375 vdd.n2125 vss 0.030582f
C2376 vdd.n2126 vss 0.005299f
C2377 vdd.n2127 vss 0.005299f
C2378 vdd.n2128 vss 0.032171f
C2379 vdd.n2129 vss 0.005299f
C2380 vdd.n2130 vss 0.005299f
C2381 vdd.n2131 vss 0.032171f
C2382 vdd.n2132 vss 0.005299f
C2383 vdd.n2133 vss 0.005299f
C2384 vdd.n2134 vss 0.032171f
C2385 vdd.n2135 vss 0.005299f
C2386 vdd.n2136 vss 0.005299f
C2387 vdd.n2137 vss 0.032171f
C2388 vdd.n2138 vss 0.005299f
C2389 vdd.n2139 vss 0.005299f
C2390 vdd.n2140 vss 0.032171f
C2391 vdd.n2141 vss 0.005299f
C2392 vdd.n2142 vss 0.005299f
C2393 vdd.n2143 vss 0.032171f
C2394 vdd.n2144 vss 0.005299f
C2395 vdd.n2145 vss 0.005299f
C2396 vdd.n2146 vss 0.032567f
C2397 vdd.n2147 vss 0.005299f
C2398 vdd.n2148 vss 0.005299f
C2399 vdd.n2149 vss 0.005299f
C2400 vdd.n2150 vss 0.03098f
C2401 vdd.n2151 vss 0.005299f
C2402 vdd.n2152 vss 0.005299f
C2403 vdd.n2153 vss 0.032171f
C2404 vdd.n2154 vss 0.005299f
C2405 vdd.n2155 vss 0.005299f
C2406 vdd.n2156 vss 0.032171f
C2407 vdd.n2157 vss 0.007009f
C2408 vdd.n2158 vss 0.044334f
C2409 vdd.n2159 vss 0.035336f
C2410 vdd.n2160 vss 0.048562f
C2411 vdd.n2161 vss 0.048863f
C2412 vdd.n2162 vss 0.048863f
C2413 vdd.n2163 vss 0.048562f
C2414 vdd.n2164 vss 0.048863f
C2415 vdd.n2165 vss 0.048562f
C2416 vdd.n2166 vss 0.048562f
C2417 vdd.n2167 vss 0.048562f
C2418 vdd.n2168 vss 0.048562f
C2419 vdd.n2169 vss 0.048863f
C2420 vdd.n2170 vss 0.048562f
C2421 vdd.n2171 vss 0.048562f
C2422 vdd.n2172 vss 0.048863f
C2423 vdd.n2173 vss 0.048863f
C2424 vdd.n2174 vss 0.048562f
C2425 vdd.n2175 vss 0.033766f
C2426 vdd.n2176 vss 0.121953f
C2427 vdd.n2177 vss 0.028305f
C2428 vdd.n2178 vss 0.035117f
C2429 vdd.t319 vss 0.009018f
C2430 vdd.t317 vss 0.008841f
C2431 vdd.n2179 vss 0.171317f
C2432 vdd.t318 vss 0.009018f
C2433 vdd.t316 vss 0.008841f
C2434 vdd.n2180 vss 0.171076f
C2435 vdd.t315 vss 0.008848f
C2436 vdd.t320 vss 0.008848f
C2437 vdd.n2181 vss 0.334604f
C2438 vdd.n2182 vss 0.216612f
C2439 vdd.n2183 vss 0.048748f
C2440 vdd.n2184 vss 0.02735f
C2441 vdd.n2185 vss 0.035117f
C2442 vdd.n2186 vss 0.071272f
C2443 vdd.n2187 vss 0.045584f
C2444 vdd.n2188 vss 0.045584f
C2445 vdd.n2189 vss 4.03e-19
C2446 vdd.n2190 vss 0.045462f
C2447 vdd.n2192 vss 0.045584f
C2448 vdd.n2195 vss 0.045584f
C2449 vdd.n2197 vss 0.045584f
C2450 vdd.n2199 vss 0.028305f
C2451 vdd.n2200 vss 0.017558f
C2452 vdd.n2201 vss 0.022213f
C2453 vdd.n2202 vss 0.064872f
C2454 vdd.n2203 vss 0.045583f
C2455 vdd.n2204 vss 0.02273f
C2456 vdd.n2205 vss 0.061117f
C2457 vdd.n2206 vss 0.017558f
C2458 vdd.n2207 vss 0.081973f
C2459 vdd.n2208 vss 0.035117f
C2460 vdd.n2209 vss 0.02735f
C2461 vdd.n2210 vss 0.121953f
C2462 vdd.n2211 vss 3.1415f
C2463 vdd.n2212 vss 3.14346f
C2464 vdd.n2213 vss 0.028701f
C2465 vdd.n2214 vss 0.02735f
C2466 vdd.n2215 vss 0.048562f
C2467 vdd.n2216 vss 0.048562f
C2468 vdd.n2217 vss 0.048562f
C2469 vdd.n2218 vss 0.048562f
C2470 vdd.n2219 vss 0.048562f
C2471 vdd.n2220 vss 0.048562f
C2472 vdd.n2221 vss 0.062653f
C2473 vdd.n2222 vss 0.048562f
C2474 vdd.n2223 vss 0.123303f
C2475 vdd.n2224 vss 0.028305f
C2476 vdd.n2225 vss 0.035117f
C2477 vdd.n2226 vss 0.048562f
C2478 vdd.n2227 vss 0.048562f
C2479 vdd.n2228 vss 0.035117f
C2480 vdd.n2229 vss 0.02735f
C2481 vdd.n2230 vss 0.120602f
C2482 vdd.n2231 vss 0.024929f
C2483 vdd.n2232 vss 0.16445f
C2484 vdd.n2233 vss 0.027279f
C2485 vdd.n2234 vss 0.048863f
C2486 vdd.n2235 vss 0.048863f
C2487 vdd.n2236 vss 0.048863f
C2488 vdd.n2237 vss 0.048562f
C2489 vdd.n2238 vss 0.048562f
C2490 vdd.n2239 vss 0.048562f
C2491 vdd.n2240 vss 0.048562f
C2492 vdd.n2241 vss 0.048562f
C2493 vdd.n2242 vss 0.048562f
C2494 vdd.n2243 vss 0.048562f
C2495 vdd.n2244 vss 0.048562f
C2496 vdd.n2245 vss 0.048863f
C2497 vdd.n2246 vss 0.048863f
C2498 vdd.n2247 vss 0.048863f
C2499 vdd.n2248 vss 0.048562f
C2500 vdd.n2249 vss 0.046764f
C2501 vdd.n2250 vss 0.048562f
C2502 vdd.n2251 vss 0.048562f
C2503 vdd.n2252 vss 0.02608f
C2504 vdd.n2253 vss 0.048562f
C2505 vdd.n2254 vss 0.044666f
C2506 vdd.n2255 vss 0.048562f
C2507 vdd.n2256 vss 0.048863f
C2508 vdd.n2257 vss 0.028478f
C2509 vdd.n2258 vss 0.048863f
C2510 vdd.n2259 vss 0.042268f
C2511 vdd.n2260 vss 0.048562f
C2512 vdd.n2261 vss 0.048562f
C2513 vdd.n2262 vss 0.030575f
C2514 vdd.n2263 vss 0.048562f
C2515 vdd.n2264 vss 0.040168f
C2516 vdd.n2265 vss 0.048562f
C2517 vdd.n2266 vss 0.048562f
C2518 vdd.n2267 vss 0.032675f
C2519 vdd.n2268 vss 0.048863f
C2520 vdd.n2269 vss 0.038071f
C2521 vdd.n2270 vss 0.048863f
C2522 vdd.n2271 vss 0.048562f
C2523 vdd.n2272 vss 0.035073f
C2524 vdd.n2273 vss 0.048562f
C2525 vdd.n2274 vss 0.035673f
C2526 vdd.n2275 vss 0.048562f
C2527 vdd.n2276 vss 0.048562f
C2528 vdd.n2277 vss 0.037171f
C2529 vdd.n2278 vss 0.048562f
C2530 vdd.n2279 vss 0.033573f
C2531 vdd.n2280 vss 0.048863f
C2532 vdd.n2281 vss 0.048863f
C2533 vdd.n2282 vss 0.039569f
C2534 vdd.n2283 vss 0.048562f
C2535 vdd.n2284 vss 0.031175f
C2536 vdd.n2285 vss 0.048562f
C2537 vdd.n2286 vss 0.048562f
C2538 vdd.n2287 vss 0.041668f
C2539 vdd.n2288 vss 0.048562f
C2540 vdd.n2289 vss 0.029078f
C2541 vdd.n2290 vss 0.048562f
C2542 vdd.n2291 vss 0.048863f
C2543 vdd.n2292 vss 0.048863f
C2544 vdd.n2293 vss 0.048863f
C2545 vdd.n2294 vss 0.026679f
C2546 vdd.n2295 vss 0.238626f
C2547 vdd.n2296 vss 0.046164f
C2548 vdd.n2297 vss 0.048562f
C2549 vdd.n2298 vss 0.048562f
C2550 vdd.n2299 vss 0.048562f
C2551 vdd.n2300 vss 0.02458f
C2552 vdd.n2301 vss 0.238626f
C2553 vdd.n2302 vss 0.048264f
C2554 vdd.n2303 vss 0.046764f
C2555 vdd.n2304 vss 0.048863f
C2556 vdd.n2305 vss 0.048863f
C2557 vdd.n2306 vss 0.026378f
C2558 vdd.n2307 vss 0.028595f
C2559 vdd.n2308 vss 0.032171f
C2560 vdd.n2309 vss 0.005299f
C2561 vdd.n2310 vss 0.005299f
C2562 vdd.n2311 vss 0.032171f
C2563 vdd.n2312 vss 0.005299f
C2564 vdd.n2313 vss 0.005299f
C2565 vdd.n2314 vss 0.028993f
C2566 vdd.n2315 vss 0.031774f
C2567 vdd.n2316 vss 0.005299f
C2568 vdd.n2317 vss 0.004121f
C2569 vdd.n2318 vss 0.032171f
C2570 vdd.n2319 vss 0.004121f
C2571 vdd.n2320 vss 0.002649f
C2572 vdd.n2321 vss 0.450127f
C2573 vdd.n2322 vss 0.182409f
C2574 vdd.n2323 vss 0.182361f
C2575 vdd.n2324 vss 2.47212f
C2576 vdd.n2325 vss 2.60984f
C2577 vdd.n2326 vss 0.182361f
C2578 vdd.n2327 vss 0.063804f
C2579 vdd.n2328 vss 0.006657f
C2580 vdd.n2329 vss 0.034552f
C2581 vdd.n2330 vss 0.002723f
C2582 vdd.n2331 vss 0.013853f
C2583 vdd.n2332 vss 0.012467f
C2584 vdd.n2333 vss 0.027705f
C2585 vdd.n2334 vss 0.027705f
C2586 vdd.n2335 vss 0.027705f
C2587 vdd.n2336 vss 0.027705f
C2588 vdd.n2337 vss 0.027705f
C2589 vdd.n2338 vss 0.027705f
C2590 vdd.n2339 vss 0.108689f
C2591 vdd.n2340 vss 0.013853f
C2592 vdd.n2341 vss 0.027705f
C2593 vdd.n2342 vss 0.094317f
C2594 vdd.n2343 vss 2.14524f
C2595 vdd.n2344 vss 0.017009f
C2596 vdd.n2345 vss 0.00449f
C2597 vdd.n2346 vss 0.034552f
C2598 vdd.n2347 vss 0.004894f
C2599 vdd.n2348 vss 0.013853f
C2600 vdd.n2349 vss 0.012467f
C2601 vdd.n2350 vss 0.027705f
C2602 vdd.t176 vss 0.018831f
C2603 vdd.t303 vss 0.018831f
C2604 vdd.n2351 vss 0.041538f
C2605 vdd.n2352 vss 0.214207f
C2606 vdd.n2353 vss 0.021125f
C2607 vdd.n2354 vss 0.012467f
C2608 vdd.n2355 vss 0.012467f
C2609 vdd.n2356 vss 0.013853f
C2610 vdd.n2357 vss 0.005299f
C2611 vdd.n2358 vss 0.005299f
C2612 vdd.n2359 vss 0.005299f
C2613 vdd.n2360 vss 0.012641f
C2614 vdd.n2361 vss 0.012467f
C2615 vdd.n2362 vss 0.027705f
C2616 vdd.t219 vss 0.018831f
C2617 vdd.t99 vss 0.018831f
C2618 vdd.n2363 vss 0.041538f
C2619 vdd.n2364 vss 0.214207f
C2620 vdd.n2365 vss 0.020433f
C2621 vdd.n2366 vss 0.012467f
C2622 vdd.n2367 vss 0.013853f
C2623 vdd.n2368 vss 0.005299f
C2624 vdd.n2369 vss 0.005299f
C2625 vdd.n2370 vss 0.013853f
C2626 vdd.n2371 vss 0.012467f
C2627 vdd.n2372 vss 0.027705f
C2628 vdd.t105 vss 0.018831f
C2629 vdd.t243 vss 0.018831f
C2630 vdd.n2373 vss 0.041538f
C2631 vdd.n2374 vss 0.214207f
C2632 vdd.n2375 vss 0.01974f
C2633 vdd.n2376 vss 0.012467f
C2634 vdd.n2377 vss 0.013853f
C2635 vdd.n2378 vss 0.005299f
C2636 vdd.n2379 vss 0.005299f
C2637 vdd.n2380 vss 0.013853f
C2638 vdd.n2381 vss 0.012467f
C2639 vdd.n2382 vss 0.027705f
C2640 vdd.t43 vss 0.018831f
C2641 vdd.t264 vss 0.018831f
C2642 vdd.n2383 vss 0.041538f
C2643 vdd.n2384 vss 0.214207f
C2644 vdd.n2385 vss 0.019047f
C2645 vdd.n2386 vss 0.012467f
C2646 vdd.n2387 vss 0.012467f
C2647 vdd.n2388 vss 0.013853f
C2648 vdd.n2389 vss 0.005299f
C2649 vdd.n2390 vss 0.005299f
C2650 vdd.n2391 vss 0.005299f
C2651 vdd.n2392 vss 0.012641f
C2652 vdd.n2393 vss 0.012467f
C2653 vdd.n2394 vss 0.027705f
C2654 vdd.t159 vss 0.018831f
C2655 vdd.t49 vss 0.018831f
C2656 vdd.n2395 vss 0.041538f
C2657 vdd.n2396 vss 0.214207f
C2658 vdd.n2397 vss 0.018355f
C2659 vdd.n2398 vss 0.012467f
C2660 vdd.n2399 vss 0.013853f
C2661 vdd.n2400 vss 0.005299f
C2662 vdd.n2401 vss 0.005299f
C2663 vdd.n2402 vss 0.013853f
C2664 vdd.n2403 vss 0.012467f
C2665 vdd.n2404 vss 0.027705f
C2666 vdd.t188 vss 0.018831f
C2667 vdd.t307 vss 0.018831f
C2668 vdd.n2405 vss 0.041538f
C2669 vdd.n2406 vss 0.214207f
C2670 vdd.n2407 vss 0.017662f
C2671 vdd.n2408 vss 0.012467f
C2672 vdd.n2409 vss 0.013853f
C2673 vdd.n2410 vss 0.005299f
C2674 vdd.n2411 vss 0.003238f
C2675 vdd.n2412 vss 0.005299f
C2676 vdd.n2413 vss 0.013853f
C2677 vdd.n2414 vss 0.012467f
C2678 vdd.n2415 vss 0.027705f
C2679 vdd.t310 vss 0.018831f
C2680 vdd.t231 vss 0.018831f
C2681 vdd.n2416 vss 0.041538f
C2682 vdd.n2417 vss 0.214207f
C2683 vdd.n2418 vss 0.01697f
C2684 vdd.n2419 vss 0.012467f
C2685 vdd.n2420 vss 0.012467f
C2686 vdd.n2421 vss 0.013853f
C2687 vdd.n2422 vss 0.00471f
C2688 vdd.n2423 vss 0.005299f
C2689 vdd.n2424 vss 0.005299f
C2690 vdd.n2425 vss 0.012641f
C2691 vdd.n2426 vss 0.012467f
C2692 vdd.n2427 vss 0.027705f
C2693 vdd.t115 vss 0.018831f
C2694 vdd.t312 vss 0.018831f
C2695 vdd.n2428 vss 0.041538f
C2696 vdd.n2429 vss 0.214207f
C2697 vdd.n2430 vss 0.016277f
C2698 vdd.n2431 vss 0.012467f
C2699 vdd.n2432 vss 0.013853f
C2700 vdd.n2433 vss 0.005299f
C2701 vdd.n2434 vss 0.005299f
C2702 vdd.n2435 vss 0.013853f
C2703 vdd.n2436 vss 0.012467f
C2704 vdd.n2437 vss 0.027705f
C2705 vdd.t53 vss 0.018831f
C2706 vdd.t266 vss 0.018831f
C2707 vdd.n2438 vss 0.041538f
C2708 vdd.n2439 vss 0.214207f
C2709 vdd.n2440 vss 0.015584f
C2710 vdd.n2441 vss 0.012467f
C2711 vdd.n2442 vss 0.013853f
C2712 vdd.n2443 vss 0.005299f
C2713 vdd.n2444 vss 0.005299f
C2714 vdd.n2445 vss 0.013853f
C2715 vdd.n2446 vss 0.012467f
C2716 vdd.n2447 vss 0.027705f
C2717 vdd.t163 vss 0.018831f
C2718 vdd.t57 vss 0.018831f
C2719 vdd.n2448 vss 0.041538f
C2720 vdd.n2449 vss 0.214207f
C2721 vdd.n2450 vss 0.014892f
C2722 vdd.n2451 vss 0.012467f
C2723 vdd.n2452 vss 0.012467f
C2724 vdd.n2453 vss 0.013853f
C2725 vdd.n2454 vss 0.005299f
C2726 vdd.n2455 vss 0.005299f
C2727 vdd.n2456 vss 0.005299f
C2728 vdd.n2457 vss 0.012641f
C2729 vdd.n2458 vss 0.012467f
C2730 vdd.n2459 vss 0.027705f
C2731 vdd.t268 vss 0.018831f
C2732 vdd.t202 vss 0.018831f
C2733 vdd.n2460 vss 0.041538f
C2734 vdd.n2461 vss 0.214207f
C2735 vdd.n2462 vss 0.014199f
C2736 vdd.n2463 vss 0.012467f
C2737 vdd.n2464 vss 0.013853f
C2738 vdd.n2465 vss 0.005299f
C2739 vdd.n2466 vss 0.005299f
C2740 vdd.n2467 vss 0.013853f
C2741 vdd.n2468 vss 0.012467f
C2742 vdd.n2469 vss 0.027359f
C2743 vdd.n2470 vss 0.214207f
C2744 vdd.n2471 vss 0.014199f
C2745 vdd.n2472 vss 0.012467f
C2746 vdd.n2473 vss 0.013853f
C2747 vdd.n2474 vss 0.005299f
C2748 vdd.n2475 vss 0.005299f
C2749 vdd.n2476 vss 0.013853f
C2750 vdd.n2477 vss 0.012467f
C2751 vdd.n2478 vss 0.026666f
C2752 vdd.n2479 vss 0.230968f
C2753 vdd.n2480 vss 0.023729f
C2754 vdd.n2481 vss 0.039118f
C2755 vdd.n2482 vss 0.070093f
C2756 vdd.n2483 vss 0.182361f
C2757 vdd.n2484 vss 2.95042f
C2758 vdd.n2485 vss 2.64283f
C2759 vdd.t133 vss 0.416023f
C2760 vdd.t269 vss 0.337394f
C2761 vdd.t169 vss 0.337394f
C2762 vdd.t291 vss 0.337394f
C2763 vdd.t203 vss 0.337394f
C2764 vdd.t124 vss 0.337394f
C2765 vdd.t185 vss 0.337394f
C2766 vdd.t4 vss 0.241607f
C2767 vdd.t246 vss 0.337394f
C2768 vdd.t223 vss 0.337394f
C2769 vdd.t8 vss 0.337394f
C2770 vdd.t122 vss 0.337394f
C2771 vdd.t288 vss 0.337394f
C2772 vdd.t183 vss 0.416023f
C2773 vdd.n2486 vss 0.033043f
C2774 vdd.n2487 vss 0.033043f
C2775 vdd.n2488 vss 0.494652f
C2776 vdd.t254 vss 0.416023f
C2777 vdd.t18 vss 0.337394f
C2778 vdd.t116 vss 0.337394f
C2779 vdd.t293 vss 0.337394f
C2780 vdd.t74 vss 0.337394f
C2781 vdd.t196 vss 0.337394f
C2782 vdd.t281 vss 0.337394f
C2783 vdd.n2489 vss 0.036165f
C2784 vdd.n2490 vss 0.049464f
C2785 vdd.n2491 vss 0.005299f
C2786 vdd.n2492 vss 0.006859f
C2787 vdd.n2493 vss 0.030896f
C2788 vdd.n2494 vss 0.006859f
C2789 vdd.n2495 vss 0.005299f
C2790 vdd.n2496 vss 0.005299f
C2791 vdd.n2497 vss 0.005299f
C2792 vdd.n2498 vss 0.005299f
C2793 vdd.n2499 vss 0.005299f
C2794 vdd.n2500 vss 0.005299f
C2795 vdd.t134 vss 0.018831f
C2796 vdd.t270 vss 0.018831f
C2797 vdd.n2501 vss 0.039834f
C2798 vdd.n2502 vss 0.137733f
C2799 vdd.n2503 vss 0.005299f
C2800 vdd.n2504 vss 0.005299f
C2801 vdd.n2505 vss 0.005299f
C2802 vdd.n2506 vss 0.005299f
C2803 vdd.n2507 vss 0.005299f
C2804 vdd.n2508 vss 0.005299f
C2805 vdd.n2509 vss 0.005299f
C2806 vdd.n2510 vss 0.005299f
C2807 vdd.n2511 vss 0.005299f
C2808 vdd.n2512 vss 0.005299f
C2809 vdd.n2513 vss 0.005299f
C2810 vdd.n2514 vss 0.028519f
C2811 vdd.n2515 vss 0.005299f
C2812 vdd.n2516 vss 0.005299f
C2813 vdd.n2517 vss 0.005299f
C2814 vdd.n2518 vss 0.005299f
C2815 vdd.n2519 vss 0.005299f
C2816 vdd.t204 vss 0.018831f
C2817 vdd.t125 vss 0.018831f
C2818 vdd.n2520 vss 0.039834f
C2819 vdd.n2521 vss 0.005299f
C2820 vdd.n2522 vss 0.005299f
C2821 vdd.n2523 vss 0.005299f
C2822 vdd.n2524 vss 0.022974f
C2823 vdd.n2525 vss 0.032084f
C2824 vdd.n2526 vss 0.005299f
C2825 vdd.n2527 vss 0.005299f
C2826 vdd.n2528 vss 0.005299f
C2827 vdd.n2529 vss 0.005299f
C2828 vdd.n2530 vss 0.03248f
C2829 vdd.n2531 vss 0.005299f
C2830 vdd.n2532 vss 0.005299f
C2831 vdd.n2533 vss 0.01624f
C2832 vdd.n2534 vss 0.143675f
C2833 vdd.n2535 vss 0.015844f
C2834 vdd.n2536 vss 0.005299f
C2835 vdd.n2537 vss 0.005299f
C2836 vdd.n2538 vss 0.032084f
C2837 vdd.n2539 vss 0.005299f
C2838 vdd.n2540 vss 0.005299f
C2839 vdd.n2541 vss 0.032084f
C2840 vdd.n2542 vss 0.005299f
C2841 vdd.n2543 vss 0.005299f
C2842 vdd.t170 vss 0.018831f
C2843 vdd.t292 vss 0.018831f
C2844 vdd.n2544 vss 0.039834f
C2845 vdd.n2545 vss 0.135753f
C2846 vdd.n2546 vss 0.018617f
C2847 vdd.n2547 vss 0.005299f
C2848 vdd.n2548 vss 0.005299f
C2849 vdd.n2549 vss 0.032084f
C2850 vdd.n2550 vss 0.005299f
C2851 vdd.n2551 vss 0.005299f
C2852 vdd.n2552 vss 0.032084f
C2853 vdd.n2553 vss 0.028519f
C2854 vdd.n2554 vss 0.010695f
C2855 vdd.n2555 vss 0.005299f
C2856 vdd.n2556 vss 0.005299f
C2857 vdd.n2557 vss 0.032084f
C2858 vdd.n2558 vss 0.005299f
C2859 vdd.n2559 vss 0.005299f
C2860 vdd.n2560 vss 0.006859f
C2861 vdd.n2561 vss 0.029707f
C2862 vdd.n2562 vss 0.003312f
C2863 vdd.n2563 vss 0.02088f
C2864 vdd.n2564 vss 0.070665f
C2865 vdd.n2565 vss 0.090428f
C2866 vdd.n2566 vss 0.090428f
C2867 vdd.t164 vss 0.337394f
C2868 vdd.n2567 vss 0.090428f
C2869 vdd.n2568 vss 0.002649f
C2870 vdd.n2569 vss 0.004305f
C2871 vdd.n2570 vss 0.019409f
C2872 vdd.n2571 vss 0.005299f
C2873 vdd.n2572 vss 0.005299f
C2874 vdd.n2573 vss 0.032084f
C2875 vdd.n2574 vss 0.005299f
C2876 vdd.n2575 vss 0.005299f
C2877 vdd.n2576 vss 0.032084f
C2878 vdd.n2577 vss 0.005299f
C2879 vdd.n2578 vss 0.005299f
C2880 vdd.t282 vss 0.018831f
C2881 vdd.t197 vss 0.018831f
C2882 vdd.n2579 vss 0.039834f
C2883 vdd.n2580 vss 0.139714f
C2884 vdd.n2581 vss 0.009902f
C2885 vdd.n2582 vss 0.005299f
C2886 vdd.n2583 vss 0.005299f
C2887 vdd.n2584 vss 0.032084f
C2888 vdd.n2585 vss 0.005299f
C2889 vdd.n2586 vss 0.005299f
C2890 vdd.n2587 vss 0.005299f
C2891 vdd.n2588 vss 0.032084f
C2892 vdd.n2589 vss 0.005299f
C2893 vdd.n2590 vss 0.005299f
C2894 vdd.n2591 vss 0.02535f
C2895 vdd.n2592 vss 0.005299f
C2896 vdd.n2593 vss 0.005299f
C2897 vdd.n2594 vss 0.032084f
C2898 vdd.n2595 vss 0.005299f
C2899 vdd.n2596 vss 0.005299f
C2900 vdd.n2597 vss 0.032084f
C2901 vdd.n2598 vss 0.005299f
C2902 vdd.n2599 vss 0.005299f
C2903 vdd.n2600 vss 0.028123f
C2904 vdd.n2601 vss 0.005299f
C2905 vdd.n2602 vss 0.005299f
C2906 vdd.n2603 vss 0.032084f
C2907 vdd.n2604 vss 0.005299f
C2908 vdd.n2605 vss 0.005299f
C2909 vdd.n2606 vss 0.032084f
C2910 vdd.n2607 vss 0.005299f
C2911 vdd.n2608 vss 0.005299f
C2912 vdd.n2609 vss 0.005299f
C2913 vdd.n2610 vss 0.028915f
C2914 vdd.n2611 vss 0.005299f
C2915 vdd.n2612 vss 0.005299f
C2916 vdd.n2613 vss 0.032084f
C2917 vdd.n2614 vss 0.003974f
C2918 vdd.n2615 vss 0.005299f
C2919 vdd.n2616 vss 0.032084f
C2920 vdd.n2617 vss 0.005299f
C2921 vdd.n2618 vss 0.005299f
C2922 vdd.n2619 vss 0.032084f
C2923 vdd.n2620 vss 0.005299f
C2924 vdd.n2621 vss 0.005299f
C2925 vdd.n2622 vss 0.022578f
C2926 vdd.n2623 vss 0.005299f
C2927 vdd.n2624 vss 0.005299f
C2928 vdd.n2625 vss 0.032084f
C2929 vdd.n2626 vss 0.005299f
C2930 vdd.n2627 vss 0.005299f
C2931 vdd.n2628 vss 0.032084f
C2932 vdd.n2629 vss 0.005299f
C2933 vdd.n2630 vss 0.005299f
C2934 vdd.n2631 vss 0.147636f
C2935 vdd.n2632 vss 0.005299f
C2936 vdd.n2633 vss 0.005299f
C2937 vdd.n2634 vss 0.005299f
C2938 vdd.n2635 vss 0.029311f
C2939 vdd.n2636 vss 0.005299f
C2940 vdd.n2637 vss 0.005299f
C2941 vdd.n2638 vss 0.032084f
C2942 vdd.n2639 vss 0.005299f
C2943 vdd.n2640 vss 0.005299f
C2944 vdd.n2641 vss 0.028519f
C2945 vdd.n2642 vss 0.005299f
C2946 vdd.n2643 vss 0.005299f
C2947 vdd.n2644 vss 0.032084f
C2948 vdd.n2645 vss 0.005299f
C2949 vdd.n2646 vss 0.003827f
C2950 vdd.n2647 vss 0.032084f
C2951 vdd.n2648 vss 0.003827f
C2952 vdd.n2649 vss -0.21879f
C2953 vdd.n2650 vss 0.004121f
C2954 vdd.n2651 vss 0.031292f
C2955 vdd.n2652 vss 0.004121f
C2956 vdd.n2653 vss 0.005299f
C2957 vdd.n2654 vss 0.005299f
C2958 vdd.t69 vss 0.018831f
C2959 vdd.t284 vss 0.018831f
C2960 vdd.n2655 vss 0.039834f
C2961 vdd.n2656 vss 0.141298f
C2962 vdd.n2657 vss 0.005299f
C2963 vdd.n2658 vss 0.004753f
C2964 vdd.n2659 vss 0.005299f
C2965 vdd.n2660 vss 0.005299f
C2966 vdd.n2661 vss 0.005299f
C2967 vdd.n2662 vss 0.005299f
C2968 vdd.n2663 vss 0.005299f
C2969 vdd.n2664 vss 0.005299f
C2970 vdd.n2665 vss 0.005299f
C2971 vdd.n2666 vss 0.005299f
C2972 vdd.n2667 vss 0.005299f
C2973 vdd.n2668 vss 0.005299f
C2974 vdd.n2669 vss 0.005299f
C2975 vdd.n2670 vss 0.028519f
C2976 vdd.n2671 vss 0.005299f
C2977 vdd.n2672 vss 0.005299f
C2978 vdd.n2673 vss 0.005299f
C2979 vdd.n2674 vss 0.005299f
C2980 vdd.n2675 vss 0.005299f
C2981 vdd.n2676 vss 0.005299f
C2982 vdd.n2677 vss 0.005299f
C2983 vdd.n2678 vss 0.005299f
C2984 vdd.n2679 vss 0.028519f
C2985 vdd.n2680 vss 0.005299f
C2986 vdd.n2681 vss 0.005299f
C2987 vdd.n2682 vss 0.005299f
C2988 vdd.t21 vss 0.070922f
C2989 vdd.n2683 vss 0.005299f
C2990 vdd.n2684 vss 0.005299f
C2991 vdd.n2685 vss 0.019171f
C2992 vdd.n2686 vss 0.005299f
C2993 vdd.n2687 vss 0.005299f
C2994 vdd.n2688 vss 0.005299f
C2995 vdd.n2689 vss 0.005299f
C2996 vdd.n2690 vss 0.005299f
C2997 vdd.n2691 vss 0.005299f
C2998 vdd.n2692 vss 0.028519f
C2999 vdd.n2693 vss 0.005299f
C3000 vdd.n2694 vss 0.005299f
C3001 vdd.n2695 vss 0.005299f
C3002 vdd.t182 vss 0.018831f
C3003 vdd.t3 vss 0.018831f
C3004 vdd.n2696 vss 0.040001f
C3005 vdd.n2697 vss 0.127877f
C3006 vdd.n2698 vss 0.005299f
C3007 vdd.n2699 vss 0.005299f
C3008 vdd.n2700 vss 0.005299f
C3009 vdd.n2701 vss 0.005299f
C3010 vdd.n2702 vss 0.005299f
C3011 vdd.n2703 vss 0.005299f
C3012 vdd.t242 vss 0.018831f
C3013 vdd.t127 vss 0.018831f
C3014 vdd.n2704 vss 0.039834f
C3015 vdd.n2705 vss 0.14209f
C3016 vdd.n2706 vss 0.005299f
C3017 vdd.n2707 vss 0.00713f
C3018 vdd.n2708 vss 0.005299f
C3019 vdd.n2709 vss 0.005299f
C3020 vdd.n2710 vss 0.005299f
C3021 vdd.n2711 vss 0.005299f
C3022 vdd.n2712 vss 0.005299f
C3023 vdd.n2713 vss 0.005299f
C3024 vdd.n2714 vss 0.005299f
C3025 vdd.n2715 vss 0.005299f
C3026 vdd.n2716 vss 0.005299f
C3027 vdd.n2717 vss 0.005299f
C3028 vdd.n2718 vss 0.005299f
C3029 vdd.n2719 vss 0.028519f
C3030 vdd.n2720 vss 0.005299f
C3031 vdd.t161 vss 0.018831f
C3032 vdd.t279 vss 0.018831f
C3033 vdd.n2721 vss 0.040001f
C3034 vdd.n2722 vss 0.131838f
C3035 vdd.n2723 vss 0.020597f
C3036 vdd.n2724 vss 0.005299f
C3037 vdd.n2725 vss 0.005299f
C3038 vdd.n2726 vss 0.005299f
C3039 vdd.n2727 vss 0.032084f
C3040 vdd.n2728 vss 0.005299f
C3041 vdd.n2729 vss 0.005299f
C3042 vdd.n2730 vss 0.03248f
C3043 vdd.n2731 vss 0.005299f
C3044 vdd.n2732 vss 0.005299f
C3045 vdd.t11 vss 0.018831f
C3046 vdd.t15 vss 0.018831f
C3047 vdd.n2733 vss 0.039834f
C3048 vdd.n2734 vss 0.124266f
C3049 vdd.n2735 vss 0.023766f
C3050 vdd.n2736 vss 0.005299f
C3051 vdd.n2737 vss 0.005299f
C3052 vdd.n2738 vss 0.032084f
C3053 vdd.n2739 vss 0.005299f
C3054 vdd.n2740 vss 0.005299f
C3055 vdd.n2741 vss 0.0305f
C3056 vdd.n2742 vss 0.030104f
C3057 vdd.n2743 vss 0.005299f
C3058 vdd.n2744 vss 0.005299f
C3059 vdd.n2745 vss 0.026539f
C3060 vdd.n2746 vss 0.005299f
C3061 vdd.n2747 vss 0.005299f
C3062 vdd.n2748 vss 0.032084f
C3063 vdd.n2749 vss 0.005299f
C3064 vdd.n2750 vss 0.005299f
C3065 vdd.n2751 vss 0.032084f
C3066 vdd.n2752 vss 0.005299f
C3067 vdd.n2753 vss 0.005299f
C3068 vdd.n2754 vss 0.029707f
C3069 vdd.n2755 vss 0.005299f
C3070 vdd.n2756 vss 0.005299f
C3071 vdd.n2757 vss 0.032084f
C3072 vdd.n2758 vss 0.005299f
C3073 vdd.n2759 vss 0.004636f
C3074 vdd.n2760 vss 0.032084f
C3075 vdd.n2761 vss 0.005299f
C3076 vdd.n2762 vss 0.005299f
C3077 vdd.n2763 vss 0.032084f
C3078 vdd.n2764 vss 0.003312f
C3079 vdd.n2765 vss 0.005299f
C3080 vdd.n2766 vss 0.011091f
C3081 vdd.n2767 vss 0.150248f
C3082 vdd.n2768 vss 0.020993f
C3083 vdd.n2769 vss 0.005299f
C3084 vdd.n2770 vss 0.005299f
C3085 vdd.n2771 vss 0.032084f
C3086 vdd.n2772 vss 0.005299f
C3087 vdd.n2773 vss 0.005299f
C3088 vdd.n2774 vss 0.032084f
C3089 vdd.n2775 vss 0.005299f
C3090 vdd.n2776 vss 0.005299f
C3091 vdd.t131 vss 0.018831f
C3092 vdd.t137 vss 0.018831f
C3093 vdd.n2777 vss 0.039834f
C3094 vdd.n2778 vss 0.134564f
C3095 vdd.n2779 vss 0.024162f
C3096 vdd.n2780 vss 0.005299f
C3097 vdd.n2781 vss 0.005299f
C3098 vdd.n2782 vss 0.032084f
C3099 vdd.n2783 vss 0.005299f
C3100 vdd.n2784 vss 0.005299f
C3101 vdd.n2785 vss 0.032084f
C3102 vdd.n2786 vss 0.005299f
C3103 vdd.n2787 vss 0.005299f
C3104 vdd.t199 vss 0.018831f
C3105 vdd.t77 vss 0.018831f
C3106 vdd.n2788 vss 0.039834f
C3107 vdd.n2789 vss 0.123474f
C3108 vdd.n2790 vss 0.026935f
C3109 vdd.n2791 vss 0.005299f
C3110 vdd.n2792 vss 0.005299f
C3111 vdd.n2793 vss 0.032084f
C3112 vdd.n2794 vss 0.005299f
C3113 vdd.n2795 vss 0.005299f
C3114 vdd.n2796 vss 0.029707f
C3115 vdd.n2797 vss 0.030896f
C3116 vdd.n2798 vss 0.005299f
C3117 vdd.n2799 vss 0.005299f
C3118 vdd.n2800 vss 0.029707f
C3119 vdd.n2801 vss 0.005299f
C3120 vdd.n2802 vss 0.005299f
C3121 vdd.n2803 vss 0.03248f
C3122 vdd.n2804 vss 0.004305f
C3123 vdd.n2805 vss 0.002649f
C3124 vdd.n2806 vss 0.073519f
C3125 vdd.t191 vss 0.264482f
C3126 vdd.n2807 vss 0.073519f
C3127 vdd.n2808 vss 0.073519f
C3128 vdd.n2809 vss 0.09004f
C3129 vdd.n2810 vss 0.022898f
C3130 vdd.n2811 vss 0.073487f
C3131 vdd.n2812 vss 0.090428f
C3132 vdd.n2813 vss 0.090428f
C3133 vdd.t278 vss 0.337394f
C3134 vdd.n2814 vss 0.090428f
C3135 vdd.n2815 vss 0.002649f
C3136 vdd.n2816 vss 0.00298f
C3137 vdd.n2817 vss 0.032084f
C3138 vdd.n2818 vss 0.005299f
C3139 vdd.n2819 vss 0.005299f
C3140 vdd.n2820 vss 0.032084f
C3141 vdd.n2821 vss 0.005299f
C3142 vdd.n2822 vss 0.005299f
C3143 vdd.n2823 vss 0.017824f
C3144 vdd.n2824 vss 0.005299f
C3145 vdd.n2825 vss 0.005299f
C3146 vdd.n2826 vss 0.01426f
C3147 vdd.n2827 vss 0.005299f
C3148 vdd.n2828 vss 0.005299f
C3149 vdd.n2829 vss 0.032084f
C3150 vdd.n2830 vss 0.005299f
C3151 vdd.n2831 vss 0.005299f
C3152 vdd.n2832 vss 0.03248f
C3153 vdd.n2833 vss 0.005299f
C3154 vdd.n2834 vss 0.005299f
C3155 vdd.n2835 vss 0.017428f
C3156 vdd.n2836 vss 0.005299f
C3157 vdd.n2837 vss 0.005299f
C3158 vdd.n2838 vss 0.032084f
C3159 vdd.n2839 vss 0.005299f
C3160 vdd.n2840 vss 0.005299f
C3161 vdd.n2841 vss 0.032084f
C3162 vdd.n2842 vss 0.005299f
C3163 vdd.n2843 vss 0.005299f
C3164 vdd.t249 vss 0.018831f
C3165 vdd.t253 vss 0.018831f
C3166 vdd.n2844 vss 0.039834f
C3167 vdd.n2845 vss 0.139318f
C3168 vdd.n2846 vss 0.011883f
C3169 vdd.n2847 vss 0.005299f
C3170 vdd.n2848 vss 0.005299f
C3171 vdd.n2849 vss 0.005299f
C3172 vdd.n2850 vss 0.032084f
C3173 vdd.n2851 vss 0.005299f
C3174 vdd.n2852 vss 0.005299f
C3175 vdd.n2853 vss 0.007009f
C3176 vdd.n2854 vss 0.031292f
C3177 vdd.t139 vss 0.070922f
C3178 vdd.n2855 vss 0.147475f
C3179 vdd.n2856 vss 0.011883f
C3180 vdd.n2857 vss 0.145367f
C3181 vdd.n2858 vss 1.40899f
C3182 vdd.n2859 vss 1.12054f
C3183 vdd.n2860 vss 0.048562f
C3184 vdd.n2861 vss 0.048562f
C3185 vdd.n2862 vss 0.048562f
C3186 vdd.n2863 vss 0.048562f
C3187 vdd.n2864 vss 0.048562f
C3188 vdd.n2865 vss 0.048562f
C3189 vdd.n2866 vss 0.048863f
C3190 vdd.n2867 vss 0.048863f
C3191 vdd.n2868 vss 0.048863f
C3192 vdd.n2869 vss 0.048562f
C3193 vdd.n2870 vss 0.048562f
C3194 vdd.n2871 vss 0.048562f
C3195 vdd.n2872 vss 0.048562f
C3196 vdd.n2873 vss 0.048562f
C3197 vdd.n2874 vss 0.048562f
C3198 vdd.n2875 vss 0.048562f
C3199 vdd.n2876 vss 0.048562f
C3200 vdd.n2877 vss 0.048863f
C3201 vdd.n2878 vss 0.048863f
C3202 vdd.n2879 vss 0.048863f
C3203 vdd.n2880 vss 0.048562f
C3204 vdd.n2881 vss 0.048562f
C3205 vdd.n2882 vss 0.048562f
C3206 vdd.n2883 vss 0.048562f
C3207 vdd.n2884 vss 0.048562f
C3208 vdd.n2885 vss 0.048562f
C3209 vdd.n2886 vss 0.048562f
C3210 vdd.n2887 vss 0.048863f
C3211 vdd.n2888 vss 0.048863f
C3212 vdd.n2889 vss 0.048863f
C3213 vdd.n2890 vss 0.048562f
C3214 vdd.n2891 vss 0.048562f
C3215 vdd.n2892 vss 0.048562f
C3216 vdd.n2893 vss 0.048562f
C3217 vdd.n2894 vss 0.048562f
C3218 vdd.n2895 vss 0.048562f
C3219 vdd.n2896 vss 0.048562f
C3220 vdd.n2897 vss 0.048562f
C3221 vdd.n2898 vss 0.048863f
C3222 vdd.n2899 vss 0.048863f
C3223 vdd.n2900 vss 0.048863f
C3224 vdd.n2901 vss 0.048562f
C3225 vdd.n2902 vss 0.048562f
C3226 vdd.n2903 vss 0.048562f
C3227 vdd.n2904 vss 0.048562f
C3228 vdd.n2905 vss 0.048562f
C3229 vdd.n2906 vss 0.048562f
C3230 vdd.n2907 vss 0.048562f
C3231 vdd.n2908 vss 0.048863f
C3232 vdd.n2909 vss 0.048863f
C3233 vdd.n2910 vss 0.048863f
C3234 vdd.n2911 vss 0.048562f
C3235 vdd.n2912 vss 0.048562f
C3236 vdd.n2913 vss 0.048562f
C3237 vdd.n2914 vss 0.048562f
C3238 vdd.n2915 vss 0.048562f
C3239 vdd.n2916 vss 0.048562f
C3240 vdd.n2917 vss 0.048562f
C3241 vdd.n2918 vss 0.048562f
C3242 vdd.n2919 vss 0.048863f
C3243 vdd.n2920 vss 0.048863f
C3244 vdd.n2921 vss 0.048863f
C3245 vdd.n2922 vss 0.048562f
C3246 vdd.n2923 vss 0.048562f
C3247 vdd.n2924 vss 0.048562f
C3248 vdd.n2925 vss 0.048562f
C3249 vdd.n2926 vss 0.048562f
C3250 vdd.n2927 vss 0.048562f
C3251 vdd.n2928 vss 0.048562f
C3252 vdd.n2929 vss 0.048863f
C3253 vdd.n2930 vss 0.048863f
C3254 vdd.n2931 vss 0.048863f
C3255 vdd.n2932 vss 0.048562f
C3256 vdd.n2933 vss 0.048562f
C3257 vdd.n2934 vss 0.048562f
C3258 vdd.n2935 vss 0.048562f
C3259 vdd.n2936 vss 0.048562f
C3260 vdd.n2937 vss 0.048562f
C3261 vdd.n2938 vss 0.048562f
C3262 vdd.n2939 vss 0.048562f
C3263 vdd.n2940 vss 0.048863f
C3264 vdd.n2941 vss 0.048863f
C3265 vdd.n2942 vss 0.048863f
C3266 vdd.n2943 vss 0.048562f
C3267 vdd.n2944 vss 0.048562f
C3268 vdd.n2945 vss 0.048562f
C3269 vdd.n2946 vss 0.048562f
C3270 vdd.n2947 vss 0.048562f
C3271 vdd.n2948 vss 0.048562f
C3272 vdd.n2949 vss 0.048562f
C3273 vdd.n2950 vss 0.048863f
C3274 vdd.n2951 vss 0.048863f
C3275 vdd.n2952 vss 0.048863f
C3276 vdd.n2953 vss 0.048562f
C3277 vdd.n2954 vss 0.048562f
C3278 vdd.n2955 vss 0.048562f
C3279 vdd.n2956 vss 0.048562f
C3280 vdd.n2957 vss 0.048562f
C3281 vdd.n2958 vss 0.048562f
C3282 vdd.n2959 vss 0.048562f
C3283 vdd.n2960 vss 0.048562f
C3284 vdd.n2961 vss 0.048863f
C3285 vdd.n2962 vss 0.048863f
C3286 vdd.n2963 vss 0.048863f
C3287 vdd.n2964 vss 0.048562f
C3288 vdd.n2965 vss 0.048562f
C3289 vdd.n2966 vss 0.048562f
C3290 vdd.n2967 vss 0.048562f
C3291 vdd.n2968 vss 0.048562f
C3292 vdd.n2969 vss 0.048562f
C3293 vdd.n2970 vss 0.048562f
C3294 vdd.n2971 vss 0.062653f
C3295 vdd.n2972 vss 0.037171f
C3296 vdd.n2973 vss 0.047887f
C3297 iref.t15 vss 0.044102f
C3298 iref.t25 vss 0.044102f
C3299 iref.n0 vss 0.096489f
C3300 iref.t1 vss 0.044102f
C3301 iref.t19 vss 0.044102f
C3302 iref.n1 vss 0.096489f
C3303 iref.t17 vss 0.044102f
C3304 iref.t9 vss 0.044102f
C3305 iref.n2 vss 0.096489f
C3306 iref.t7 vss 0.044102f
C3307 iref.t5 vss 0.044102f
C3308 iref.n3 vss 0.096489f
C3309 iref.t27 vss 0.044102f
C3310 iref.t21 vss 0.044102f
C3311 iref.n4 vss 0.096489f
C3312 iref.t23 vss 0.044102f
C3313 iref.t11 vss 0.044102f
C3314 iref.n5 vss 0.096489f
C3315 iref.t3 vss 0.044102f
C3316 iref.t13 vss 0.044102f
C3317 iref.n6 vss 0.096489f
C3318 iref.t29 vss 0.168976f
C3319 iref.t58 vss 0.158044f
C3320 iref.t108 vss 0.158044f
C3321 iref.n7 vss 0.174251f
C3322 iref.t117 vss 0.158044f
C3323 iref.t172 vss 0.158044f
C3324 iref.n8 vss 0.170249f
C3325 iref.n9 vss 0.209101f
C3326 iref.t35 vss 0.158044f
C3327 iref.t90 vss 0.158044f
C3328 iref.n10 vss 0.170249f
C3329 iref.n11 vss 0.103482f
C3330 iref.t152 vss 0.158044f
C3331 iref.t202 vss 0.158044f
C3332 iref.n12 vss 0.170249f
C3333 iref.n13 vss 0.103482f
C3334 iref.t206 vss 0.158044f
C3335 iref.t79 vss 0.158044f
C3336 iref.n14 vss 0.170249f
C3337 iref.n15 vss 0.103482f
C3338 iref.t84 vss 0.158044f
C3339 iref.t143 vss 0.158044f
C3340 iref.n16 vss 0.170249f
C3341 iref.n17 vss 0.103482f
C3342 iref.t82 vss 0.158044f
C3343 iref.t139 vss 0.158044f
C3344 iref.n18 vss 0.170249f
C3345 iref.n19 vss 0.103482f
C3346 iref.t185 vss 0.158044f
C3347 iref.t61 vss 0.158044f
C3348 iref.n20 vss 0.170249f
C3349 iref.n21 vss 0.103482f
C3350 iref.t114 vss 0.158044f
C3351 iref.t169 vss 0.158044f
C3352 iref.n22 vss 0.170249f
C3353 iref.n23 vss 0.103482f
C3354 iref.t177 vss 0.158044f
C3355 iref.t45 vss 0.158044f
C3356 iref.n24 vss 0.170249f
C3357 iref.n25 vss 0.103482f
C3358 iref.t54 vss 0.158044f
C3359 iref.t102 vss 0.158044f
C3360 iref.n26 vss 0.170249f
C3361 iref.n27 vss 0.103482f
C3362 iref.t111 vss 0.158044f
C3363 iref.t166 vss 0.158044f
C3364 iref.n28 vss 0.170249f
C3365 iref.n29 vss 0.103482f
C3366 iref.t173 vss 0.158044f
C3367 iref.t43 vss 0.158044f
C3368 iref.n30 vss 0.170249f
C3369 iref.n31 vss 0.103482f
C3370 iref.t148 vss 0.158044f
C3371 iref.t197 vss 0.158044f
C3372 iref.n32 vss 0.170249f
C3373 iref.n33 vss 0.103482f
C3374 iref.t144 vss 0.158044f
C3375 iref.t195 vss 0.158044f
C3376 iref.n34 vss 0.170249f
C3377 iref.n35 vss 0.103482f
C3378 iref.t201 vss 0.158044f
C3379 iref.t74 vss 0.158044f
C3380 iref.n36 vss 0.170249f
C3381 iref.n37 vss 0.103482f
C3382 iref.t78 vss 0.158044f
C3383 iref.t134 vss 0.158044f
C3384 iref.n38 vss 0.170249f
C3385 iref.n39 vss 0.103482f
C3386 iref.t141 vss 0.158044f
C3387 iref.t193 vss 0.158044f
C3388 iref.n40 vss 0.170249f
C3389 iref.n41 vss 0.103482f
C3390 iref.t63 vss 0.158044f
C3391 iref.t121 vss 0.158044f
C3392 iref.n42 vss 0.170249f
C3393 iref.n43 vss 0.103482f
C3394 iref.t171 vss 0.158044f
C3395 iref.t40 vss 0.158044f
C3396 iref.n44 vss 0.170249f
C3397 iref.n45 vss 0.103482f
C3398 iref.t47 vss 0.158044f
C3399 iref.t96 vss 0.158044f
C3400 iref.n46 vss 0.170249f
C3401 iref.n47 vss 0.103482f
C3402 iref.t103 vss 0.158044f
C3403 iref.t160 vss 0.158044f
C3404 iref.n48 vss 0.170249f
C3405 iref.n49 vss 0.103482f
C3406 iref.t167 vss 0.158044f
C3407 iref.t39 vss 0.158044f
C3408 iref.n50 vss 0.170249f
C3409 iref.n51 vss 0.103482f
C3410 iref.t208 vss 0.158044f
C3411 iref.t86 vss 0.158044f
C3412 iref.n52 vss 0.170249f
C3413 iref.n53 vss 0.103482f
C3414 iref.t138 vss 0.158044f
C3415 iref.t188 vss 0.158044f
C3416 iref.n54 vss 0.170249f
C3417 iref.n55 vss 0.617821f
C3418 iref.t70 vss 0.158044f
C3419 iref.t127 vss 0.158044f
C3420 iref.n56 vss 0.170249f
C3421 iref.n57 vss 0.617821f
C3422 iref.t181 vss 0.158044f
C3423 iref.t49 vss 0.158044f
C3424 iref.n58 vss 0.170249f
C3425 iref.n59 vss 0.103482f
C3426 iref.t57 vss 0.158044f
C3427 iref.t107 vss 0.158044f
C3428 iref.n60 vss 0.170249f
C3429 iref.n61 vss 0.103482f
C3430 iref.t116 vss 0.158044f
C3431 iref.t170 vss 0.158044f
C3432 iref.n62 vss 0.170249f
C3433 iref.n63 vss 0.103482f
C3434 iref.t179 vss 0.158044f
C3435 iref.t46 vss 0.158044f
C3436 iref.n64 vss 0.170249f
C3437 iref.n65 vss 0.103482f
C3438 iref.t33 vss 0.158044f
C3439 iref.t89 vss 0.158044f
C3440 iref.n66 vss 0.170249f
C3441 iref.n67 vss 0.103482f
C3442 iref.t151 vss 0.158044f
C3443 iref.t199 vss 0.158044f
C3444 iref.n68 vss 0.170249f
C3445 iref.n69 vss 0.103482f
C3446 iref.t205 vss 0.158044f
C3447 iref.t76 vss 0.158044f
C3448 iref.n70 vss 0.170249f
C3449 iref.n71 vss 0.103482f
C3450 iref.t81 vss 0.158044f
C3451 iref.t137 vss 0.158044f
C3452 iref.n72 vss 0.170249f
C3453 iref.n73 vss 0.103482f
C3454 iref.t146 vss 0.158044f
C3455 iref.t196 vss 0.158044f
C3456 iref.n74 vss 0.170249f
C3457 iref.n75 vss 0.103482f
C3458 iref.t68 vss 0.158044f
C3459 iref.t124 vss 0.158044f
C3460 iref.n76 vss 0.170249f
C3461 iref.n77 vss 0.103482f
C3462 iref.t128 vss 0.158044f
C3463 iref.t183 vss 0.158044f
C3464 iref.n78 vss 0.170249f
C3465 iref.n79 vss 0.103482f
C3466 iref.t53 vss 0.158044f
C3467 iref.t101 vss 0.158044f
C3468 iref.n80 vss 0.170249f
C3469 iref.n81 vss 0.103482f
C3470 iref.t48 vss 0.158044f
C3471 iref.t97 vss 0.158044f
C3472 iref.n82 vss 0.170249f
C3473 iref.n83 vss 0.103482f
C3474 iref.t105 vss 0.158044f
C3475 iref.t162 vss 0.158044f
C3476 iref.n84 vss 0.170249f
C3477 iref.n85 vss 0.103482f
C3478 iref.t30 vss 0.158044f
C3479 iref.t88 vss 0.158044f
C3480 iref.n86 vss 0.170249f
C3481 iref.n87 vss 0.103482f
C3482 iref.t91 vss 0.158044f
C3483 iref.t154 vss 0.158044f
C3484 iref.n88 vss 0.170249f
C3485 iref.n89 vss 0.103482f
C3486 iref.t200 vss 0.158044f
C3487 iref.t73 vss 0.158044f
C3488 iref.n90 vss 0.170249f
C3489 iref.n91 vss 0.103482f
C3490 iref.t77 vss 0.158044f
C3491 iref.t133 vss 0.158044f
C3492 iref.n92 vss 0.170249f
C3493 iref.n93 vss 0.103482f
C3494 iref.t140 vss 0.158044f
C3495 iref.t190 vss 0.158044f
C3496 iref.n94 vss 0.170249f
C3497 iref.n95 vss 0.103482f
C3498 iref.t62 vss 0.158044f
C3499 iref.t120 vss 0.158044f
C3500 iref.n96 vss 0.170249f
C3501 iref.n97 vss 0.103482f
C3502 iref.t125 vss 0.158044f
C3503 iref.t182 vss 0.158044f
C3504 iref.n98 vss 0.170249f
C3505 iref.n99 vss 0.103482f
C3506 iref.t123 vss 0.158044f
C3507 iref.t180 vss 0.158044f
C3508 iref.n100 vss 0.170249f
C3509 iref.n101 vss 0.103482f
C3510 iref.t44 vss 0.158044f
C3511 iref.t94 vss 0.158044f
C3512 iref.n102 vss 0.170249f
C3513 iref.n103 vss 0.103482f
C3514 iref.t100 vss 0.158044f
C3515 iref.t158 vss 0.158044f
C3516 iref.n104 vss 0.170249f
C3517 iref.n105 vss 0.617821f
C3518 iref.t64 vss 0.158044f
C3519 iref.t122 vss 0.158044f
C3520 iref.n106 vss 0.170249f
C3521 iref.n107 vss 0.617821f
C3522 iref.t174 vss 0.158044f
C3523 iref.t42 vss 0.158044f
C3524 iref.n108 vss 0.170249f
C3525 iref.n109 vss 0.103482f
C3526 iref.t50 vss 0.158044f
C3527 iref.t99 vss 0.158044f
C3528 iref.n110 vss 0.170249f
C3529 iref.n111 vss 0.103482f
C3530 iref.t106 vss 0.158044f
C3531 iref.t164 vss 0.158044f
C3532 iref.n112 vss 0.170249f
C3533 iref.n113 vss 0.103482f
C3534 iref.t104 vss 0.158044f
C3535 iref.t161 vss 0.158044f
C3536 iref.n114 vss 0.170249f
C3537 iref.n115 vss 0.103482f
C3538 iref.t209 vss 0.158044f
C3539 iref.t87 vss 0.158044f
C3540 iref.n116 vss 0.170249f
C3541 iref.n117 vss 0.103482f
C3542 iref.t142 vss 0.158044f
C3543 iref.t192 vss 0.158044f
C3544 iref.n118 vss 0.170249f
C3545 iref.n119 vss 0.103482f
C3546 iref.t198 vss 0.158044f
C3547 iref.t71 vss 0.158044f
C3548 iref.n120 vss 0.170249f
C3549 iref.n121 vss 0.103482f
C3550 iref.t75 vss 0.158044f
C3551 iref.t131 vss 0.158044f
C3552 iref.n122 vss 0.170249f
C3553 iref.n123 vss 0.103482f
C3554 iref.t136 vss 0.158044f
C3555 iref.t189 vss 0.158044f
C3556 iref.n124 vss 0.170249f
C3557 iref.n125 vss 0.103482f
C3558 iref.t60 vss 0.158044f
C3559 iref.t118 vss 0.158044f
C3560 iref.n126 vss 0.170249f
C3561 iref.n127 vss 0.103482f
C3562 iref.t168 vss 0.158044f
C3563 iref.t38 vss 0.158044f
C3564 iref.n128 vss 0.170249f
C3565 iref.n129 vss 0.103482f
C3566 iref.t165 vss 0.158044f
C3567 iref.t34 vss 0.158044f
C3568 iref.n130 vss 0.170249f
C3569 iref.n131 vss 0.103482f
C3570 iref.t41 vss 0.158044f
C3571 iref.t93 vss 0.158044f
C3572 iref.n132 vss 0.170249f
C3573 iref.n133 vss 0.103482f
C3574 iref.t98 vss 0.158044f
C3575 iref.t157 vss 0.158044f
C3576 iref.n134 vss 0.170249f
C3577 iref.n135 vss 0.103482f
C3578 iref.t163 vss 0.158044f
C3579 iref.t32 vss 0.158044f
C3580 iref.n136 vss 0.170249f
C3581 iref.n137 vss 0.103482f
C3582 iref.t135 vss 0.158044f
C3583 iref.t187 vss 0.158044f
C3584 iref.n138 vss 0.170249f
C3585 iref.n139 vss 0.103482f
C3586 iref.t194 vss 0.158044f
C3587 iref.t69 vss 0.158044f
C3588 iref.n140 vss 0.170249f
C3589 iref.n141 vss 0.103482f
C3590 iref.t72 vss 0.158044f
C3591 iref.t130 vss 0.158044f
C3592 iref.n142 vss 0.170249f
C3593 iref.n143 vss 0.103482f
C3594 iref.t132 vss 0.158044f
C3595 iref.t184 vss 0.158044f
C3596 iref.n144 vss 0.170249f
C3597 iref.n145 vss 0.103482f
C3598 iref.t191 vss 0.158044f
C3599 iref.t66 vss 0.158044f
C3600 iref.n146 vss 0.170249f
C3601 iref.n147 vss 0.103482f
C3602 iref.t59 vss 0.158044f
C3603 iref.t110 vss 0.158044f
C3604 iref.n148 vss 0.170249f
C3605 iref.n149 vss 0.103482f
C3606 iref.t159 vss 0.158044f
C3607 iref.t31 vss 0.158044f
C3608 iref.n150 vss 0.170249f
C3609 iref.n151 vss 0.103482f
C3610 iref.t37 vss 0.158044f
C3611 iref.t92 vss 0.158044f
C3612 iref.n152 vss 0.170249f
C3613 iref.n153 vss 0.103482f
C3614 iref.t95 vss 0.158044f
C3615 iref.t155 vss 0.158044f
C3616 iref.n154 vss 0.170249f
C3617 iref.n155 vss 0.947124f
C3618 iref.t147 vss 0.158929f
C3619 iref.n156 vss 1.03671f
C3620 iref.t65 vss 0.158929f
C3621 iref.n157 vss 0.193065f
C3622 iref.t126 vss 0.158929f
C3623 iref.n158 vss 0.193065f
C3624 iref.t52 vss 0.158929f
C3625 iref.n159 vss 0.193065f
C3626 iref.t109 vss 0.158929f
C3627 iref.n160 vss 0.193065f
C3628 iref.t150 vss 0.158929f
C3629 iref.n161 vss 0.193065f
C3630 iref.t67 vss 0.158929f
C3631 iref.n162 vss 0.193065f
C3632 iref.t129 vss 0.158929f
C3633 iref.n163 vss 0.193065f
C3634 iref.t56 vss 0.158929f
C3635 iref.n164 vss 0.193065f
C3636 iref.t113 vss 0.158929f
C3637 iref.n165 vss 0.193065f
C3638 iref.t176 vss 0.158929f
C3639 iref.n166 vss 0.193065f
C3640 iref.t51 vss 0.158929f
C3641 iref.n167 vss 0.193065f
C3642 iref.t156 vss 0.158929f
C3643 iref.n168 vss 0.193065f
C3644 iref.t204 vss 0.202595f
C3645 iref.n169 vss 0.193065f
C3646 iref.t80 vss 0.158929f
C3647 iref.n170 vss 0.293039f
C3648 iref.t119 vss 0.158929f
C3649 iref.n171 vss 0.293039f
C3650 iref.t36 vss 0.158929f
C3651 iref.n172 vss 0.193065f
C3652 iref.t153 vss 0.158929f
C3653 iref.n173 vss 0.193065f
C3654 iref.t207 vss 0.158929f
C3655 iref.n174 vss 0.193065f
C3656 iref.t85 vss 0.158929f
C3657 iref.n175 vss 0.193065f
C3658 iref.t83 vss 0.158929f
C3659 iref.n176 vss 0.193065f
C3660 iref.t186 vss 0.158929f
C3661 iref.n177 vss 0.193065f
C3662 iref.t115 vss 0.158929f
C3663 iref.n178 vss 0.193065f
C3664 iref.t178 vss 0.158929f
C3665 iref.n179 vss 0.193065f
C3666 iref.t55 vss 0.158929f
C3667 iref.n180 vss 0.193065f
C3668 iref.t112 vss 0.158929f
C3669 iref.n181 vss 0.193065f
C3670 iref.t175 vss 0.158929f
C3671 iref.n182 vss 0.193065f
C3672 iref.t149 vss 0.158929f
C3673 iref.n183 vss 0.193065f
C3674 iref.t145 vss 0.202595f
C3675 iref.n184 vss 0.193065f
C3676 iref.t203 vss 0.158929f
C3677 iref.n185 vss 0.267166f
C3678 iref.n186 vss 0.623214f
C3679 iref.t28 vss 0.158929f
C3680 iref.n187 vss 0.167191f
C3681 iref.t2 vss 0.158929f
C3682 iref.n188 vss 0.167191f
C3683 iref.n189 vss 0.507523f
C3684 iref.t12 vss 0.158929f
C3685 iref.n190 vss 0.167191f
C3686 iref.t22 vss 0.158929f
C3687 iref.n191 vss 0.167191f
C3688 iref.n192 vss 0.507523f
C3689 iref.t10 vss 0.158929f
C3690 iref.n193 vss 0.167191f
C3691 iref.t26 vss 0.158929f
C3692 iref.n194 vss 0.167191f
C3693 iref.n195 vss 0.507523f
C3694 iref.t20 vss 0.158929f
C3695 iref.n196 vss 0.167191f
C3696 iref.t6 vss 0.158929f
C3697 iref.n197 vss 0.167191f
C3698 iref.n198 vss 0.507523f
C3699 iref.t4 vss 0.158929f
C3700 iref.n199 vss 0.167191f
C3701 iref.t16 vss 0.158929f
C3702 iref.n200 vss 0.167191f
C3703 iref.n201 vss 0.507523f
C3704 iref.t8 vss 0.158929f
C3705 iref.n202 vss 0.167191f
C3706 iref.t0 vss 0.158929f
C3707 iref.n203 vss 0.167191f
C3708 iref.n204 vss 0.507523f
C3709 iref.t18 vss 0.158929f
C3710 iref.n205 vss 0.167191f
C3711 iref.t14 vss 0.202595f
C3712 iref.n206 vss 0.167191f
C3713 iref.n207 vss 0.507523f
C3714 iref.t24 vss 0.158929f
C3715 iref.n208 vss 1.35066f
C3716 vin_p.t182 vss 0.127716f
C3717 vin_p.t181 vss 0.127716f
C3718 vin_p.n0 vss 0.125934f
C3719 vin_p.t128 vss 0.127716f
C3720 vin_p.t127 vss 0.127716f
C3721 vin_p.n1 vss 0.125751f
C3722 vin_p.n2 vss 0.301849f
C3723 vin_p.t120 vss 0.127716f
C3724 vin_p.t119 vss 0.127716f
C3725 vin_p.n3 vss 0.125751f
C3726 vin_p.n4 vss 0.162518f
C3727 vin_p.t56 vss 0.127716f
C3728 vin_p.t55 vss 0.127716f
C3729 vin_p.n5 vss 0.125751f
C3730 vin_p.n6 vss 0.162518f
C3731 vin_p.t46 vss 0.127716f
C3732 vin_p.t45 vss 0.127716f
C3733 vin_p.n7 vss 0.125751f
C3734 vin_p.n8 vss 0.162518f
C3735 vin_p.t40 vss 0.127716f
C3736 vin_p.t39 vss 0.127716f
C3737 vin_p.n9 vss 0.125751f
C3738 vin_p.n10 vss 0.162518f
C3739 vin_p.t172 vss 0.127716f
C3740 vin_p.t170 vss 0.127716f
C3741 vin_p.n11 vss 0.125751f
C3742 vin_p.n12 vss 0.162518f
C3743 vin_p.t164 vss 0.127716f
C3744 vin_p.t163 vss 0.127716f
C3745 vin_p.n13 vss 0.125751f
C3746 vin_p.n14 vss 0.162518f
C3747 vin_p.t98 vss 0.127716f
C3748 vin_p.t97 vss 0.127716f
C3749 vin_p.n15 vss 0.125751f
C3750 vin_p.n16 vss 0.162518f
C3751 vin_p.t94 vss 0.127716f
C3752 vin_p.t93 vss 0.127716f
C3753 vin_p.n17 vss 0.125751f
C3754 vin_p.n18 vss 0.162518f
C3755 vin_p.t91 vss 0.127716f
C3756 vin_p.t89 vss 0.127716f
C3757 vin_p.n19 vss 0.125751f
C3758 vin_p.n20 vss 0.162518f
C3759 vin_p.t32 vss 0.127716f
C3760 vin_p.t30 vss 0.127716f
C3761 vin_p.n21 vss 0.125751f
C3762 vin_p.n22 vss 0.162518f
C3763 vin_p.t26 vss 0.127716f
C3764 vin_p.t25 vss 0.127716f
C3765 vin_p.n23 vss 0.125751f
C3766 vin_p.n24 vss 0.162518f
C3767 vin_p.t24 vss 0.127716f
C3768 vin_p.t23 vss 0.127716f
C3769 vin_p.n25 vss 0.125751f
C3770 vin_p.n26 vss 0.162518f
C3771 vin_p.t177 vss 0.127716f
C3772 vin_p.t174 vss 0.127716f
C3773 vin_p.n27 vss 0.125751f
C3774 vin_p.n28 vss 0.162518f
C3775 vin_p.t167 vss 0.127716f
C3776 vin_p.t166 vss 0.127716f
C3777 vin_p.n29 vss 0.125751f
C3778 vin_p.n30 vss 0.162518f
C3779 vin_p.t116 vss 0.127716f
C3780 vin_p.t115 vss 0.127716f
C3781 vin_p.n31 vss 0.125751f
C3782 vin_p.n32 vss 0.162518f
C3783 vin_p.t109 vss 0.127716f
C3784 vin_p.t107 vss 0.127716f
C3785 vin_p.n33 vss 0.125751f
C3786 vin_p.n34 vss 0.162518f
C3787 vin_p.t103 vss 0.127716f
C3788 vin_p.t101 vss 0.127716f
C3789 vin_p.n35 vss 0.125751f
C3790 vin_p.n36 vss 0.162518f
C3791 vin_p.t35 vss 0.127716f
C3792 vin_p.t33 vss 0.127716f
C3793 vin_p.n37 vss 0.125751f
C3794 vin_p.n38 vss 0.162518f
C3795 vin_p.t28 vss 0.127716f
C3796 vin_p.t27 vss 0.127716f
C3797 vin_p.n39 vss 0.125751f
C3798 vin_p.n40 vss 0.162518f
C3799 vin_p.t180 vss 0.127716f
C3800 vin_p.t179 vss 0.127716f
C3801 vin_p.n41 vss 0.125751f
C3802 vin_p.n42 vss 0.162518f
C3803 vin_p.t171 vss 0.127716f
C3804 vin_p.t169 vss 0.127716f
C3805 vin_p.n43 vss 0.125751f
C3806 vin_p.n44 vss 0.162518f
C3807 vin_p.t191 vss 0.127716f
C3808 vin_p.t188 vss 0.127716f
C3809 vin_p.n45 vss 0.125751f
C3810 vin_p.n46 vss 0.162518f
C3811 vin_p.t185 vss 0.127716f
C3812 vin_p.t183 vss 0.127716f
C3813 vin_p.n47 vss 0.125751f
C3814 vin_p.n48 vss 0.162518f
C3815 vin_p.t113 vss 0.127716f
C3816 vin_p.t112 vss 0.127716f
C3817 vin_p.n49 vss 0.125751f
C3818 vin_p.n50 vss 0.162518f
C3819 vin_p.t66 vss 0.127716f
C3820 vin_p.t65 vss 0.127716f
C3821 vin_p.n51 vss 0.125751f
C3822 vin_p.n52 vss 0.162518f
C3823 vin_p.t63 vss 0.127716f
C3824 vin_p.t62 vss 0.127716f
C3825 vin_p.n53 vss 0.125751f
C3826 vin_p.n54 vss 0.162518f
C3827 vin_p.t52 vss 0.127716f
C3828 vin_p.t49 vss 0.127716f
C3829 vin_p.n55 vss 0.125751f
C3830 vin_p.n56 vss 0.162518f
C3831 vin_p.t43 vss 0.127716f
C3832 vin_p.t41 vss 0.127716f
C3833 vin_p.n57 vss 0.125751f
C3834 vin_p.n58 vss 0.162518f
C3835 vin_p.t176 vss 0.127716f
C3836 vin_p.t175 vss 0.127716f
C3837 vin_p.n59 vss 0.125751f
C3838 vin_p.n60 vss 0.162518f
C3839 vin_p.t146 vss 0.127716f
C3840 vin_p.t143 vss 0.127716f
C3841 vin_p.n61 vss 0.125751f
C3842 vin_p.n62 vss 0.162518f
C3843 vin_p.t141 vss 0.127716f
C3844 vin_p.t140 vss 0.127716f
C3845 vin_p.n63 vss 0.125751f
C3846 vin_p.n64 vss 0.162518f
C3847 vin_p.t137 vss 0.127716f
C3848 vin_p.t136 vss 0.127716f
C3849 vin_p.n65 vss 0.125751f
C3850 vin_p.n66 vss 0.162518f
C3851 vin_p.t131 vss 0.127716f
C3852 vin_p.t130 vss 0.127716f
C3853 vin_p.n67 vss 0.125751f
C3854 vin_p.n68 vss 0.162518f
C3855 vin_p.t123 vss 0.127716f
C3856 vin_p.t122 vss 0.127716f
C3857 vin_p.n69 vss 0.125751f
C3858 vin_p.n70 vss 0.162518f
C3859 vin_p.t4 vss 0.127716f
C3860 vin_p.t2 vss 0.127716f
C3861 vin_p.n71 vss 0.125751f
C3862 vin_p.n72 vss 0.162518f
C3863 vin_p.t0 vss 0.127716f
C3864 vin_p.t199 vss 0.127716f
C3865 vin_p.n73 vss 0.125751f
C3866 vin_p.n74 vss 0.162518f
C3867 vin_p.t197 vss 0.127716f
C3868 vin_p.t196 vss 0.127716f
C3869 vin_p.n75 vss 0.125751f
C3870 vin_p.n76 vss 0.162518f
C3871 vin_p.t190 vss 0.127716f
C3872 vin_p.t189 vss 0.127716f
C3873 vin_p.n77 vss 0.125751f
C3874 vin_p.n78 vss 0.162518f
C3875 vin_p.t11 vss 0.127716f
C3876 vin_p.t10 vss 0.127716f
C3877 vin_p.n79 vss 0.125751f
C3878 vin_p.n80 vss 0.162518f
C3879 vin_p.t152 vss 0.127716f
C3880 vin_p.t151 vss 0.127716f
C3881 vin_p.n81 vss 0.125751f
C3882 vin_p.n82 vss 0.162518f
C3883 vin_p.t87 vss 0.127716f
C3884 vin_p.t86 vss 0.127716f
C3885 vin_p.n83 vss 0.125751f
C3886 vin_p.n84 vss 0.162518f
C3887 vin_p.t83 vss 0.127716f
C3888 vin_p.t82 vss 0.127716f
C3889 vin_p.n85 vss 0.125751f
C3890 vin_p.n86 vss 0.162518f
C3891 vin_p.t79 vss 0.127716f
C3892 vin_p.t78 vss 0.127716f
C3893 vin_p.n87 vss 0.125751f
C3894 vin_p.n88 vss 0.162518f
C3895 vin_p.t74 vss 0.127716f
C3896 vin_p.t73 vss 0.127716f
C3897 vin_p.n89 vss 0.125751f
C3898 vin_p.n90 vss 0.162518f
C3899 vin_p.t16 vss 0.127716f
C3900 vin_p.t15 vss 0.127716f
C3901 vin_p.n91 vss 0.125751f
C3902 vin_p.n92 vss 0.162518f
C3903 vin_p.t145 vss 0.127716f
C3904 vin_p.t144 vss 0.127716f
C3905 vin_p.n93 vss 0.125751f
C3906 vin_p.n94 vss 0.162518f
C3907 vin_p.t159 vss 0.127716f
C3908 vin_p.t158 vss 0.127716f
C3909 vin_p.n95 vss 0.125751f
C3910 vin_p.n96 vss 0.162518f
C3911 vin_p.t155 vss 0.127716f
C3912 vin_p.t154 vss 0.127716f
C3913 vin_p.n97 vss 0.125751f
C3914 vin_p.n98 vss 0.725129f
C3915 vin_p.t68 vss 0.127716f
C3916 vin_p.t67 vss 0.127716f
C3917 vin_p.n99 vss 0.125934f
C3918 vin_p.t8 vss 0.127716f
C3919 vin_p.t7 vss 0.127716f
C3920 vin_p.n100 vss 0.125751f
C3921 vin_p.n101 vss 0.301849f
C3922 vin_p.t3 vss 0.127716f
C3923 vin_p.t1 vss 0.127716f
C3924 vin_p.n102 vss 0.125751f
C3925 vin_p.n103 vss 0.162518f
C3926 vin_p.t134 vss 0.127716f
C3927 vin_p.t133 vss 0.127716f
C3928 vin_p.n104 vss 0.125751f
C3929 vin_p.n105 vss 0.162518f
C3930 vin_p.t126 vss 0.127716f
C3931 vin_p.t125 vss 0.127716f
C3932 vin_p.n106 vss 0.125751f
C3933 vin_p.n107 vss 0.162518f
C3934 vin_p.t118 vss 0.127716f
C3935 vin_p.t117 vss 0.127716f
C3936 vin_p.n108 vss 0.125751f
C3937 vin_p.n109 vss 0.162518f
C3938 vin_p.t53 vss 0.127716f
C3939 vin_p.t50 vss 0.127716f
C3940 vin_p.n110 vss 0.125751f
C3941 vin_p.n111 vss 0.162518f
C3942 vin_p.t44 vss 0.127716f
C3943 vin_p.t42 vss 0.127716f
C3944 vin_p.n112 vss 0.125751f
C3945 vin_p.n113 vss 0.162518f
C3946 vin_p.t178 vss 0.127716f
C3947 vin_p.t173 vss 0.127716f
C3948 vin_p.n114 vss 0.125751f
C3949 vin_p.n115 vss 0.162518f
C3950 vin_p.t168 vss 0.127716f
C3951 vin_p.t165 vss 0.127716f
C3952 vin_p.n116 vss 0.125751f
C3953 vin_p.n117 vss 0.162518f
C3954 vin_p.t162 vss 0.127716f
C3955 vin_p.t161 vss 0.127716f
C3956 vin_p.n118 vss 0.125751f
C3957 vin_p.n119 vss 0.162518f
C3958 vin_p.t110 vss 0.127716f
C3959 vin_p.t108 vss 0.127716f
C3960 vin_p.n120 vss 0.125751f
C3961 vin_p.n121 vss 0.162518f
C3962 vin_p.t104 vss 0.127716f
C3963 vin_p.t102 vss 0.127716f
C3964 vin_p.n122 vss 0.125751f
C3965 vin_p.n123 vss 0.162518f
C3966 vin_p.t100 vss 0.127716f
C3967 vin_p.t99 vss 0.127716f
C3968 vin_p.n124 vss 0.125751f
C3969 vin_p.n125 vss 0.162518f
C3970 vin_p.t59 vss 0.127716f
C3971 vin_p.t57 vss 0.127716f
C3972 vin_p.n126 vss 0.125751f
C3973 vin_p.n127 vss 0.162518f
C3974 vin_p.t48 vss 0.127716f
C3975 vin_p.t47 vss 0.127716f
C3976 vin_p.n128 vss 0.125751f
C3977 vin_p.n129 vss 0.162518f
C3978 vin_p.t198 vss 0.127716f
C3979 vin_p.t195 vss 0.127716f
C3980 vin_p.n130 vss 0.125751f
C3981 vin_p.n131 vss 0.162518f
C3982 vin_p.t192 vss 0.127716f
C3983 vin_p.t187 vss 0.127716f
C3984 vin_p.n132 vss 0.125751f
C3985 vin_p.n133 vss 0.162518f
C3986 vin_p.t186 vss 0.127716f
C3987 vin_p.t184 vss 0.127716f
C3988 vin_p.n134 vss 0.125751f
C3989 vin_p.n135 vss 0.162518f
C3990 vin_p.t114 vss 0.127716f
C3991 vin_p.t111 vss 0.127716f
C3992 vin_p.n136 vss 0.125751f
C3993 vin_p.n137 vss 0.162518f
C3994 vin_p.t106 vss 0.127716f
C3995 vin_p.t105 vss 0.127716f
C3996 vin_p.n138 vss 0.125751f
C3997 vin_p.n139 vss 0.162518f
C3998 vin_p.t64 vss 0.127716f
C3999 vin_p.t61 vss 0.127716f
C4000 vin_p.n140 vss 0.125751f
C4001 vin_p.n141 vss 0.162518f
C4002 vin_p.t54 vss 0.127716f
C4003 vin_p.t51 vss 0.127716f
C4004 vin_p.n142 vss 0.125751f
C4005 vin_p.n143 vss 0.162518f
C4006 vin_p.t75 vss 0.127716f
C4007 vin_p.t71 vss 0.127716f
C4008 vin_p.n144 vss 0.125751f
C4009 vin_p.n145 vss 0.162518f
C4010 vin_p.t70 vss 0.127716f
C4011 vin_p.t69 vss 0.127716f
C4012 vin_p.n146 vss 0.125751f
C4013 vin_p.n147 vss 0.162518f
C4014 vin_p.t194 vss 0.127716f
C4015 vin_p.t193 vss 0.127716f
C4016 vin_p.n148 vss 0.125751f
C4017 vin_p.n149 vss 0.162518f
C4018 vin_p.t142 vss 0.127716f
C4019 vin_p.t139 vss 0.127716f
C4020 vin_p.n150 vss 0.125751f
C4021 vin_p.n151 vss 0.162518f
C4022 vin_p.t138 vss 0.127716f
C4023 vin_p.t135 vss 0.127716f
C4024 vin_p.n152 vss 0.125751f
C4025 vin_p.n153 vss 0.162518f
C4026 vin_p.t132 vss 0.127716f
C4027 vin_p.t129 vss 0.127716f
C4028 vin_p.n154 vss 0.125751f
C4029 vin_p.n155 vss 0.162518f
C4030 vin_p.t124 vss 0.127716f
C4031 vin_p.t121 vss 0.127716f
C4032 vin_p.n156 vss 0.125751f
C4033 vin_p.n157 vss 0.162518f
C4034 vin_p.t60 vss 0.127716f
C4035 vin_p.t58 vss 0.127716f
C4036 vin_p.n158 vss 0.125751f
C4037 vin_p.n159 vss 0.162518f
C4038 vin_p.t21 vss 0.127716f
C4039 vin_p.t19 vss 0.127716f
C4040 vin_p.n160 vss 0.125751f
C4041 vin_p.n161 vss 0.162518f
C4042 vin_p.t18 vss 0.127716f
C4043 vin_p.t17 vss 0.127716f
C4044 vin_p.n162 vss 0.125751f
C4045 vin_p.n163 vss 0.162518f
C4046 vin_p.t14 vss 0.127716f
C4047 vin_p.t13 vss 0.127716f
C4048 vin_p.n164 vss 0.125751f
C4049 vin_p.n165 vss 0.162518f
C4050 vin_p.t12 vss 0.127716f
C4051 vin_p.t9 vss 0.127716f
C4052 vin_p.n166 vss 0.125751f
C4053 vin_p.n167 vss 0.162518f
C4054 vin_p.t6 vss 0.127716f
C4055 vin_p.t5 vss 0.127716f
C4056 vin_p.n168 vss 0.125751f
C4057 vin_p.n169 vss 0.162518f
C4058 vin_p.t88 vss 0.127716f
C4059 vin_p.t85 vss 0.127716f
C4060 vin_p.n170 vss 0.125751f
C4061 vin_p.n171 vss 0.162518f
C4062 vin_p.t84 vss 0.127716f
C4063 vin_p.t81 vss 0.127716f
C4064 vin_p.n172 vss 0.125751f
C4065 vin_p.n173 vss 0.162518f
C4066 vin_p.t80 vss 0.127716f
C4067 vin_p.t77 vss 0.127716f
C4068 vin_p.n174 vss 0.125751f
C4069 vin_p.n175 vss 0.162518f
C4070 vin_p.t76 vss 0.127716f
C4071 vin_p.t72 vss 0.127716f
C4072 vin_p.n176 vss 0.125751f
C4073 vin_p.n177 vss 0.162518f
C4074 vin_p.t92 vss 0.127716f
C4075 vin_p.t90 vss 0.127716f
C4076 vin_p.n178 vss 0.125751f
C4077 vin_p.n179 vss 0.162518f
C4078 vin_p.t31 vss 0.127716f
C4079 vin_p.t29 vss 0.127716f
C4080 vin_p.n180 vss 0.125751f
C4081 vin_p.n181 vss 0.162518f
C4082 vin_p.t160 vss 0.127716f
C4083 vin_p.t157 vss 0.127716f
C4084 vin_p.n182 vss 0.125751f
C4085 vin_p.n183 vss 0.162518f
C4086 vin_p.t156 vss 0.127716f
C4087 vin_p.t153 vss 0.127716f
C4088 vin_p.n184 vss 0.125751f
C4089 vin_p.n185 vss 0.162518f
C4090 vin_p.t150 vss 0.127716f
C4091 vin_p.t149 vss 0.127716f
C4092 vin_p.n186 vss 0.125751f
C4093 vin_p.n187 vss 0.162518f
C4094 vin_p.t148 vss 0.127716f
C4095 vin_p.t147 vss 0.127716f
C4096 vin_p.n188 vss 0.125751f
C4097 vin_p.n189 vss 0.162518f
C4098 vin_p.t96 vss 0.127716f
C4099 vin_p.t95 vss 0.127716f
C4100 vin_p.n190 vss 0.125751f
C4101 vin_p.n191 vss 0.162518f
C4102 vin_p.t22 vss 0.127716f
C4103 vin_p.t20 vss 0.127716f
C4104 vin_p.n192 vss 0.125751f
C4105 vin_p.n193 vss 0.162482f
C4106 vin_p.t38 vss 0.127716f
C4107 vin_p.t37 vss 0.127716f
C4108 vin_p.n194 vss 0.125751f
C4109 vin_p.n195 vss 0.162935f
C4110 vin_p.t36 vss 0.127716f
C4111 vin_p.t34 vss 0.127716f
C4112 vin_p.n196 vss 0.125751f
C4113 vin_p.n197 vss 0.724796f
C4114 vin_p.n198 vss 1.97419f
C4115 w_4660_n6791.n0 vss 0.697187f
C4116 w_4660_n6791.n1 vss 0.075269f
C4117 w_4660_n6791.n2 vss 0.007326f
C4118 w_4660_n6791.n3 vss 0.078245f
C4119 w_4660_n6791.n4 vss 0.696682f
C4120 w_4660_n6791.n5 vss 0.064443f
C4121 w_4660_n6791.n6 vss 0.065338f
C4122 w_4660_n6791.n7 vss 0.008764f
C4123 w_4660_n6791.n8 vss 0.065338f
C4124 w_4660_n6791.n9 vss 0.008764f
C4125 w_4660_n6791.n10 vss 0.065338f
C4126 w_4660_n6791.n11 vss 0.008764f
C4127 w_4660_n6791.n12 vss 0.065338f
C4128 w_4660_n6791.n13 vss 0.008764f
C4129 w_4660_n6791.n14 vss 0.065338f
C4130 w_4660_n6791.n15 vss 0.008764f
C4131 w_4660_n6791.n16 vss 0.065338f
C4132 w_4660_n6791.n17 vss 0.008764f
C4133 w_4660_n6791.n18 vss 0.065338f
C4134 w_4660_n6791.n19 vss 0.008764f
C4135 w_4660_n6791.n20 vss 0.065338f
C4136 w_4660_n6791.n21 vss 0.063548f
C4137 w_4660_n6791.n22 vss 0.065338f
C4138 w_4660_n6791.n23 vss 0.008764f
C4139 w_4660_n6791.n24 vss 0.065338f
C4140 w_4660_n6791.n25 vss 0.063548f
C4141 w_4660_n6791.n26 vss 0.065338f
C4142 w_4660_n6791.n27 vss 0.008764f
C4143 w_4660_n6791.n28 vss 0.065338f
C4144 w_4660_n6791.n29 vss 0.063548f
C4145 w_4660_n6791.n30 vss 0.065338f
C4146 w_4660_n6791.n31 vss 0.065338f
C4147 w_4660_n6791.n32 vss 0.063548f
C4148 w_4660_n6791.n33 vss 0.065338f
C4149 w_4660_n6791.n34 vss 0.081778f
C4150 w_4660_n6791.n35 vss 0.707001f
C4151 w_4660_n6791.n36 vss 0.032221f
C4152 w_4660_n6791.n37 vss 0.421054f
C4153 w_4660_n6791.n38 vss 0.693654f
C4154 w_4660_n6791.n40 vss 0.313182f
C4155 w_4660_n6791.t266 vss 0.031147f
C4156 w_4660_n6791.n41 vss 0.073197f
C4157 w_4660_n6791.n42 vss 0.032221f
C4158 w_4660_n6791.t346 vss 0.120265f
C4159 w_4660_n6791.n43 vss 0.508901f
C4160 w_4660_n6791.n44 vss 0.092379f
C4161 w_4660_n6791.t274 vss 0.031147f
C4162 w_4660_n6791.t248 vss 0.031147f
C4163 w_4660_n6791.n45 vss 0.069153f
C4164 w_4660_n6791.n46 vss 0.087331f
C4165 w_4660_n6791.n47 vss 0.059968f
C4166 w_4660_n6791.n48 vss 0.008764f
C4167 w_4660_n6791.n49 vss 0.064443f
C4168 w_4660_n6791.n50 vss 0.008764f
C4169 w_4660_n6791.n51 vss 0.008764f
C4170 w_4660_n6791.n52 vss 0.008764f
C4171 w_4660_n6791.n53 vss 0.008764f
C4172 w_4660_n6791.n54 vss 0.008764f
C4173 w_4660_n6791.n55 vss 0.036697f
C4174 w_4660_n6791.n56 vss 0.008764f
C4175 w_4660_n6791.n57 vss 0.008764f
C4176 w_4660_n6791.n58 vss 0.008764f
C4177 w_4660_n6791.n59 vss 0.008764f
C4178 w_4660_n6791.n60 vss 0.064443f
C4179 w_4660_n6791.n61 vss 0.00773f
C4180 w_4660_n6791.n62 vss 0.008764f
C4181 w_4660_n6791.n63 vss 0.008764f
C4182 w_4660_n6791.n64 vss 0.028194f
C4183 w_4660_n6791.n65 vss 0.012964f
C4184 w_4660_n6791.n66 vss 0.060863f
C4185 w_4660_n6791.n67 vss 0.008764f
C4186 w_4660_n6791.n68 vss 0.043363f
C4187 w_4660_n6791.n69 vss 0.068999f
C4188 w_4660_n6791.n70 vss 0.008764f
C4189 w_4660_n6791.n71 vss 0.010661f
C4190 w_4660_n6791.n72 vss 0.009834f
C4191 w_4660_n6791.n73 vss 0.008374f
C4192 w_4660_n6791.n74 vss 0.061865f
C4193 w_4660_n6791.n75 vss 0.010661f
C4194 w_4660_n6791.n76 vss 0.008764f
C4195 w_4660_n6791.n77 vss 0.008764f
C4196 w_4660_n6791.n78 vss 0.051497f
C4197 w_4660_n6791.n79 vss 0.008764f
C4198 w_4660_n6791.n80 vss 0.008764f
C4199 w_4660_n6791.n81 vss 0.037132f
C4200 w_4660_n6791.n82 vss 0.008825f
C4201 w_4660_n6791.n83 vss 0.012355f
C4202 w_4660_n6791.n84 vss 0.009022f
C4203 w_4660_n6791.n85 vss 0.008764f
C4204 w_4660_n6791.n86 vss 0.008764f
C4205 w_4660_n6791.n87 vss 0.061865f
C4206 w_4660_n6791.n88 vss 0.008764f
C4207 w_4660_n6791.n89 vss 0.008764f
C4208 w_4660_n6791.n90 vss 0.008764f
C4209 w_4660_n6791.n91 vss 0.061865f
C4210 w_4660_n6791.n92 vss 0.009022f
C4211 w_4660_n6791.n93 vss 0.009022f
C4212 w_4660_n6791.n94 vss 0.008764f
C4213 w_4660_n6791.n95 vss 0.008764f
C4214 w_4660_n6791.n96 vss 0.061865f
C4215 w_4660_n6791.n97 vss 0.008764f
C4216 w_4660_n6791.n98 vss 0.008764f
C4217 w_4660_n6791.n99 vss 0.008764f
C4218 w_4660_n6791.n100 vss 0.061865f
C4219 w_4660_n6791.n101 vss 0.009022f
C4220 w_4660_n6791.n102 vss 0.008764f
C4221 w_4660_n6791.n103 vss 0.008764f
C4222 w_4660_n6791.n104 vss 0.061865f
C4223 w_4660_n6791.n105 vss 0.008764f
C4224 w_4660_n6791.n106 vss 0.008764f
C4225 w_4660_n6791.n107 vss 0.008764f
C4226 w_4660_n6791.n108 vss 0.061865f
C4227 w_4660_n6791.n109 vss 0.00595f
C4228 w_4660_n6791.n110 vss 0.479417f
C4229 w_4660_n6791.n111 vss 0.479417f
C4230 w_4660_n6791.t77 vss 4.35485f
C4231 w_4660_n6791.n112 vss 0.48173f
C4232 w_4660_n6791.n113 vss 0.48173f
C4233 w_4660_n6791.n114 vss 0.479417f
C4234 w_4660_n6791.n115 vss 0.479417f
C4235 w_4660_n6791.n116 vss 0.007329f
C4236 w_4660_n6791.n117 vss 0.009022f
C4237 w_4660_n6791.n118 vss 0.061865f
C4238 w_4660_n6791.n119 vss 0.008764f
C4239 w_4660_n6791.n120 vss 0.061865f
C4240 w_4660_n6791.n121 vss 0.008764f
C4241 w_4660_n6791.n122 vss 0.008764f
C4242 w_4660_n6791.n123 vss 0.008764f
C4243 w_4660_n6791.n124 vss 0.008764f
C4244 w_4660_n6791.n125 vss 0.061865f
C4245 w_4660_n6791.n126 vss 0.009022f
C4246 w_4660_n6791.n127 vss 0.008764f
C4247 w_4660_n6791.n128 vss 0.008764f
C4248 w_4660_n6791.n129 vss 0.061865f
C4249 w_4660_n6791.n130 vss 0.008764f
C4250 w_4660_n6791.n131 vss 0.008764f
C4251 w_4660_n6791.n132 vss 0.008764f
C4252 w_4660_n6791.n133 vss 0.061865f
C4253 w_4660_n6791.n134 vss 0.009022f
C4254 w_4660_n6791.n135 vss 0.008764f
C4255 w_4660_n6791.n136 vss 0.008764f
C4256 w_4660_n6791.n137 vss 0.061865f
C4257 w_4660_n6791.n138 vss 0.010849f
C4258 w_4660_n6791.n139 vss 0.008764f
C4259 w_4660_n6791.n140 vss 0.008764f
C4260 w_4660_n6791.n141 vss 0.042962f
C4261 w_4660_n6791.n142 vss 0.00773f
C4262 w_4660_n6791.n143 vss 0.069813f
C4263 w_4660_n6791.n144 vss 0.008825f
C4264 w_4660_n6791.n145 vss 0.005404f
C4265 w_4660_n6791.n146 vss 0.008764f
C4266 w_4660_n6791.n147 vss 0.045647f
C4267 w_4660_n6791.t434 vss 0.121336f
C4268 w_4660_n6791.t78 vss 0.120265f
C4269 w_4660_n6791.t111 vss 0.031147f
C4270 w_4660_n6791.t436 vss 0.031147f
C4271 w_4660_n6791.n148 vss 0.07032f
C4272 w_4660_n6791.t171 vss 0.031147f
C4273 w_4660_n6791.t151 vss 0.031147f
C4274 w_4660_n6791.n149 vss 0.069153f
C4275 w_4660_n6791.t28 vss 0.031147f
C4276 w_4660_n6791.t183 vss 0.031147f
C4277 w_4660_n6791.n150 vss 0.07032f
C4278 w_4660_n6791.t139 vss 0.031147f
C4279 w_4660_n6791.t390 vss 0.031147f
C4280 w_4660_n6791.n151 vss 0.069153f
C4281 w_4660_n6791.n152 vss 0.90734f
C4282 w_4660_n6791.n153 vss 0.036697f
C4283 w_4660_n6791.n154 vss 0.008764f
C4284 w_4660_n6791.n155 vss 0.008764f
C4285 w_4660_n6791.n156 vss 0.008764f
C4286 w_4660_n6791.n157 vss 0.064443f
C4287 w_4660_n6791.n158 vss 0.008764f
C4288 w_4660_n6791.n159 vss 0.008764f
C4289 w_4660_n6791.n160 vss 0.008764f
C4290 w_4660_n6791.n161 vss 0.064443f
C4291 w_4660_n6791.n162 vss 0.008764f
C4292 w_4660_n6791.n163 vss 0.008764f
C4293 w_4660_n6791.n164 vss 0.008764f
C4294 w_4660_n6791.n165 vss 0.032221f
C4295 w_4660_n6791.n166 vss 0.008764f
C4296 w_4660_n6791.n167 vss 0.008764f
C4297 w_4660_n6791.n168 vss 0.008764f
C4298 w_4660_n6791.n169 vss 0.064443f
C4299 w_4660_n6791.n170 vss 0.008764f
C4300 w_4660_n6791.n171 vss 0.032221f
C4301 w_4660_n6791.n172 vss 0.008764f
C4302 w_4660_n6791.n173 vss 0.008764f
C4303 w_4660_n6791.n174 vss 0.008764f
C4304 w_4660_n6791.n175 vss 0.064443f
C4305 w_4660_n6791.n176 vss 0.008764f
C4306 w_4660_n6791.n177 vss 0.032221f
C4307 w_4660_n6791.n178 vss 0.008764f
C4308 w_4660_n6791.n179 vss 0.008764f
C4309 w_4660_n6791.n180 vss 0.008764f
C4310 w_4660_n6791.n181 vss 0.064443f
C4311 w_4660_n6791.n182 vss 0.008764f
C4312 w_4660_n6791.n183 vss 0.008764f
C4313 w_4660_n6791.n184 vss 0.008764f
C4314 w_4660_n6791.n185 vss 0.064443f
C4315 w_4660_n6791.n186 vss 0.008764f
C4316 w_4660_n6791.n187 vss 0.040277f
C4317 w_4660_n6791.n188 vss 0.008764f
C4318 w_4660_n6791.n189 vss 0.008764f
C4319 w_4660_n6791.n190 vss 0.008764f
C4320 w_4660_n6791.n191 vss 0.064443f
C4321 w_4660_n6791.n192 vss 0.008764f
C4322 w_4660_n6791.n193 vss 0.008764f
C4323 w_4660_n6791.n194 vss 0.032221f
C4324 w_4660_n6791.n195 vss 0.008764f
C4325 w_4660_n6791.n196 vss 0.032221f
C4326 w_4660_n6791.n197 vss 0.008764f
C4327 w_4660_n6791.n198 vss 0.008764f
C4328 w_4660_n6791.n199 vss 0.008764f
C4329 w_4660_n6791.n200 vss 0.064443f
C4330 w_4660_n6791.n201 vss 0.008764f
C4331 w_4660_n6791.n202 vss 0.032221f
C4332 w_4660_n6791.n203 vss 0.008764f
C4333 w_4660_n6791.n204 vss 0.008764f
C4334 w_4660_n6791.n205 vss 0.008764f
C4335 w_4660_n6791.n206 vss 0.064443f
C4336 w_4660_n6791.n207 vss 0.008764f
C4337 w_4660_n6791.n208 vss 0.034907f
C4338 w_4660_n6791.n209 vss 0.008764f
C4339 w_4660_n6791.n210 vss 0.008764f
C4340 w_4660_n6791.n211 vss 0.008764f
C4341 w_4660_n6791.n212 vss 0.064443f
C4342 w_4660_n6791.n213 vss 0.008764f
C4343 w_4660_n6791.n214 vss 0.008764f
C4344 w_4660_n6791.n215 vss 0.032221f
C4345 w_4660_n6791.n216 vss 0.008764f
C4346 w_4660_n6791.n217 vss 0.032221f
C4347 w_4660_n6791.n218 vss 0.008764f
C4348 w_4660_n6791.n219 vss 0.008764f
C4349 w_4660_n6791.n220 vss 0.008764f
C4350 w_4660_n6791.n221 vss 0.064443f
C4351 w_4660_n6791.n222 vss 0.008764f
C4352 w_4660_n6791.n223 vss 0.032221f
C4353 w_4660_n6791.n224 vss 0.008764f
C4354 w_4660_n6791.n225 vss 0.008764f
C4355 w_4660_n6791.n226 vss 0.008764f
C4356 w_4660_n6791.n227 vss 0.064443f
C4357 w_4660_n6791.n228 vss 0.008764f
C4358 w_4660_n6791.n229 vss 0.032221f
C4359 w_4660_n6791.n230 vss 0.008764f
C4360 w_4660_n6791.n231 vss 0.008764f
C4361 w_4660_n6791.n232 vss 0.006817f
C4362 w_4660_n6791.n233 vss 0.064443f
C4363 w_4660_n6791.n234 vss 0.00633f
C4364 w_4660_n6791.t79 vss 2.64882f
C4365 w_4660_n6791.n235 vss -0.361891f
C4366 w_4660_n6791.n236 vss -0.361891f
C4367 w_4660_n6791.n237 vss -0.361891f
C4368 w_4660_n6791.n238 vss 0.479417f
C4369 w_4660_n6791.n239 vss 0.479417f
C4370 w_4660_n6791.n240 vss -0.361891f
C4371 w_4660_n6791.n241 vss -0.361891f
C4372 w_4660_n6791.n242 vss 0.006817f
C4373 w_4660_n6791.n243 vss -0.361891f
C4374 w_4660_n6791.n244 vss 0.479417f
C4375 w_4660_n6791.n245 vss -0.361891f
C4376 w_4660_n6791.t148 vss 3.53177f
C4377 w_4660_n6791.t109 vss 3.53177f
C4378 w_4660_n6791.t92 vss 3.53177f
C4379 w_4660_n6791.t13 vss 3.53177f
C4380 w_4660_n6791.t130 vss 3.53177f
C4381 w_4660_n6791.t45 vss 3.53177f
C4382 w_4660_n6791.t39 vss 3.53177f
C4383 w_4660_n6791.t5 vss 3.53177f
C4384 w_4660_n6791.t64 vss 3.53177f
C4385 w_4660_n6791.t23 vss 3.53177f
C4386 w_4660_n6791.t52 vss 3.53177f
C4387 w_4660_n6791.t41 vss 3.53177f
C4388 w_4660_n6791.t141 vss 3.53177f
C4389 w_4660_n6791.t15 vss 3.53177f
C4390 w_4660_n6791.t98 vss 3.53177f
C4391 w_4660_n6791.t72 vss 3.53177f
C4392 w_4660_n6791.t35 vss 3.53177f
C4393 w_4660_n6791.t0 vss 3.53177f
C4394 w_4660_n6791.t50 vss 3.53177f
C4395 w_4660_n6791.t168 vss 3.53177f
C4396 w_4660_n6791.t112 vss 3.53177f
C4397 w_4660_n6791.t11 vss 3.53177f
C4398 w_4660_n6791.t163 vss 3.53177f
C4399 w_4660_n6791.t43 vss 2.64882f
C4400 w_4660_n6791.n246 vss 0.48173f
C4401 w_4660_n6791.n247 vss 0.294894f
C4402 w_4660_n6791.n248 vss 0.009022f
C4403 w_4660_n6791.n249 vss 0.035229f
C4404 w_4660_n6791.n250 vss 0.008764f
C4405 w_4660_n6791.n251 vss 0.061865f
C4406 w_4660_n6791.n252 vss 0.010849f
C4407 w_4660_n6791.n253 vss 0.028693f
C4408 w_4660_n6791.n254 vss 0.154304f
C4409 w_4660_n6791.n255 vss 0.010849f
C4410 w_4660_n6791.n256 vss 0.022123f
C4411 w_4660_n6791.n257 vss 0.010849f
C4412 w_4660_n6791.n258 vss 0.008764f
C4413 w_4660_n6791.n259 vss 0.008764f
C4414 w_4660_n6791.n260 vss 0.008764f
C4415 w_4660_n6791.n261 vss 0.061865f
C4416 w_4660_n6791.n262 vss 0.009022f
C4417 w_4660_n6791.n263 vss 0.008764f
C4418 w_4660_n6791.n264 vss 0.008764f
C4419 w_4660_n6791.n265 vss 0.061865f
C4420 w_4660_n6791.n266 vss 0.008764f
C4421 w_4660_n6791.n267 vss 0.008764f
C4422 w_4660_n6791.n268 vss 0.008764f
C4423 w_4660_n6791.n269 vss 0.061865f
C4424 w_4660_n6791.n270 vss 0.009022f
C4425 w_4660_n6791.n271 vss 0.008764f
C4426 w_4660_n6791.n272 vss 0.008764f
C4427 w_4660_n6791.n273 vss 0.061865f
C4428 w_4660_n6791.n274 vss 0.008764f
C4429 w_4660_n6791.n275 vss 0.008764f
C4430 w_4660_n6791.n276 vss 0.008764f
C4431 w_4660_n6791.n277 vss 0.061865f
C4432 w_4660_n6791.n278 vss 0.004507f
C4433 w_4660_n6791.n279 vss 0.008764f
C4434 w_4660_n6791.n280 vss 0.008764f
C4435 w_4660_n6791.n281 vss 0.061865f
C4436 w_4660_n6791.n282 vss 0.008764f
C4437 w_4660_n6791.n283 vss 0.008764f
C4438 w_4660_n6791.n284 vss 0.008764f
C4439 w_4660_n6791.n285 vss 0.061865f
C4440 w_4660_n6791.n286 vss 0.008582f
C4441 w_4660_n6791.n287 vss 0.009022f
C4442 w_4660_n6791.n288 vss 0.008764f
C4443 w_4660_n6791.n289 vss 0.008764f
C4444 w_4660_n6791.n290 vss 0.061865f
C4445 w_4660_n6791.n291 vss 0.008764f
C4446 w_4660_n6791.n292 vss 0.008764f
C4447 w_4660_n6791.n293 vss 0.008764f
C4448 w_4660_n6791.n294 vss 0.061865f
C4449 w_4660_n6791.n295 vss 0.009022f
C4450 w_4660_n6791.n296 vss 0.008764f
C4451 w_4660_n6791.n297 vss 0.008764f
C4452 w_4660_n6791.n298 vss 0.061865f
C4453 w_4660_n6791.n299 vss 0.111491f
C4454 w_4660_n6791.n300 vss 0.008764f
C4455 w_4660_n6791.n301 vss 0.011345f
C4456 w_4660_n6791.n302 vss 0.008764f
C4457 w_4660_n6791.n303 vss 0.032221f
C4458 w_4660_n6791.n304 vss 0.008764f
C4459 w_4660_n6791.n305 vss 0.059968f
C4460 w_4660_n6791.n306 vss 0.008764f
C4461 w_4660_n6791.n307 vss 0.064443f
C4462 w_4660_n6791.n308 vss 0.008764f
C4463 w_4660_n6791.n309 vss 0.008764f
C4464 w_4660_n6791.t410 vss 0.031147f
C4465 w_4660_n6791.t435 vss 0.031147f
C4466 w_4660_n6791.n310 vss 0.069153f
C4467 w_4660_n6791.t14 vss 0.031147f
C4468 w_4660_n6791.t93 vss 0.031147f
C4469 w_4660_n6791.n311 vss 0.069153f
C4470 w_4660_n6791.t134 vss 0.031147f
C4471 w_4660_n6791.t131 vss 0.031147f
C4472 w_4660_n6791.n312 vss 0.069153f
C4473 w_4660_n6791.n313 vss 0.549171f
C4474 w_4660_n6791.n314 vss 0.059968f
C4475 w_4660_n6791.n315 vss 0.008764f
C4476 w_4660_n6791.n316 vss 0.008764f
C4477 w_4660_n6791.n317 vss 0.008764f
C4478 w_4660_n6791.n318 vss 0.064443f
C4479 w_4660_n6791.n319 vss 0.008764f
C4480 w_4660_n6791.n320 vss 0.045647f
C4481 w_4660_n6791.n321 vss 0.008764f
C4482 w_4660_n6791.n322 vss 0.064443f
C4483 w_4660_n6791.n323 vss 0.032221f
C4484 w_4660_n6791.n324 vss 0.008764f
C4485 w_4660_n6791.n325 vss 0.032221f
C4486 w_4660_n6791.n326 vss 0.008764f
C4487 w_4660_n6791.n327 vss 0.008764f
C4488 w_4660_n6791.n328 vss 0.064443f
C4489 w_4660_n6791.n329 vss 0.008764f
C4490 w_4660_n6791.n330 vss 0.008764f
C4491 w_4660_n6791.t143 vss 0.031147f
C4492 w_4660_n6791.t65 vss 0.031147f
C4493 w_4660_n6791.n331 vss 0.069153f
C4494 w_4660_n6791.t42 vss 0.031147f
C4495 w_4660_n6791.t137 vss 0.031147f
C4496 w_4660_n6791.n332 vss 0.069153f
C4497 w_4660_n6791.t55 vss 0.031147f
C4498 w_4660_n6791.t142 vss 0.031147f
C4499 w_4660_n6791.n333 vss 0.069153f
C4500 w_4660_n6791.n334 vss 0.549171f
C4501 w_4660_n6791.n335 vss 0.056388f
C4502 w_4660_n6791.n336 vss 0.008764f
C4503 w_4660_n6791.n337 vss 0.008764f
C4504 w_4660_n6791.n338 vss 0.008764f
C4505 w_4660_n6791.n339 vss 0.064443f
C4506 w_4660_n6791.n340 vss 0.008764f
C4507 w_4660_n6791.n341 vss 0.049227f
C4508 w_4660_n6791.n342 vss 0.008764f
C4509 w_4660_n6791.n343 vss 0.064443f
C4510 w_4660_n6791.n344 vss 0.032221f
C4511 w_4660_n6791.n345 vss 0.008764f
C4512 w_4660_n6791.n346 vss 0.032221f
C4513 w_4660_n6791.n347 vss 0.008764f
C4514 w_4660_n6791.n348 vss 0.064443f
C4515 w_4660_n6791.n349 vss 0.008764f
C4516 w_4660_n6791.n350 vss 0.032221f
C4517 w_4660_n6791.n351 vss 0.008764f
C4518 w_4660_n6791.n352 vss 0.043857f
C4519 w_4660_n6791.n353 vss 0.008764f
C4520 w_4660_n6791.n354 vss 0.064443f
C4521 w_4660_n6791.n355 vss 0.008764f
C4522 w_4660_n6791.n356 vss 0.008764f
C4523 w_4660_n6791.t415 vss 0.031147f
C4524 w_4660_n6791.t165 vss 0.031147f
C4525 w_4660_n6791.n357 vss 0.069153f
C4526 w_4660_n6791.t12 vss 0.031147f
C4527 w_4660_n6791.t113 vss 0.031147f
C4528 w_4660_n6791.n358 vss 0.069153f
C4529 w_4660_n6791.t450 vss 0.031147f
C4530 w_4660_n6791.t409 vss 0.031147f
C4531 w_4660_n6791.n359 vss 0.069153f
C4532 w_4660_n6791.n360 vss 0.549171f
C4533 w_4660_n6791.n361 vss 0.043857f
C4534 w_4660_n6791.n362 vss 0.008764f
C4535 w_4660_n6791.n363 vss 0.008764f
C4536 w_4660_n6791.n364 vss 0.008764f
C4537 w_4660_n6791.n365 vss 0.061758f
C4538 w_4660_n6791.n366 vss 0.006817f
C4539 w_4660_n6791.n367 vss 0.064443f
C4540 w_4660_n6791.n368 vss 0.032221f
C4541 w_4660_n6791.n369 vss 0.008764f
C4542 w_4660_n6791.n370 vss 0.038487f
C4543 w_4660_n6791.n371 vss 0.008764f
C4544 w_4660_n6791.n372 vss 0.064443f
C4545 w_4660_n6791.n373 vss 0.032221f
C4546 w_4660_n6791.n374 vss 0.008764f
C4547 w_4660_n6791.n375 vss 0.032221f
C4548 w_4660_n6791.n376 vss 0.008764f
C4549 w_4660_n6791.n377 vss 0.056388f
C4550 w_4660_n6791.n378 vss 0.008764f
C4551 w_4660_n6791.n379 vss 0.064443f
C4552 w_4660_n6791.n380 vss 0.008764f
C4553 w_4660_n6791.n381 vss 0.008764f
C4554 w_4660_n6791.t449 vss 0.031147f
C4555 w_4660_n6791.t402 vss 0.031147f
C4556 w_4660_n6791.n382 vss 0.069153f
C4557 w_4660_n6791.t152 vss 0.031147f
C4558 w_4660_n6791.t462 vss 0.031147f
C4559 w_4660_n6791.n383 vss 0.069153f
C4560 w_4660_n6791.t445 vss 0.031147f
C4561 w_4660_n6791.t121 vss 0.031147f
C4562 w_4660_n6791.n384 vss 0.069153f
C4563 w_4660_n6791.n385 vss 0.549171f
C4564 w_4660_n6791.n386 vss 0.063548f
C4565 w_4660_n6791.n387 vss 0.008764f
C4566 w_4660_n6791.n388 vss 0.008764f
C4567 w_4660_n6791.n389 vss 0.008764f
C4568 w_4660_n6791.n390 vss 0.064443f
C4569 w_4660_n6791.n391 vss 0.008764f
C4570 w_4660_n6791.n392 vss 0.042067f
C4571 w_4660_n6791.n393 vss 0.008764f
C4572 w_4660_n6791.n394 vss 0.064443f
C4573 w_4660_n6791.n395 vss 0.032221f
C4574 w_4660_n6791.n396 vss 0.008764f
C4575 w_4660_n6791.n397 vss 0.032221f
C4576 w_4660_n6791.n398 vss 0.008764f
C4577 w_4660_n6791.n399 vss 0.059968f
C4578 w_4660_n6791.n400 vss 0.008764f
C4579 w_4660_n6791.n401 vss 0.064443f
C4580 w_4660_n6791.n402 vss 0.008764f
C4581 w_4660_n6791.n403 vss 0.008764f
C4582 w_4660_n6791.t105 vss 0.031147f
C4583 w_4660_n6791.t442 vss 0.031147f
C4584 w_4660_n6791.n404 vss 0.069153f
C4585 w_4660_n6791.t108 vss 0.031147f
C4586 w_4660_n6791.t427 vss 0.031147f
C4587 w_4660_n6791.n405 vss 0.069153f
C4588 w_4660_n6791.t429 vss 0.031147f
C4589 w_4660_n6791.t180 vss 0.031147f
C4590 w_4660_n6791.n406 vss 0.069153f
C4591 w_4660_n6791.n407 vss 0.549171f
C4592 w_4660_n6791.n408 vss 0.059968f
C4593 w_4660_n6791.n409 vss 0.008764f
C4594 w_4660_n6791.n410 vss 0.008764f
C4595 w_4660_n6791.n411 vss 0.008764f
C4596 w_4660_n6791.n412 vss 0.064443f
C4597 w_4660_n6791.n413 vss 0.008764f
C4598 w_4660_n6791.n414 vss 0.045647f
C4599 w_4660_n6791.n415 vss 0.008764f
C4600 w_4660_n6791.n416 vss 0.064443f
C4601 w_4660_n6791.n417 vss 0.032221f
C4602 w_4660_n6791.n418 vss 0.008764f
C4603 w_4660_n6791.n419 vss 0.032221f
C4604 w_4660_n6791.n420 vss 0.008764f
C4605 w_4660_n6791.n421 vss 0.008764f
C4606 w_4660_n6791.n422 vss 0.064443f
C4607 w_4660_n6791.n423 vss 0.008764f
C4608 w_4660_n6791.n424 vss 0.008764f
C4609 w_4660_n6791.t456 vss 0.031147f
C4610 w_4660_n6791.t469 vss 0.031147f
C4611 w_4660_n6791.n425 vss 0.069153f
C4612 w_4660_n6791.t96 vss 0.031147f
C4613 w_4660_n6791.t404 vss 0.031147f
C4614 w_4660_n6791.n426 vss 0.069153f
C4615 w_4660_n6791.t136 vss 0.120265f
C4616 w_4660_n6791.t159 vss 0.121336f
C4617 w_4660_n6791.t123 vss 0.120265f
C4618 w_4660_n6791.n427 vss 0.875204f
C4619 w_4660_n6791.t463 vss 0.121336f
C4620 w_4660_n6791.t221 vss 0.120256f
C4621 w_4660_n6791.n428 vss 0.875654f
C4622 w_4660_n6791.t220 vss 0.121325f
C4623 w_4660_n6791.t273 vss 0.120265f
C4624 w_4660_n6791.n429 vss 0.875655f
C4625 w_4660_n6791.n430 vss 0.081778f
C4626 w_4660_n6791.n431 vss 0.081778f
C4627 w_4660_n6791.n432 vss 0.081778f
C4628 w_4660_n6791.n433 vss 0.081273f
C4629 w_4660_n6791.n435 vss 0.081273f
C4630 w_4660_n6791.n436 vss 0.081778f
C4631 w_4660_n6791.n437 vss 0.081778f
C4632 w_4660_n6791.n445 vss 0.081778f
C4633 w_4660_n6791.t349 vss 0.120265f
C4634 w_4660_n6791.n446 vss 0.06512f
C4635 w_4660_n6791.n447 vss 0.072327f
C4636 w_4660_n6791.n448 vss 0.011345f
C4637 w_4660_n6791.n449 vss 0.064443f
C4638 w_4660_n6791.n450 vss 0.011345f
C4639 w_4660_n6791.n451 vss 0.063443f
C4640 w_4660_n6791.n452 vss 0.48173f
C4641 w_4660_n6791.t83 vss 3.53177f
C4642 w_4660_n6791.t88 vss 3.53177f
C4643 w_4660_n6791.t67 vss 3.53177f
C4644 w_4660_n6791.t37 vss 3.53177f
C4645 w_4660_n6791.t86 vss 3.53177f
C4646 w_4660_n6791.t102 vss 3.53177f
C4647 w_4660_n6791.t62 vss 3.53177f
C4648 w_4660_n6791.t30 vss 3.53177f
C4649 w_4660_n6791.t47 vss 3.53177f
C4650 w_4660_n6791.t70 vss 3.53177f
C4651 w_4660_n6791.t2 vss 3.53177f
C4652 w_4660_n6791.t33 vss 3.53177f
C4653 w_4660_n6791.t7 vss 3.53177f
C4654 w_4660_n6791.t94 vss 3.53177f
C4655 w_4660_n6791.t107 vss 3.53177f
C4656 w_4660_n6791.t60 vss 3.53177f
C4657 w_4660_n6791.t118 vss 3.53177f
C4658 w_4660_n6791.t144 vss 3.53177f
C4659 w_4660_n6791.t240 vss 3.53177f
C4660 w_4660_n6791.t166 vss 3.53177f
C4661 w_4660_n6791.t25 vss 3.53177f
C4662 w_4660_n6791.t291 vss 3.53177f
C4663 w_4660_n6791.t17 vss 3.53177f
C4664 w_4660_n6791.t122 vss 4.35485f
C4665 w_4660_n6791.n453 vss 0.005426f
C4666 w_4660_n6791.n454 vss 0.009022f
C4667 w_4660_n6791.n455 vss 0.049836f
C4668 w_4660_n6791.n456 vss 0.008764f
C4669 w_4660_n6791.n457 vss 0.061865f
C4670 w_4660_n6791.n458 vss 0.168931f
C4671 w_4660_n6791.n459 vss 0.008764f
C4672 w_4660_n6791.n460 vss 0.061865f
C4673 w_4660_n6791.n461 vss 0.009022f
C4674 w_4660_n6791.n462 vss 0.008764f
C4675 w_4660_n6791.n463 vss 0.061865f
C4676 w_4660_n6791.n464 vss 0.008764f
C4677 w_4660_n6791.n465 vss 0.009022f
C4678 w_4660_n6791.n466 vss 0.061865f
C4679 w_4660_n6791.n467 vss 0.008764f
C4680 w_4660_n6791.n468 vss 0.008764f
C4681 w_4660_n6791.n469 vss 0.061865f
C4682 w_4660_n6791.n470 vss 0.008764f
C4683 w_4660_n6791.n471 vss 0.008764f
C4684 w_4660_n6791.n472 vss 0.009022f
C4685 w_4660_n6791.n473 vss 0.061865f
C4686 w_4660_n6791.n474 vss 0.008764f
C4687 w_4660_n6791.n475 vss 0.008764f
C4688 w_4660_n6791.n476 vss 0.008764f
C4689 w_4660_n6791.n477 vss 0.061865f
C4690 w_4660_n6791.n478 vss 0.008764f
C4691 w_4660_n6791.n479 vss 0.008764f
C4692 w_4660_n6791.n480 vss 0.009022f
C4693 w_4660_n6791.n481 vss 0.061865f
C4694 w_4660_n6791.n482 vss 0.008764f
C4695 w_4660_n6791.n483 vss 0.008764f
C4696 w_4660_n6791.n484 vss 0.008764f
C4697 w_4660_n6791.n485 vss 0.061865f
C4698 w_4660_n6791.n486 vss 0.008764f
C4699 w_4660_n6791.n487 vss 0.008764f
C4700 w_4660_n6791.n488 vss 0.009022f
C4701 w_4660_n6791.n489 vss 0.061865f
C4702 w_4660_n6791.n490 vss 0.008764f
C4703 w_4660_n6791.n491 vss 0.008764f
C4704 w_4660_n6791.n492 vss 0.008764f
C4705 w_4660_n6791.n493 vss 0.061865f
C4706 w_4660_n6791.n494 vss 0.008764f
C4707 w_4660_n6791.n495 vss 0.008764f
C4708 w_4660_n6791.n496 vss 0.009022f
C4709 w_4660_n6791.n497 vss 0.061865f
C4710 w_4660_n6791.n498 vss 0.008764f
C4711 w_4660_n6791.n499 vss 0.008764f
C4712 w_4660_n6791.n500 vss 0.008764f
C4713 w_4660_n6791.n501 vss 0.061865f
C4714 w_4660_n6791.n502 vss 0.008764f
C4715 w_4660_n6791.n503 vss 0.008764f
C4716 w_4660_n6791.n504 vss 0.008764f
C4717 w_4660_n6791.n505 vss 0.032221f
C4718 w_4660_n6791.n506 vss 0.010661f
C4719 w_4660_n6791.n507 vss 0.008764f
C4720 w_4660_n6791.n508 vss 0.008764f
C4721 w_4660_n6791.n509 vss 0.059968f
C4722 w_4660_n6791.n510 vss 0.008764f
C4723 w_4660_n6791.n511 vss 0.032221f
C4724 w_4660_n6791.n512 vss 0.008764f
C4725 w_4660_n6791.n513 vss 0.008764f
C4726 w_4660_n6791.n514 vss 0.064443f
C4727 w_4660_n6791.n515 vss 0.008764f
C4728 w_4660_n6791.n516 vss 0.008764f
C4729 w_4660_n6791.n517 vss 0.008764f
C4730 w_4660_n6791.n518 vss 0.008764f
C4731 w_4660_n6791.n519 vss 0.036697f
C4732 w_4660_n6791.n520 vss 0.008764f
C4733 w_4660_n6791.n521 vss 0.032221f
C4734 w_4660_n6791.n522 vss 0.008764f
C4735 w_4660_n6791.n523 vss 0.008764f
C4736 w_4660_n6791.n524 vss 0.064443f
C4737 w_4660_n6791.n525 vss 0.008764f
C4738 w_4660_n6791.n526 vss 0.008764f
C4739 w_4660_n6791.n527 vss 0.008764f
C4740 w_4660_n6791.n528 vss 0.032221f
C4741 w_4660_n6791.n529 vss 0.008764f
C4742 w_4660_n6791.n530 vss 0.008764f
C4743 w_4660_n6791.n531 vss 0.008764f
C4744 w_4660_n6791.n532 vss 0.054598f
C4745 w_4660_n6791.n533 vss 0.008764f
C4746 w_4660_n6791.n534 vss 0.032221f
C4747 w_4660_n6791.n535 vss 0.008764f
C4748 w_4660_n6791.n536 vss 0.008764f
C4749 w_4660_n6791.n537 vss 0.064443f
C4750 w_4660_n6791.n538 vss 0.008764f
C4751 w_4660_n6791.n539 vss 0.008764f
C4752 w_4660_n6791.n540 vss 0.008764f
C4753 w_4660_n6791.n541 vss 0.008764f
C4754 w_4660_n6791.n542 vss 0.008764f
C4755 w_4660_n6791.n543 vss 0.008764f
C4756 w_4660_n6791.n544 vss 0.064443f
C4757 w_4660_n6791.n545 vss 0.008764f
C4758 w_4660_n6791.n546 vss 0.008764f
C4759 w_4660_n6791.n547 vss 0.008764f
C4760 w_4660_n6791.n548 vss 0.032221f
C4761 w_4660_n6791.n549 vss 0.008764f
C4762 w_4660_n6791.n550 vss 0.008764f
C4763 w_4660_n6791.n551 vss 0.008764f
C4764 w_4660_n6791.n552 vss 0.008764f
C4765 w_4660_n6791.n553 vss 0.049227f
C4766 w_4660_n6791.n554 vss 0.008764f
C4767 w_4660_n6791.n555 vss 0.032221f
C4768 w_4660_n6791.n556 vss 0.008764f
C4769 w_4660_n6791.n557 vss 0.008764f
C4770 w_4660_n6791.n558 vss 0.064443f
C4771 w_4660_n6791.n559 vss 0.008764f
C4772 w_4660_n6791.n560 vss 0.008764f
C4773 w_4660_n6791.n561 vss 0.008764f
C4774 w_4660_n6791.n562 vss 0.008764f
C4775 w_4660_n6791.n563 vss 0.032221f
C4776 w_4660_n6791.n564 vss 0.008764f
C4777 w_4660_n6791.n565 vss 0.008764f
C4778 w_4660_n6791.n566 vss 0.008764f
C4779 w_4660_n6791.n567 vss 0.064443f
C4780 w_4660_n6791.n568 vss 0.008764f
C4781 w_4660_n6791.n569 vss 0.008764f
C4782 w_4660_n6791.n570 vss 0.008764f
C4783 w_4660_n6791.n571 vss 0.032221f
C4784 w_4660_n6791.n572 vss 0.008764f
C4785 w_4660_n6791.n573 vss 0.008764f
C4786 w_4660_n6791.n574 vss 0.008764f
C4787 w_4660_n6791.n575 vss 0.008764f
C4788 w_4660_n6791.n576 vss 0.043857f
C4789 w_4660_n6791.n577 vss 0.008764f
C4790 w_4660_n6791.n578 vss 0.032221f
C4791 w_4660_n6791.n579 vss 0.008764f
C4792 w_4660_n6791.n580 vss 0.008764f
C4793 w_4660_n6791.n581 vss 0.064443f
C4794 w_4660_n6791.n582 vss 0.008764f
C4795 w_4660_n6791.n583 vss 0.008764f
C4796 w_4660_n6791.n584 vss 0.008764f
C4797 w_4660_n6791.n585 vss 0.008764f
C4798 w_4660_n6791.n586 vss 0.032221f
C4799 w_4660_n6791.n587 vss 0.008764f
C4800 w_4660_n6791.n588 vss 0.008764f
C4801 w_4660_n6791.n589 vss 0.008764f
C4802 w_4660_n6791.n590 vss 0.061758f
C4803 w_4660_n6791.n591 vss 0.006817f
C4804 w_4660_n6791.n592 vss 0.032221f
C4805 w_4660_n6791.n593 vss 0.008764f
C4806 w_4660_n6791.n594 vss 0.008764f
C4807 w_4660_n6791.n595 vss 0.006817f
C4808 w_4660_n6791.n596 vss 0.004382f
C4809 w_4660_n6791.n597 vss 0.00633f
C4810 w_4660_n6791.n598 vss 0.038487f
C4811 w_4660_n6791.n599 vss 0.00633f
C4812 w_4660_n6791.n600 vss 0.008764f
C4813 w_4660_n6791.n601 vss 0.032221f
C4814 w_4660_n6791.n602 vss 0.008764f
C4815 w_4660_n6791.n603 vss 0.008764f
C4816 w_4660_n6791.n604 vss 0.064443f
C4817 w_4660_n6791.n605 vss 0.008764f
C4818 w_4660_n6791.n606 vss 0.008764f
C4819 w_4660_n6791.n607 vss 0.008764f
C4820 w_4660_n6791.n608 vss 0.008764f
C4821 w_4660_n6791.n609 vss 0.032221f
C4822 w_4660_n6791.n610 vss 0.008764f
C4823 w_4660_n6791.n611 vss 0.008764f
C4824 w_4660_n6791.n612 vss 0.008764f
C4825 w_4660_n6791.n613 vss 0.056388f
C4826 w_4660_n6791.n614 vss 0.008764f
C4827 w_4660_n6791.n615 vss 0.032221f
C4828 w_4660_n6791.n616 vss 0.008764f
C4829 w_4660_n6791.n617 vss 0.008764f
C4830 w_4660_n6791.n618 vss 0.064443f
C4831 w_4660_n6791.n619 vss 0.008764f
C4832 w_4660_n6791.n620 vss 0.008764f
C4833 w_4660_n6791.n621 vss 0.008764f
C4834 w_4660_n6791.n622 vss 0.008764f
C4835 w_4660_n6791.n623 vss 0.008764f
C4836 w_4660_n6791.n624 vss 0.008764f
C4837 w_4660_n6791.n625 vss 0.064443f
C4838 w_4660_n6791.n626 vss 0.008764f
C4839 w_4660_n6791.n627 vss 0.008764f
C4840 w_4660_n6791.n628 vss 0.008764f
C4841 w_4660_n6791.n629 vss 0.032221f
C4842 w_4660_n6791.n630 vss 0.008764f
C4843 w_4660_n6791.n631 vss 0.008764f
C4844 w_4660_n6791.n632 vss 0.008764f
C4845 w_4660_n6791.n633 vss 0.051017f
C4846 w_4660_n6791.n634 vss 0.008764f
C4847 w_4660_n6791.n635 vss 0.032221f
C4848 w_4660_n6791.n636 vss 0.008764f
C4849 w_4660_n6791.n637 vss 0.008764f
C4850 w_4660_n6791.n638 vss 0.064443f
C4851 w_4660_n6791.n639 vss 0.008764f
C4852 w_4660_n6791.n640 vss 0.008764f
C4853 w_4660_n6791.n641 vss 0.008764f
C4854 w_4660_n6791.n642 vss 0.008764f
C4855 w_4660_n6791.n643 vss 0.032221f
C4856 w_4660_n6791.n644 vss 0.008764f
C4857 w_4660_n6791.n645 vss 0.008764f
C4858 w_4660_n6791.n646 vss 0.008764f
C4859 w_4660_n6791.n647 vss 0.064443f
C4860 w_4660_n6791.n648 vss 0.008764f
C4861 w_4660_n6791.n649 vss 0.008764f
C4862 w_4660_n6791.n650 vss 0.008764f
C4863 w_4660_n6791.n651 vss 0.032221f
C4864 w_4660_n6791.n652 vss 0.008764f
C4865 w_4660_n6791.n653 vss 0.008764f
C4866 w_4660_n6791.n654 vss 0.008764f
C4867 w_4660_n6791.n655 vss 0.008764f
C4868 w_4660_n6791.n656 vss 0.045647f
C4869 w_4660_n6791.n657 vss 0.008764f
C4870 w_4660_n6791.n658 vss 0.032221f
C4871 w_4660_n6791.n659 vss 0.008764f
C4872 w_4660_n6791.n660 vss 0.008764f
C4873 w_4660_n6791.n661 vss 0.064443f
C4874 w_4660_n6791.n662 vss 0.008764f
C4875 w_4660_n6791.n663 vss 0.008764f
C4876 w_4660_n6791.n664 vss 0.008764f
C4877 w_4660_n6791.n665 vss 0.008764f
C4878 w_4660_n6791.n666 vss 0.032221f
C4879 w_4660_n6791.n667 vss 0.008764f
C4880 w_4660_n6791.n668 vss 0.008764f
C4881 w_4660_n6791.n669 vss 0.008764f
C4882 w_4660_n6791.n670 vss 0.008764f
C4883 w_4660_n6791.n671 vss 0.008764f
C4884 w_4660_n6791.n672 vss 0.008764f
C4885 w_4660_n6791.n673 vss 0.064443f
C4886 w_4660_n6791.n674 vss 0.008764f
C4887 w_4660_n6791.n675 vss 0.008764f
C4888 w_4660_n6791.n676 vss 0.008764f
C4889 w_4660_n6791.n677 vss 0.008764f
C4890 w_4660_n6791.n678 vss 0.040277f
C4891 w_4660_n6791.n679 vss 0.008764f
C4892 w_4660_n6791.n680 vss 0.032221f
C4893 w_4660_n6791.n681 vss 0.008764f
C4894 w_4660_n6791.n682 vss 0.008764f
C4895 w_4660_n6791.n683 vss 0.064443f
C4896 w_4660_n6791.n684 vss 0.009312f
C4897 w_4660_n6791.n685 vss 0.008764f
C4898 w_4660_n6791.n686 vss 0.008764f
C4899 w_4660_n6791.t447 vss 0.121336f
C4900 w_4660_n6791.t257 vss 0.120256f
C4901 w_4660_n6791.t110 vss 0.031147f
C4902 w_4660_n6791.t149 vss 0.031147f
C4903 w_4660_n6791.n687 vss 0.07032f
C4904 w_4660_n6791.t270 vss 0.031147f
C4905 w_4660_n6791.t252 vss 0.031147f
C4906 w_4660_n6791.n688 vss 0.069142f
C4907 w_4660_n6791.t471 vss 0.031147f
C4908 w_4660_n6791.t186 vss 0.031147f
C4909 w_4660_n6791.n689 vss 0.07032f
C4910 w_4660_n6791.t344 vss 0.031147f
C4911 w_4660_n6791.t197 vss 0.031147f
C4912 w_4660_n6791.n690 vss 0.069142f
C4913 w_4660_n6791.t181 vss 0.031147f
C4914 w_4660_n6791.t138 vss 0.031147f
C4915 w_4660_n6791.n691 vss 0.07032f
C4916 w_4660_n6791.t335 vss 0.031147f
C4917 w_4660_n6791.t339 vss 0.031147f
C4918 w_4660_n6791.n692 vss 0.069142f
C4919 w_4660_n6791.t420 vss 0.031147f
C4920 w_4660_n6791.t40 vss 0.031147f
C4921 w_4660_n6791.n693 vss 0.07032f
C4922 w_4660_n6791.t260 vss 0.031147f
C4923 w_4660_n6791.t329 vss 0.031147f
C4924 w_4660_n6791.n694 vss 0.069142f
C4925 w_4660_n6791.t458 vss 0.031147f
C4926 w_4660_n6791.t389 vss 0.031147f
C4927 w_4660_n6791.n695 vss 0.07032f
C4928 w_4660_n6791.t216 vss 0.031147f
C4929 w_4660_n6791.t201 vss 0.031147f
C4930 w_4660_n6791.n696 vss 0.069142f
C4931 w_4660_n6791.t476 vss 0.031147f
C4932 w_4660_n6791.t53 vss 0.031147f
C4933 w_4660_n6791.n697 vss 0.07032f
C4934 w_4660_n6791.t207 vss 0.031147f
C4935 w_4660_n6791.t210 vss 0.031147f
C4936 w_4660_n6791.n698 vss 0.069142f
C4937 w_4660_n6791.t29 vss 0.031147f
C4938 w_4660_n6791.t454 vss 0.031147f
C4939 w_4660_n6791.n699 vss 0.07032f
C4940 w_4660_n6791.t289 vss 0.031147f
C4941 w_4660_n6791.t205 vss 0.031147f
C4942 w_4660_n6791.n700 vss 0.069142f
C4943 w_4660_n6791.t175 vss 0.031147f
C4944 w_4660_n6791.t172 vss 0.031147f
C4945 w_4660_n6791.n701 vss 0.07032f
C4946 w_4660_n6791.t281 vss 0.031147f
C4947 w_4660_n6791.t285 vss 0.031147f
C4948 w_4660_n6791.n702 vss 0.069142f
C4949 w_4660_n6791.t153 vss 0.031147f
C4950 w_4660_n6791.t185 vss 0.031147f
C4951 w_4660_n6791.n703 vss 0.07032f
C4952 w_4660_n6791.t269 vss 0.031147f
C4953 w_4660_n6791.t277 vss 0.031147f
C4954 w_4660_n6791.n704 vss 0.069142f
C4955 w_4660_n6791.t446 vss 0.031147f
C4956 w_4660_n6791.t51 vss 0.031147f
C4957 w_4660_n6791.n705 vss 0.07032f
C4958 w_4660_n6791.t371 vss 0.031147f
C4959 w_4660_n6791.t231 vss 0.031147f
C4960 w_4660_n6791.n706 vss 0.069142f
C4961 w_4660_n6791.t158 vss 0.031147f
C4962 w_4660_n6791.t170 vss 0.031147f
C4963 w_4660_n6791.n707 vss 0.07032f
C4964 w_4660_n6791.t357 vss 0.031147f
C4965 w_4660_n6791.t362 vss 0.031147f
C4966 w_4660_n6791.n708 vss 0.069142f
C4967 w_4660_n6791.t394 vss 0.031147f
C4968 w_4660_n6791.t178 vss 0.031147f
C4969 w_4660_n6791.n709 vss 0.07032f
C4970 w_4660_n6791.t302 vss 0.031147f
C4971 w_4660_n6791.t350 vss 0.031147f
C4972 w_4660_n6791.n710 vss 0.069142f
C4973 w_4660_n6791.t84 vss 0.031147f
C4974 w_4660_n6791.t80 vss 0.031147f
C4975 w_4660_n6791.n711 vss 0.07032f
C4976 w_4660_n6791.t215 vss 0.031147f
C4977 w_4660_n6791.t219 vss 0.031147f
C4978 w_4660_n6791.n712 vss 0.069142f
C4979 w_4660_n6791.t115 vss 0.031147f
C4980 w_4660_n6791.t421 vss 0.031147f
C4981 w_4660_n6791.n713 vss 0.07032f
C4982 w_4660_n6791.t227 vss 0.031147f
C4983 w_4660_n6791.t238 vss 0.031147f
C4984 w_4660_n6791.n714 vss 0.069142f
C4985 w_4660_n6791.t444 vss 0.031147f
C4986 w_4660_n6791.t59 vss 0.031147f
C4987 w_4660_n6791.n715 vss 0.07032f
C4988 w_4660_n6791.t382 vss 0.031147f
C4989 w_4660_n6791.t387 vss 0.031147f
C4990 w_4660_n6791.n716 vss 0.069142f
C4991 w_4660_n6791.t63 vss 0.031147f
C4992 w_4660_n6791.t103 vss 0.031147f
C4993 w_4660_n6791.n717 vss 0.07032f
C4994 w_4660_n6791.t306 vss 0.031147f
C4995 w_4660_n6791.t309 vss 0.031147f
C4996 w_4660_n6791.n718 vss 0.069142f
C4997 w_4660_n6791.t106 vss 0.031147f
C4998 w_4660_n6791.t399 vss 0.031147f
C4999 w_4660_n6791.n719 vss 0.07032f
C5000 w_4660_n6791.t243 vss 0.031147f
C5001 w_4660_n6791.t299 vss 0.031147f
C5002 w_4660_n6791.n720 vss 0.069142f
C5003 w_4660_n6791.t3 vss 0.031147f
C5004 w_4660_n6791.t439 vss 0.031147f
C5005 w_4660_n6791.n721 vss 0.07032f
C5006 w_4660_n6791.t190 vss 0.031147f
C5007 w_4660_n6791.t230 vss 0.031147f
C5008 w_4660_n6791.n722 vss 0.069142f
C5009 w_4660_n6791.t32 vss 0.031147f
C5010 w_4660_n6791.t423 vss 0.031147f
C5011 w_4660_n6791.n723 vss 0.07032f
C5012 w_4660_n6791.t384 vss 0.031147f
C5013 w_4660_n6791.t188 vss 0.031147f
C5014 w_4660_n6791.n724 vss 0.069142f
C5015 w_4660_n6791.t182 vss 0.031147f
C5016 w_4660_n6791.t419 vss 0.031147f
C5017 w_4660_n6791.n725 vss 0.07032f
C5018 w_4660_n6791.t320 vss 0.031147f
C5019 w_4660_n6791.t324 vss 0.031147f
C5020 w_4660_n6791.n726 vss 0.069142f
C5021 w_4660_n6791.t132 vss 0.031147f
C5022 w_4660_n6791.t401 vss 0.031147f
C5023 w_4660_n6791.n727 vss 0.07032f
C5024 w_4660_n6791.t246 vss 0.031147f
C5025 w_4660_n6791.t318 vss 0.031147f
C5026 w_4660_n6791.n728 vss 0.069142f
C5027 w_4660_n6791.t437 vss 0.031147f
C5028 w_4660_n6791.t145 vss 0.031147f
C5029 w_4660_n6791.n729 vss 0.07032f
C5030 w_4660_n6791.t375 vss 0.031147f
C5031 w_4660_n6791.t237 vss 0.031147f
C5032 w_4660_n6791.n730 vss 0.069142f
C5033 w_4660_n6791.t27 vss 0.031147f
C5034 w_4660_n6791.t424 vss 0.031147f
C5035 w_4660_n6791.n731 vss 0.07032f
C5036 w_4660_n6791.t360 vss 0.031147f
C5037 w_4660_n6791.t368 vss 0.031147f
C5038 w_4660_n6791.n732 vss 0.069142f
C5039 w_4660_n6791.t116 vss 0.031147f
C5040 w_4660_n6791.t395 vss 0.031147f
C5041 w_4660_n6791.n733 vss 0.07032f
C5042 w_4660_n6791.t287 vss 0.031147f
C5043 w_4660_n6791.t293 vss 0.031147f
C5044 w_4660_n6791.n734 vss 0.069142f
C5045 w_4660_n6791.n735 vss 0.908009f
C5046 w_4660_n6791.n736 vss 0.908009f
C5047 w_4660_n6791.n737 vss 0.908009f
C5048 w_4660_n6791.n738 vss 0.908009f
C5049 w_4660_n6791.n739 vss 0.908009f
C5050 w_4660_n6791.n740 vss 0.908009f
C5051 w_4660_n6791.n741 vss 0.908009f
C5052 w_4660_n6791.n742 vss 0.908009f
C5053 w_4660_n6791.n743 vss 0.908009f
C5054 w_4660_n6791.n744 vss 0.908009f
C5055 w_4660_n6791.n745 vss 0.908009f
C5056 w_4660_n6791.n746 vss 0.908009f
C5057 w_4660_n6791.n747 vss 0.908009f
C5058 w_4660_n6791.n748 vss 0.908009f
C5059 w_4660_n6791.n749 vss 0.908009f
C5060 w_4660_n6791.n750 vss 0.908009f
C5061 w_4660_n6791.n751 vss 0.908009f
C5062 w_4660_n6791.n752 vss 0.908009f
C5063 w_4660_n6791.n753 vss 0.908009f
C5064 w_4660_n6791.n754 vss 0.908009f
C5065 w_4660_n6791.n755 vss 0.908009f
C5066 w_4660_n6791.n756 vss 0.908009f
C5067 w_4660_n6791.n757 vss 0.908009f
C5068 w_4660_n6791.n758 vss 0.908009f
C5069 w_4660_n6791.n759 vss 0.897221f
C5070 w_4660_n6791.n760 vss 0.032221f
C5071 w_4660_n6791.n761 vss 0.013694f
C5072 w_4660_n6791.n762 vss 0.008216f
C5073 w_4660_n6791.n763 vss 0.004315f
C5074 w_4660_n6791.n764 vss 0.008333f
C5075 w_4660_n6791.n765 vss 0.006451f
C5076 w_4660_n6791.n766 vss 0.011278f
C5077 w_4660_n6791.n767 vss 0.00132f
C5078 w_4660_n6791.n768 vss 0.073394f
C5079 w_4660_n6791.n769 vss 0.051465f
C5080 w_4660_n6791.n770 vss 0.009312f
C5081 w_4660_n6791.n771 vss 0.008764f
C5082 w_4660_n6791.n772 vss 0.049227f
C5083 w_4660_n6791.n773 vss 0.008764f
C5084 w_4660_n6791.n774 vss 0.008764f
C5085 w_4660_n6791.n775 vss 0.008764f
C5086 w_4660_n6791.n776 vss 0.056388f
C5087 w_4660_n6791.n777 vss 0.008764f
C5088 w_4660_n6791.n778 vss 0.008764f
C5089 w_4660_n6791.n779 vss 0.008764f
C5090 w_4660_n6791.n780 vss 0.064443f
C5091 w_4660_n6791.n781 vss 0.008764f
C5092 w_4660_n6791.n782 vss 0.008764f
C5093 w_4660_n6791.n783 vss 0.008764f
C5094 w_4660_n6791.n784 vss 0.008764f
C5095 w_4660_n6791.n785 vss 0.008764f
C5096 w_4660_n6791.n786 vss 0.008764f
C5097 w_4660_n6791.n787 vss 0.064443f
C5098 w_4660_n6791.n788 vss 0.042067f
C5099 w_4660_n6791.n789 vss 0.008764f
C5100 w_4660_n6791.n790 vss 0.008764f
C5101 w_4660_n6791.n791 vss 0.054598f
C5102 w_4660_n6791.n792 vss 0.008764f
C5103 w_4660_n6791.n793 vss 0.008764f
C5104 w_4660_n6791.n794 vss 0.008764f
C5105 w_4660_n6791.n795 vss 0.051017f
C5106 w_4660_n6791.n796 vss 0.008764f
C5107 w_4660_n6791.n797 vss 0.008764f
C5108 w_4660_n6791.n798 vss 0.008764f
C5109 w_4660_n6791.n799 vss 0.064443f
C5110 w_4660_n6791.n800 vss 0.059968f
C5111 w_4660_n6791.n801 vss 0.008764f
C5112 w_4660_n6791.n802 vss 0.008764f
C5113 w_4660_n6791.n803 vss 0.036697f
C5114 w_4660_n6791.n804 vss 0.008764f
C5115 w_4660_n6791.n805 vss 0.008764f
C5116 w_4660_n6791.n806 vss 0.008764f
C5117 w_4660_n6791.n807 vss 0.064443f
C5118 w_4660_n6791.n808 vss 0.036697f
C5119 w_4660_n6791.n809 vss 0.008764f
C5120 w_4660_n6791.n810 vss 0.008764f
C5121 w_4660_n6791.n811 vss 0.059968f
C5122 w_4660_n6791.n812 vss 0.008764f
C5123 w_4660_n6791.n813 vss 0.008764f
C5124 w_4660_n6791.n814 vss 0.008764f
C5125 w_4660_n6791.n815 vss 0.045647f
C5126 w_4660_n6791.n816 vss 0.008764f
C5127 w_4660_n6791.n817 vss 0.008764f
C5128 w_4660_n6791.n818 vss 0.008764f
C5129 w_4660_n6791.n819 vss 0.064443f
C5130 w_4660_n6791.n820 vss 0.054598f
C5131 w_4660_n6791.n821 vss 0.008764f
C5132 w_4660_n6791.n822 vss 0.008764f
C5133 w_4660_n6791.n823 vss 0.042067f
C5134 w_4660_n6791.n824 vss 0.008764f
C5135 w_4660_n6791.n825 vss 0.008764f
C5136 w_4660_n6791.n826 vss 0.008764f
C5137 w_4660_n6791.n827 vss 0.063548f
C5138 w_4660_n6791.n828 vss 0.008764f
C5139 w_4660_n6791.n829 vss 0.008764f
C5140 w_4660_n6791.n830 vss 0.008764f
C5141 w_4660_n6791.n831 vss 0.064443f
C5142 w_4660_n6791.n832 vss 0.008764f
C5143 w_4660_n6791.n833 vss 0.008764f
C5144 w_4660_n6791.n834 vss 0.008764f
C5145 w_4660_n6791.n835 vss 0.040277f
C5146 w_4660_n6791.n836 vss 0.008764f
C5147 w_4660_n6791.n837 vss 0.008764f
C5148 w_4660_n6791.n838 vss 0.008764f
C5149 w_4660_n6791.n839 vss 0.064443f
C5150 w_4660_n6791.n840 vss 0.049227f
C5151 w_4660_n6791.n841 vss 0.008764f
C5152 w_4660_n6791.n842 vss 0.008764f
C5153 w_4660_n6791.n843 vss 0.047437f
C5154 w_4660_n6791.n844 vss 0.008764f
C5155 w_4660_n6791.n845 vss 0.008764f
C5156 w_4660_n6791.n846 vss 0.008764f
C5157 w_4660_n6791.n847 vss 0.058178f
C5158 w_4660_n6791.n848 vss 0.008764f
C5159 w_4660_n6791.n849 vss 0.008764f
C5160 w_4660_n6791.n850 vss 0.00633f
C5161 w_4660_n6791.n851 vss 0.064443f
C5162 w_4660_n6791.n852 vss 0.064443f
C5163 w_4660_n6791.n853 vss 0.008764f
C5164 w_4660_n6791.n854 vss 0.006817f
C5165 w_4660_n6791.n855 vss 0.008764f
C5166 w_4660_n6791.n856 vss 0.034907f
C5167 w_4660_n6791.n857 vss 0.008764f
C5168 w_4660_n6791.n858 vss 0.008764f
C5169 w_4660_n6791.n859 vss 0.008764f
C5170 w_4660_n6791.n860 vss 0.064443f
C5171 w_4660_n6791.n861 vss 0.043857f
C5172 w_4660_n6791.n862 vss 0.008764f
C5173 w_4660_n6791.n863 vss 0.008764f
C5174 w_4660_n6791.n864 vss 0.052807f
C5175 w_4660_n6791.n865 vss 0.008764f
C5176 w_4660_n6791.n866 vss 0.008764f
C5177 w_4660_n6791.n867 vss 0.008764f
C5178 w_4660_n6791.n868 vss 0.052807f
C5179 w_4660_n6791.n869 vss 0.008764f
C5180 w_4660_n6791.n870 vss 0.008764f
C5181 w_4660_n6791.n871 vss 0.008764f
C5182 w_4660_n6791.n872 vss 0.064443f
C5183 w_4660_n6791.n873 vss 0.061758f
C5184 w_4660_n6791.n874 vss 0.008764f
C5185 w_4660_n6791.n875 vss 0.008764f
C5186 w_4660_n6791.n876 vss 0.034907f
C5187 w_4660_n6791.n877 vss 0.008764f
C5188 w_4660_n6791.n878 vss 0.008764f
C5189 w_4660_n6791.n879 vss 0.008764f
C5190 w_4660_n6791.n880 vss 0.064443f
C5191 w_4660_n6791.n881 vss 0.038487f
C5192 w_4660_n6791.n882 vss 0.008764f
C5193 w_4660_n6791.n883 vss 0.008764f
C5194 w_4660_n6791.n884 vss 0.058178f
C5195 w_4660_n6791.n885 vss 0.008764f
C5196 w_4660_n6791.n886 vss 0.008764f
C5197 w_4660_n6791.n887 vss 0.008764f
C5198 w_4660_n6791.n888 vss 0.047437f
C5199 w_4660_n6791.n889 vss 0.008764f
C5200 w_4660_n6791.n890 vss 0.008764f
C5201 w_4660_n6791.n891 vss 0.008764f
C5202 w_4660_n6791.n892 vss 0.064443f
C5203 w_4660_n6791.n893 vss 0.056388f
C5204 w_4660_n6791.n894 vss 0.008764f
C5205 w_4660_n6791.n895 vss 0.008764f
C5206 w_4660_n6791.n896 vss 0.040277f
C5207 w_4660_n6791.n897 vss 0.008764f
C5208 w_4660_n6791.n898 vss 0.008764f
C5209 w_4660_n6791.n899 vss 0.008764f
C5210 w_4660_n6791.n900 vss 0.064443f
C5211 w_4660_n6791.n901 vss 0.008764f
C5212 w_4660_n6791.n902 vss 0.008764f
C5213 w_4660_n6791.n903 vss 0.063548f
C5214 w_4660_n6791.n904 vss 0.008764f
C5215 w_4660_n6791.n905 vss 0.008764f
C5216 w_4660_n6791.n906 vss 0.008764f
C5217 w_4660_n6791.n907 vss 0.042067f
C5218 w_4660_n6791.n908 vss 0.008764f
C5219 w_4660_n6791.n909 vss 0.008764f
C5220 w_4660_n6791.n910 vss 0.008764f
C5221 w_4660_n6791.n911 vss 0.064443f
C5222 w_4660_n6791.n912 vss 0.051017f
C5223 w_4660_n6791.n913 vss 0.008764f
C5224 w_4660_n6791.n914 vss 0.008764f
C5225 w_4660_n6791.n915 vss 0.045647f
C5226 w_4660_n6791.n916 vss 0.008764f
C5227 w_4660_n6791.n917 vss 0.008764f
C5228 w_4660_n6791.n918 vss 0.008764f
C5229 w_4660_n6791.n919 vss 0.059968f
C5230 w_4660_n6791.n920 vss 0.008764f
C5231 w_4660_n6791.n921 vss 0.008764f
C5232 w_4660_n6791.n922 vss 0.008764f
C5233 w_4660_n6791.n923 vss 0.064443f
C5234 w_4660_n6791.n924 vss 0.008764f
C5235 w_4660_n6791.n925 vss 0.008764f
C5236 w_4660_n6791.n926 vss 0.008764f
C5237 w_4660_n6791.n927 vss 0.036697f
C5238 w_4660_n6791.n928 vss 0.008764f
C5239 w_4660_n6791.n929 vss 0.008764f
C5240 w_4660_n6791.n930 vss 0.008764f
C5241 w_4660_n6791.n931 vss 0.064443f
C5242 w_4660_n6791.n932 vss 0.045647f
C5243 w_4660_n6791.n933 vss 0.010661f
C5244 w_4660_n6791.n934 vss 0.052229f
C5245 w_4660_n6791.n935 vss 0.063443f
C5246 w_4660_n6791.n936 vss 0.298174f
C5247 w_4660_n6791.n937 vss 0.425158f
C5248 w_4660_n6791.n938 vss 0.01091f
C5249 w_4660_n6791.n939 vss 0.154304f
C5250 w_4660_n6791.n940 vss 0.008764f
C5251 w_4660_n6791.n941 vss 0.010849f
C5252 w_4660_n6791.n942 vss 0.008764f
C5253 w_4660_n6791.n943 vss 0.061865f
C5254 w_4660_n6791.n944 vss 0.022123f
C5255 w_4660_n6791.n945 vss 0.010849f
C5256 w_4660_n6791.n946 vss 0.009022f
C5257 w_4660_n6791.n947 vss 0.061865f
C5258 w_4660_n6791.n948 vss 0.008764f
C5259 w_4660_n6791.n949 vss 0.008764f
C5260 w_4660_n6791.n950 vss 0.061865f
C5261 w_4660_n6791.n951 vss 0.008764f
C5262 w_4660_n6791.n952 vss 0.008764f
C5263 w_4660_n6791.n953 vss 0.009022f
C5264 w_4660_n6791.n954 vss 0.061865f
C5265 w_4660_n6791.n955 vss 0.008764f
C5266 w_4660_n6791.n956 vss 0.008764f
C5267 w_4660_n6791.n957 vss 0.008764f
C5268 w_4660_n6791.n958 vss 0.061865f
C5269 w_4660_n6791.n959 vss 0.008764f
C5270 w_4660_n6791.n960 vss 0.008764f
C5271 w_4660_n6791.n961 vss 0.008764f
C5272 w_4660_n6791.n962 vss 0.008764f
C5273 w_4660_n6791.n963 vss 0.008764f
C5274 w_4660_n6791.n964 vss 0.008764f
C5275 w_4660_n6791.n965 vss 0.061865f
C5276 w_4660_n6791.n966 vss 0.009022f
C5277 w_4660_n6791.n967 vss 0.009022f
C5278 w_4660_n6791.n968 vss 0.009022f
C5279 w_4660_n6791.n969 vss 0.061865f
C5280 w_4660_n6791.n970 vss 0.008764f
C5281 w_4660_n6791.n971 vss 0.008764f
C5282 w_4660_n6791.n972 vss 0.008764f
C5283 w_4660_n6791.n973 vss 0.061865f
C5284 w_4660_n6791.n974 vss 0.009022f
C5285 w_4660_n6791.n975 vss 0.009022f
C5286 w_4660_n6791.n976 vss 0.009022f
C5287 w_4660_n6791.n977 vss 0.061865f
C5288 w_4660_n6791.n978 vss 0.008764f
C5289 w_4660_n6791.n979 vss 0.008764f
C5290 w_4660_n6791.n980 vss 0.008764f
C5291 w_4660_n6791.n981 vss 0.008764f
C5292 w_4660_n6791.n982 vss 0.061865f
C5293 w_4660_n6791.n983 vss 0.009022f
C5294 w_4660_n6791.n984 vss 0.009022f
C5295 w_4660_n6791.n985 vss 0.004389f
C5296 w_4660_n6791.n986 vss 0.008764f
C5297 w_4660_n6791.n987 vss 0.032221f
C5298 w_4660_n6791.n988 vss 0.073394f
C5299 w_4660_n6791.n989 vss 0.001689f
C5300 w_4660_n6791.n990 vss 0.01368f
C5301 w_4660_n6791.n991 vss 0.009312f
C5302 w_4660_n6791.n992 vss 0.008764f
C5303 w_4660_n6791.n993 vss 0.064443f
C5304 w_4660_n6791.n994 vss 0.008764f
C5305 w_4660_n6791.n995 vss 0.032221f
C5306 w_4660_n6791.n996 vss 0.008764f
C5307 w_4660_n6791.n997 vss 0.008764f
C5308 w_4660_n6791.n998 vss 0.008764f
C5309 w_4660_n6791.n999 vss 0.064443f
C5310 w_4660_n6791.n1000 vss 0.008764f
C5311 w_4660_n6791.n1001 vss 0.008764f
C5312 w_4660_n6791.n1002 vss 0.008764f
C5313 w_4660_n6791.n1003 vss 0.064443f
C5314 w_4660_n6791.n1004 vss 0.008764f
C5315 w_4660_n6791.n1005 vss 0.008764f
C5316 w_4660_n6791.n1006 vss 0.032221f
C5317 w_4660_n6791.n1007 vss 0.008764f
C5318 w_4660_n6791.n1008 vss 0.008764f
C5319 w_4660_n6791.n1009 vss 0.008764f
C5320 w_4660_n6791.n1010 vss 0.064443f
C5321 w_4660_n6791.n1011 vss 0.008764f
C5322 w_4660_n6791.n1012 vss 0.032221f
C5323 w_4660_n6791.n1013 vss 0.008764f
C5324 w_4660_n6791.n1014 vss 0.008764f
C5325 w_4660_n6791.n1015 vss 0.008764f
C5326 w_4660_n6791.n1016 vss 0.064443f
C5327 w_4660_n6791.n1017 vss 0.008764f
C5328 w_4660_n6791.n1018 vss 0.032221f
C5329 w_4660_n6791.n1019 vss 0.008764f
C5330 w_4660_n6791.n1020 vss 0.008764f
C5331 w_4660_n6791.n1021 vss 0.008764f
C5332 w_4660_n6791.n1022 vss 0.064443f
C5333 w_4660_n6791.n1023 vss 0.008764f
C5334 w_4660_n6791.n1024 vss 0.036697f
C5335 w_4660_n6791.n1025 vss 0.008764f
C5336 w_4660_n6791.n1026 vss 0.008764f
C5337 w_4660_n6791.n1027 vss 0.008764f
C5338 w_4660_n6791.n1028 vss 0.064443f
C5339 w_4660_n6791.n1029 vss 0.008764f
C5340 w_4660_n6791.n1030 vss 0.032221f
C5341 w_4660_n6791.n1031 vss 0.008764f
C5342 w_4660_n6791.n1032 vss 0.032221f
C5343 w_4660_n6791.n1033 vss 0.008764f
C5344 w_4660_n6791.n1034 vss 0.008764f
C5345 w_4660_n6791.n1035 vss 0.008764f
C5346 w_4660_n6791.n1036 vss 0.064443f
C5347 w_4660_n6791.n1037 vss 0.008764f
C5348 w_4660_n6791.n1038 vss 0.032221f
C5349 w_4660_n6791.n1039 vss 0.008764f
C5350 w_4660_n6791.n1040 vss 0.008764f
C5351 w_4660_n6791.n1041 vss 0.008764f
C5352 w_4660_n6791.n1042 vss 0.064443f
C5353 w_4660_n6791.n1043 vss 0.008764f
C5354 w_4660_n6791.n1044 vss 0.008764f
C5355 w_4660_n6791.n1045 vss 0.008764f
C5356 w_4660_n6791.n1046 vss 0.064443f
C5357 w_4660_n6791.n1047 vss 0.008764f
C5358 w_4660_n6791.n1048 vss 0.040277f
C5359 w_4660_n6791.n1049 vss 0.008764f
C5360 w_4660_n6791.n1050 vss 0.008764f
C5361 w_4660_n6791.n1051 vss 0.008764f
C5362 w_4660_n6791.n1052 vss 0.064443f
C5363 w_4660_n6791.n1053 vss 0.008764f
C5364 w_4660_n6791.n1054 vss 0.032221f
C5365 w_4660_n6791.n1055 vss 0.008764f
C5366 w_4660_n6791.n1056 vss 0.032221f
C5367 w_4660_n6791.n1057 vss 0.008764f
C5368 w_4660_n6791.n1058 vss 0.008764f
C5369 w_4660_n6791.n1059 vss 0.008764f
C5370 w_4660_n6791.n1060 vss 0.064443f
C5371 w_4660_n6791.n1061 vss 0.008764f
C5372 w_4660_n6791.n1062 vss 0.032221f
C5373 w_4660_n6791.n1063 vss 0.008764f
C5374 w_4660_n6791.n1064 vss 0.008764f
C5375 w_4660_n6791.n1065 vss 0.00633f
C5376 w_4660_n6791.n1066 vss 0.064443f
C5377 w_4660_n6791.n1067 vss 0.008764f
C5378 w_4660_n6791.n1068 vss 0.032221f
C5379 w_4660_n6791.n1069 vss 0.006817f
C5380 w_4660_n6791.n1070 vss 0.008764f
C5381 w_4660_n6791.n1071 vss 0.008764f
C5382 w_4660_n6791.n1072 vss 0.064443f
C5383 w_4660_n6791.n1073 vss 0.008764f
C5384 w_4660_n6791.n1074 vss 0.032221f
C5385 w_4660_n6791.n1075 vss 0.008764f
C5386 w_4660_n6791.n1076 vss 0.008764f
C5387 w_4660_n6791.n1077 vss 0.008764f
C5388 w_4660_n6791.n1078 vss 0.064443f
C5389 w_4660_n6791.n1079 vss 0.008764f
C5390 w_4660_n6791.n1080 vss 0.032221f
C5391 w_4660_n6791.n1081 vss 0.008764f
C5392 w_4660_n6791.n1082 vss 0.008764f
C5393 w_4660_n6791.n1083 vss 0.008764f
C5394 w_4660_n6791.n1084 vss 0.064443f
C5395 w_4660_n6791.n1085 vss 0.008764f
C5396 w_4660_n6791.n1086 vss 0.032221f
C5397 w_4660_n6791.n1087 vss 0.008764f
C5398 w_4660_n6791.n1088 vss 0.008764f
C5399 w_4660_n6791.n1089 vss 0.008764f
C5400 w_4660_n6791.n1090 vss 0.064443f
C5401 w_4660_n6791.n1091 vss 0.008764f
C5402 w_4660_n6791.n1092 vss 0.038487f
C5403 w_4660_n6791.n1093 vss 0.008764f
C5404 w_4660_n6791.n1094 vss 0.008764f
C5405 w_4660_n6791.n1095 vss 0.008764f
C5406 w_4660_n6791.n1096 vss 0.064443f
C5407 w_4660_n6791.n1097 vss 0.008764f
C5408 w_4660_n6791.n1098 vss 0.032221f
C5409 w_4660_n6791.n1099 vss 0.008764f
C5410 w_4660_n6791.n1100 vss 0.032221f
C5411 w_4660_n6791.n1101 vss 0.008764f
C5412 w_4660_n6791.n1102 vss 0.008764f
C5413 w_4660_n6791.n1103 vss 0.008764f
C5414 w_4660_n6791.n1104 vss 0.064443f
C5415 w_4660_n6791.n1105 vss 0.008764f
C5416 w_4660_n6791.n1106 vss 0.032221f
C5417 w_4660_n6791.n1107 vss 0.008764f
C5418 w_4660_n6791.n1108 vss 0.008764f
C5419 w_4660_n6791.n1109 vss 0.008764f
C5420 w_4660_n6791.n1110 vss 0.064443f
C5421 w_4660_n6791.n1111 vss 0.008764f
C5422 w_4660_n6791.n1112 vss 0.008764f
C5423 w_4660_n6791.n1113 vss 0.008764f
C5424 w_4660_n6791.n1114 vss 0.064443f
C5425 w_4660_n6791.n1115 vss 0.008764f
C5426 w_4660_n6791.n1116 vss 0.008764f
C5427 w_4660_n6791.n1117 vss 0.008764f
C5428 w_4660_n6791.n1118 vss 0.032221f
C5429 w_4660_n6791.n1119 vss 0.008764f
C5430 w_4660_n6791.n1120 vss 0.008764f
C5431 w_4660_n6791.n1121 vss 0.008764f
C5432 w_4660_n6791.n1122 vss 0.064443f
C5433 w_4660_n6791.n1123 vss 0.008764f
C5434 w_4660_n6791.n1124 vss 0.032221f
C5435 w_4660_n6791.n1125 vss 0.008764f
C5436 w_4660_n6791.n1126 vss 0.008764f
C5437 w_4660_n6791.n1127 vss 0.008764f
C5438 w_4660_n6791.n1128 vss 0.064443f
C5439 w_4660_n6791.n1129 vss 0.008764f
C5440 w_4660_n6791.n1130 vss 0.032221f
C5441 w_4660_n6791.n1131 vss 0.008764f
C5442 w_4660_n6791.n1132 vss 0.008764f
C5443 w_4660_n6791.n1133 vss 0.008764f
C5444 w_4660_n6791.n1134 vss 0.064443f
C5445 w_4660_n6791.n1135 vss 0.008764f
C5446 w_4660_n6791.n1136 vss 0.036697f
C5447 w_4660_n6791.n1137 vss 0.008764f
C5448 w_4660_n6791.n1138 vss 0.008764f
C5449 w_4660_n6791.n1139 vss 0.008764f
C5450 w_4660_n6791.n1140 vss 0.064443f
C5451 w_4660_n6791.n1141 vss 0.008764f
C5452 w_4660_n6791.t286 vss 0.031147f
C5453 w_4660_n6791.t292 vss 0.031147f
C5454 w_4660_n6791.n1142 vss 0.070309f
C5455 w_4660_n6791.t352 vss 0.031147f
C5456 w_4660_n6791.t294 vss 0.031147f
C5457 w_4660_n6791.n1143 vss 0.069153f
C5458 w_4660_n6791.t359 vss 0.031147f
C5459 w_4660_n6791.t365 vss 0.031147f
C5460 w_4660_n6791.n1144 vss 0.070309f
C5461 w_4660_n6791.t379 vss 0.031147f
C5462 w_4660_n6791.t313 vss 0.031147f
C5463 w_4660_n6791.n1145 vss 0.069153f
C5464 w_4660_n6791.t373 vss 0.031147f
C5465 w_4660_n6791.t233 vss 0.031147f
C5466 w_4660_n6791.n1146 vss 0.070309f
C5467 w_4660_n6791.t241 vss 0.031147f
C5468 w_4660_n6791.t351 vss 0.031147f
C5469 w_4660_n6791.n1147 vss 0.069153f
C5470 w_4660_n6791.t244 vss 0.031147f
C5471 w_4660_n6791.t317 vss 0.031147f
C5472 w_4660_n6791.n1148 vss 0.070309f
C5473 w_4660_n6791.t290 vss 0.031147f
C5474 w_4660_n6791.t377 vss 0.031147f
C5475 w_4660_n6791.n1149 vss 0.069153f
C5476 w_4660_n6791.t319 vss 0.031147f
C5477 w_4660_n6791.t323 vss 0.031147f
C5478 w_4660_n6791.n1150 vss 0.070309f
C5479 w_4660_n6791.t310 vss 0.031147f
C5480 w_4660_n6791.t234 vss 0.031147f
C5481 w_4660_n6791.n1151 vss 0.069153f
C5482 w_4660_n6791.t383 vss 0.031147f
C5483 w_4660_n6791.t187 vss 0.031147f
C5484 w_4660_n6791.n1152 vss 0.070309f
C5485 w_4660_n6791.t321 vss 0.031147f
C5486 w_4660_n6791.t255 vss 0.031147f
C5487 w_4660_n6791.n1153 vss 0.069153f
C5488 w_4660_n6791.t189 vss 0.031147f
C5489 w_4660_n6791.t228 vss 0.031147f
C5490 w_4660_n6791.n1154 vss 0.070309f
C5491 w_4660_n6791.t193 vss 0.031147f
C5492 w_4660_n6791.t342 vss 0.031147f
C5493 w_4660_n6791.n1155 vss 0.069153f
C5494 w_4660_n6791.t242 vss 0.031147f
C5495 w_4660_n6791.t297 vss 0.031147f
C5496 w_4660_n6791.n1156 vss 0.070309f
C5497 w_4660_n6791.t278 vss 0.031147f
C5498 w_4660_n6791.t358 vss 0.031147f
C5499 w_4660_n6791.n1157 vss 0.069153f
C5500 w_4660_n6791.t304 vss 0.031147f
C5501 w_4660_n6791.t307 vss 0.031147f
C5502 w_4660_n6791.n1158 vss 0.070309f
C5503 w_4660_n6791.t295 vss 0.031147f
C5504 w_4660_n6791.t218 vss 0.031147f
C5505 w_4660_n6791.n1159 vss 0.069153f
C5506 w_4660_n6791.t381 vss 0.031147f
C5507 w_4660_n6791.t385 vss 0.031147f
C5508 w_4660_n6791.n1160 vss 0.070309f
C5509 w_4660_n6791.t314 vss 0.031147f
C5510 w_4660_n6791.t245 vss 0.031147f
C5511 w_4660_n6791.n1161 vss 0.069153f
C5512 w_4660_n6791.t226 vss 0.031147f
C5513 w_4660_n6791.t235 vss 0.031147f
C5514 w_4660_n6791.n1162 vss 0.070309f
C5515 w_4660_n6791.t325 vss 0.031147f
C5516 w_4660_n6791.t261 vss 0.031147f
C5517 w_4660_n6791.n1163 vss 0.069153f
C5518 w_4660_n6791.t212 vss 0.031147f
C5519 w_4660_n6791.t217 vss 0.031147f
C5520 w_4660_n6791.n1164 vss 0.070309f
C5521 w_4660_n6791.t262 vss 0.031147f
C5522 w_4660_n6791.t194 vss 0.031147f
C5523 w_4660_n6791.n1165 vss 0.069153f
C5524 w_4660_n6791.t301 vss 0.031147f
C5525 w_4660_n6791.t348 vss 0.031147f
C5526 w_4660_n6791.n1166 vss 0.070309f
C5527 w_4660_n6791.t282 vss 0.031147f
C5528 w_4660_n6791.t363 vss 0.031147f
C5529 w_4660_n6791.n1167 vss 0.069153f
C5530 w_4660_n6791.t356 vss 0.031147f
C5531 w_4660_n6791.t361 vss 0.031147f
C5532 w_4660_n6791.n1168 vss 0.070309f
C5533 w_4660_n6791.t298 vss 0.031147f
C5534 w_4660_n6791.t222 vss 0.031147f
C5535 w_4660_n6791.n1169 vss 0.069153f
C5536 w_4660_n6791.t369 vss 0.031147f
C5537 w_4660_n6791.t229 vss 0.031147f
C5538 w_4660_n6791.n1170 vss 0.070309f
C5539 w_4660_n6791.t366 vss 0.031147f
C5540 w_4660_n6791.t249 vss 0.031147f
C5541 w_4660_n6791.n1171 vss 0.069153f
C5542 w_4660_n6791.t267 vss 0.031147f
C5543 w_4660_n6791.t275 vss 0.031147f
C5544 w_4660_n6791.n1172 vss 0.070309f
C5545 w_4660_n6791.t198 vss 0.031147f
C5546 w_4660_n6791.t331 vss 0.031147f
C5547 w_4660_n6791.n1173 vss 0.069153f
C5548 w_4660_n6791.t279 vss 0.031147f
C5549 w_4660_n6791.t284 vss 0.031147f
C5550 w_4660_n6791.n1174 vss 0.070309f
C5551 w_4660_n6791.t265 vss 0.031147f
C5552 w_4660_n6791.t199 vss 0.031147f
C5553 w_4660_n6791.n1175 vss 0.069153f
C5554 w_4660_n6791.t288 vss 0.031147f
C5555 w_4660_n6791.t204 vss 0.031147f
C5556 w_4660_n6791.n1176 vss 0.070309f
C5557 w_4660_n6791.t334 vss 0.031147f
C5558 w_4660_n6791.t372 vss 0.031147f
C5559 w_4660_n6791.n1177 vss 0.069153f
C5560 w_4660_n6791.t206 vss 0.031147f
C5561 w_4660_n6791.t209 vss 0.031147f
C5562 w_4660_n6791.n1178 vss 0.070309f
C5563 w_4660_n6791.t305 vss 0.031147f
C5564 w_4660_n6791.t225 vss 0.031147f
C5565 w_4660_n6791.n1179 vss 0.069153f
C5566 w_4660_n6791.t213 vss 0.031147f
C5567 w_4660_n6791.t200 vss 0.031147f
C5568 w_4660_n6791.n1180 vss 0.070309f
C5569 w_4660_n6791.t374 vss 0.031147f
C5570 w_4660_n6791.t376 vss 0.031147f
C5571 w_4660_n6791.n1181 vss 0.069153f
C5572 w_4660_n6791.t259 vss 0.031147f
C5573 w_4660_n6791.t327 vss 0.031147f
C5574 w_4660_n6791.n1182 vss 0.070309f
C5575 w_4660_n6791.t253 vss 0.031147f
C5576 w_4660_n6791.t336 vss 0.031147f
C5577 w_4660_n6791.n1183 vss 0.069153f
C5578 w_4660_n6791.t333 vss 0.031147f
C5579 w_4660_n6791.t337 vss 0.031147f
C5580 w_4660_n6791.n1184 vss 0.070309f
C5581 w_4660_n6791.t271 vss 0.031147f
C5582 w_4660_n6791.t202 vss 0.031147f
C5583 w_4660_n6791.n1185 vss 0.069153f
C5584 w_4660_n6791.t343 vss 0.031147f
C5585 w_4660_n6791.t195 vss 0.031147f
C5586 w_4660_n6791.n1186 vss 0.070309f
C5587 w_4660_n6791.t338 vss 0.031147f
C5588 w_4660_n6791.t211 vss 0.031147f
C5589 w_4660_n6791.n1187 vss 0.069153f
C5590 w_4660_n6791.t268 vss 0.031147f
C5591 w_4660_n6791.t251 vss 0.031147f
C5592 w_4660_n6791.n1188 vss 0.070309f
C5593 w_4660_n6791.t308 vss 0.031147f
C5594 w_4660_n6791.t311 vss 0.031147f
C5595 w_4660_n6791.n1189 vss 0.069153f
C5596 w_4660_n6791.t254 vss 0.121325f
C5597 w_4660_n6791.t239 vss 0.120265f
C5598 w_4660_n6791.n1190 vss 0.897222f
C5599 w_4660_n6791.n1191 vss 0.90801f
C5600 w_4660_n6791.n1192 vss 0.90801f
C5601 w_4660_n6791.n1193 vss 0.90801f
C5602 w_4660_n6791.n1194 vss 0.90801f
C5603 w_4660_n6791.n1195 vss 0.90801f
C5604 w_4660_n6791.n1196 vss 0.90801f
C5605 w_4660_n6791.n1197 vss 0.90801f
C5606 w_4660_n6791.n1198 vss 0.90801f
C5607 w_4660_n6791.n1199 vss 0.90801f
C5608 w_4660_n6791.n1200 vss 0.90801f
C5609 w_4660_n6791.n1201 vss 0.90801f
C5610 w_4660_n6791.n1202 vss 0.90801f
C5611 w_4660_n6791.n1203 vss 0.90801f
C5612 w_4660_n6791.n1204 vss 0.90801f
C5613 w_4660_n6791.n1205 vss 0.90801f
C5614 w_4660_n6791.n1206 vss 0.90801f
C5615 w_4660_n6791.n1207 vss 0.90801f
C5616 w_4660_n6791.n1208 vss 0.90801f
C5617 w_4660_n6791.n1209 vss 0.90801f
C5618 w_4660_n6791.n1210 vss 0.90801f
C5619 w_4660_n6791.n1211 vss 0.90801f
C5620 w_4660_n6791.n1212 vss 0.90801f
C5621 w_4660_n6791.n1213 vss 0.90801f
C5622 w_4660_n6791.n1214 vss 0.90801f
C5623 w_4660_n6791.n1215 vss 0.032221f
C5624 w_4660_n6791.n1216 vss 0.052229f
C5625 w_4660_n6791.n1217 vss 0.032221f
C5626 w_4660_n6791.n1218 vss 0.008764f
C5627 w_4660_n6791.n1219 vss 0.008764f
C5628 w_4660_n6791.n1220 vss 0.010661f
C5629 w_4660_n6791.n1221 vss 0.045647f
C5630 w_4660_n6791.n1222 vss 0.010661f
C5631 w_4660_n6791.n1223 vss 0.008764f
C5632 w_4660_n6791.n1224 vss 0.008764f
C5633 w_4660_n6791.n1225 vss 0.008764f
C5634 w_4660_n6791.n1226 vss 0.059968f
C5635 w_4660_n6791.n1227 vss 0.008764f
C5636 w_4660_n6791.n1228 vss 0.008764f
C5637 w_4660_n6791.n1229 vss 0.008764f
C5638 w_4660_n6791.n1230 vss 0.064443f
C5639 w_4660_n6791.n1231 vss 0.008764f
C5640 w_4660_n6791.n1232 vss 0.008764f
C5641 w_4660_n6791.n1233 vss 0.008764f
C5642 w_4660_n6791.n1234 vss 0.036697f
C5643 w_4660_n6791.n1235 vss 0.008764f
C5644 w_4660_n6791.n1236 vss 0.008764f
C5645 w_4660_n6791.n1237 vss 0.059968f
C5646 w_4660_n6791.n1238 vss 0.008764f
C5647 w_4660_n6791.n1239 vss 0.008764f
C5648 w_4660_n6791.n1240 vss 0.008764f
C5649 w_4660_n6791.n1241 vss 0.045647f
C5650 w_4660_n6791.n1242 vss 0.008764f
C5651 w_4660_n6791.n1243 vss 0.008764f
C5652 w_4660_n6791.n1244 vss 0.051017f
C5653 w_4660_n6791.n1245 vss 0.008764f
C5654 w_4660_n6791.n1246 vss 0.008764f
C5655 w_4660_n6791.n1247 vss 0.008764f
C5656 w_4660_n6791.n1248 vss 0.054598f
C5657 w_4660_n6791.n1249 vss 0.008764f
C5658 w_4660_n6791.n1250 vss 0.008764f
C5659 w_4660_n6791.n1251 vss 0.042067f
C5660 w_4660_n6791.n1252 vss 0.008764f
C5661 w_4660_n6791.n1253 vss 0.008764f
C5662 w_4660_n6791.n1254 vss 0.008764f
C5663 w_4660_n6791.n1255 vss 0.063548f
C5664 w_4660_n6791.n1256 vss 0.008764f
C5665 w_4660_n6791.n1257 vss 0.008764f
C5666 w_4660_n6791.n1258 vss 0.008764f
C5667 w_4660_n6791.n1259 vss 0.064443f
C5668 w_4660_n6791.n1260 vss 0.008764f
C5669 w_4660_n6791.n1261 vss 0.008764f
C5670 w_4660_n6791.n1262 vss 0.008764f
C5671 w_4660_n6791.n1263 vss 0.040277f
C5672 w_4660_n6791.n1264 vss 0.008764f
C5673 w_4660_n6791.n1265 vss 0.008764f
C5674 w_4660_n6791.n1266 vss 0.056388f
C5675 w_4660_n6791.n1267 vss 0.008764f
C5676 w_4660_n6791.n1268 vss 0.008764f
C5677 w_4660_n6791.n1269 vss 0.008764f
C5678 w_4660_n6791.n1270 vss 0.049227f
C5679 w_4660_n6791.n1271 vss 0.008764f
C5680 w_4660_n6791.n1272 vss 0.008764f
C5681 w_4660_n6791.n1273 vss 0.047437f
C5682 w_4660_n6791.n1274 vss 0.008764f
C5683 w_4660_n6791.n1275 vss 0.008764f
C5684 w_4660_n6791.n1276 vss 0.008764f
C5685 w_4660_n6791.n1277 vss 0.008764f
C5686 w_4660_n6791.n1278 vss 0.058178f
C5687 w_4660_n6791.n1279 vss 0.008764f
C5688 w_4660_n6791.n1280 vss 0.008764f
C5689 w_4660_n6791.n1281 vss 0.008764f
C5690 w_4660_n6791.n1282 vss 0.064443f
C5691 w_4660_n6791.n1283 vss 0.008764f
C5692 w_4660_n6791.n1284 vss 0.008764f
C5693 w_4660_n6791.n1285 vss 0.008764f
C5694 w_4660_n6791.n1286 vss 0.034907f
C5695 w_4660_n6791.n1287 vss 0.008764f
C5696 w_4660_n6791.n1288 vss 0.008764f
C5697 w_4660_n6791.n1289 vss 0.061758f
C5698 w_4660_n6791.n1290 vss 0.008764f
C5699 w_4660_n6791.n1291 vss 0.008764f
C5700 w_4660_n6791.n1292 vss 0.008764f
C5701 w_4660_n6791.n1293 vss 0.043857f
C5702 w_4660_n6791.n1294 vss 0.008764f
C5703 w_4660_n6791.n1295 vss 0.008764f
C5704 w_4660_n6791.n1296 vss 0.052807f
C5705 w_4660_n6791.n1297 vss 0.008764f
C5706 w_4660_n6791.n1298 vss 0.008764f
C5707 w_4660_n6791.n1299 vss 0.008764f
C5708 w_4660_n6791.n1300 vss 0.052807f
C5709 w_4660_n6791.n1301 vss 0.008764f
C5710 w_4660_n6791.n1302 vss 0.008764f
C5711 w_4660_n6791.n1303 vss 0.043857f
C5712 w_4660_n6791.n1304 vss 0.008764f
C5713 w_4660_n6791.n1305 vss 0.008764f
C5714 w_4660_n6791.n1306 vss 0.008764f
C5715 w_4660_n6791.n1307 vss 0.061758f
C5716 w_4660_n6791.n1308 vss 0.008764f
C5717 w_4660_n6791.n1309 vss 0.006817f
C5718 w_4660_n6791.n1310 vss 0.008764f
C5719 w_4660_n6791.n1311 vss 0.034907f
C5720 w_4660_n6791.n1312 vss 0.008764f
C5721 w_4660_n6791.n1313 vss 0.006817f
C5722 w_4660_n6791.n1314 vss 0.004382f
C5723 w_4660_n6791.n1315 vss 0.00633f
C5724 w_4660_n6791.n1316 vss 0.064443f
C5725 w_4660_n6791.n1317 vss 0.00633f
C5726 w_4660_n6791.n1318 vss 0.008764f
C5727 w_4660_n6791.n1319 vss 0.038487f
C5728 w_4660_n6791.n1320 vss 0.008764f
C5729 w_4660_n6791.n1321 vss 0.008764f
C5730 w_4660_n6791.n1322 vss 0.058178f
C5731 w_4660_n6791.n1323 vss 0.008764f
C5732 w_4660_n6791.n1324 vss 0.008764f
C5733 w_4660_n6791.n1325 vss 0.008764f
C5734 w_4660_n6791.n1326 vss 0.047437f
C5735 w_4660_n6791.n1327 vss 0.008764f
C5736 w_4660_n6791.n1328 vss 0.008764f
C5737 w_4660_n6791.n1329 vss 0.049227f
C5738 w_4660_n6791.n1330 vss 0.008764f
C5739 w_4660_n6791.n1331 vss 0.008764f
C5740 w_4660_n6791.n1332 vss 0.008764f
C5741 w_4660_n6791.n1333 vss 0.008764f
C5742 w_4660_n6791.n1334 vss 0.056388f
C5743 w_4660_n6791.n1335 vss 0.008764f
C5744 w_4660_n6791.n1336 vss 0.008764f
C5745 w_4660_n6791.n1337 vss 0.008764f
C5746 w_4660_n6791.n1338 vss 0.064443f
C5747 w_4660_n6791.n1339 vss 0.008764f
C5748 w_4660_n6791.n1340 vss 0.008764f
C5749 w_4660_n6791.n1341 vss 0.008764f
C5750 w_4660_n6791.n1342 vss 0.008764f
C5751 w_4660_n6791.n1343 vss 0.008764f
C5752 w_4660_n6791.n1344 vss 0.063548f
C5753 w_4660_n6791.n1345 vss 0.008764f
C5754 w_4660_n6791.n1346 vss 0.008764f
C5755 w_4660_n6791.n1347 vss 0.008764f
C5756 w_4660_n6791.n1348 vss 0.042067f
C5757 w_4660_n6791.n1349 vss 0.008764f
C5758 w_4660_n6791.n1350 vss 0.008764f
C5759 w_4660_n6791.n1351 vss 0.054598f
C5760 w_4660_n6791.n1352 vss 0.008764f
C5761 w_4660_n6791.n1353 vss 0.008764f
C5762 w_4660_n6791.n1354 vss 0.008764f
C5763 w_4660_n6791.n1355 vss 0.051017f
C5764 w_4660_n6791.n1356 vss 0.008764f
C5765 w_4660_n6791.n1357 vss 0.008764f
C5766 w_4660_n6791.n1358 vss 0.045647f
C5767 w_4660_n6791.n1359 vss 0.008764f
C5768 w_4660_n6791.n1360 vss 0.008764f
C5769 w_4660_n6791.n1361 vss 0.008764f
C5770 w_4660_n6791.n1362 vss 0.008764f
C5771 w_4660_n6791.n1363 vss 0.059968f
C5772 w_4660_n6791.n1364 vss 0.008764f
C5773 w_4660_n6791.n1365 vss 0.008764f
C5774 w_4660_n6791.n1366 vss 0.008764f
C5775 w_4660_n6791.n1367 vss 0.064443f
C5776 w_4660_n6791.n1368 vss 0.008764f
C5777 w_4660_n6791.n1369 vss 0.008764f
C5778 w_4660_n6791.n1370 vss 0.008764f
C5779 w_4660_n6791.n1371 vss 0.036697f
C5780 w_4660_n6791.n1372 vss 0.008764f
C5781 w_4660_n6791.n1373 vss 0.008764f
C5782 w_4660_n6791.n1374 vss 0.059968f
C5783 w_4660_n6791.n1375 vss 0.008764f
C5784 w_4660_n6791.n1376 vss 0.008764f
C5785 w_4660_n6791.n1377 vss 0.008764f
C5786 w_4660_n6791.n1378 vss 0.045647f
C5787 w_4660_n6791.n1379 vss 0.008764f
C5788 w_4660_n6791.n1380 vss 0.008764f
C5789 w_4660_n6791.n1381 vss 0.051017f
C5790 w_4660_n6791.n1382 vss 0.008764f
C5791 w_4660_n6791.n1383 vss 0.008764f
C5792 w_4660_n6791.n1384 vss 0.008764f
C5793 w_4660_n6791.n1385 vss 0.054598f
C5794 w_4660_n6791.n1386 vss 0.008764f
C5795 w_4660_n6791.n1387 vss 0.008764f
C5796 w_4660_n6791.n1388 vss 0.042067f
C5797 w_4660_n6791.n1389 vss 0.008764f
C5798 w_4660_n6791.n1390 vss 0.008764f
C5799 w_4660_n6791.n1391 vss 0.008764f
C5800 w_4660_n6791.n1392 vss 0.008764f
C5801 w_4660_n6791.n1393 vss 0.063548f
C5802 w_4660_n6791.n1394 vss 0.008764f
C5803 w_4660_n6791.n1395 vss 0.008764f
C5804 w_4660_n6791.n1396 vss 0.008764f
C5805 w_4660_n6791.n1397 vss 0.064443f
C5806 w_4660_n6791.n1398 vss 0.008764f
C5807 w_4660_n6791.n1399 vss 0.008764f
C5808 w_4660_n6791.n1400 vss 0.008764f
C5809 w_4660_n6791.n1401 vss 0.040277f
C5810 w_4660_n6791.n1402 vss 0.008764f
C5811 w_4660_n6791.n1403 vss 0.008764f
C5812 w_4660_n6791.n1404 vss 0.056388f
C5813 w_4660_n6791.n1405 vss 0.008764f
C5814 w_4660_n6791.n1406 vss 0.008764f
C5815 w_4660_n6791.n1407 vss 0.008764f
C5816 w_4660_n6791.n1408 vss 0.049227f
C5817 w_4660_n6791.n1409 vss 0.008764f
C5818 w_4660_n6791.n1410 vss 0.009312f
C5819 w_4660_n6791.n1411 vss 0.051465f
C5820 w_4660_n6791.n1412 vss 0.008216f
C5821 w_4660_n6791.n1413 vss 0.008342f
C5822 w_4660_n6791.n1414 vss 0.008832f
C5823 w_4660_n6791.n1415 vss 0.044681f
C5824 w_4660_n6791.n1416 vss 0.010849f
C5825 w_4660_n6791.n1417 vss 0.028693f
C5826 w_4660_n6791.n1418 vss 0.010849f
C5827 w_4660_n6791.n1419 vss 0.03351f
C5828 w_4660_n6791.n1420 vss 0.005403f
C5829 w_4660_n6791.n1421 vss 0.189917f
C5830 w_4660_n6791.n1422 vss 0.005073f
C5831 w_4660_n6791.n1423 vss 0.009022f
C5832 w_4660_n6791.n1424 vss 0.061865f
C5833 w_4660_n6791.n1425 vss 0.008764f
C5834 w_4660_n6791.n1426 vss 0.008764f
C5835 w_4660_n6791.n1427 vss 0.008764f
C5836 w_4660_n6791.n1428 vss 0.061865f
C5837 w_4660_n6791.n1429 vss 0.009022f
C5838 w_4660_n6791.n1430 vss 0.009022f
C5839 w_4660_n6791.n1431 vss 0.009022f
C5840 w_4660_n6791.n1432 vss 0.061865f
C5841 w_4660_n6791.n1433 vss 0.008764f
C5842 w_4660_n6791.n1434 vss 0.008764f
C5843 w_4660_n6791.n1435 vss 0.008764f
C5844 w_4660_n6791.n1436 vss 0.061865f
C5845 w_4660_n6791.n1437 vss 0.009022f
C5846 w_4660_n6791.n1438 vss 0.009022f
C5847 w_4660_n6791.n1439 vss 0.009022f
C5848 w_4660_n6791.n1440 vss 0.061865f
C5849 w_4660_n6791.n1441 vss 0.008764f
C5850 w_4660_n6791.n1442 vss 0.008764f
C5851 w_4660_n6791.n1443 vss 0.008764f
C5852 w_4660_n6791.n1444 vss 0.061865f
C5853 w_4660_n6791.n1445 vss 0.009022f
C5854 w_4660_n6791.n1446 vss 0.005198f
C5855 w_4660_n6791.n1447 vss 0.004507f
C5856 w_4660_n6791.n1448 vss 0.008331f
C5857 w_4660_n6791.n1449 vss 0.061865f
C5858 w_4660_n6791.n1450 vss 0.008764f
C5859 w_4660_n6791.n1451 vss 0.008764f
C5860 w_4660_n6791.n1452 vss 0.008764f
C5861 w_4660_n6791.n1453 vss 0.061865f
C5862 w_4660_n6791.n1454 vss 0.009022f
C5863 w_4660_n6791.n1455 vss 0.009022f
C5864 w_4660_n6791.n1456 vss 0.009022f
C5865 w_4660_n6791.n1457 vss 0.061865f
C5866 w_4660_n6791.n1458 vss 0.008764f
C5867 w_4660_n6791.n1459 vss 0.008764f
C5868 w_4660_n6791.n1460 vss 0.008764f
C5869 w_4660_n6791.n1461 vss 0.008764f
C5870 w_4660_n6791.n1462 vss 0.061865f
C5871 w_4660_n6791.n1463 vss 0.009022f
C5872 w_4660_n6791.n1464 vss 0.009022f
C5873 w_4660_n6791.n1465 vss 0.009022f
C5874 w_4660_n6791.n1466 vss 0.009022f
C5875 w_4660_n6791.n1467 vss 0.061865f
C5876 w_4660_n6791.n1468 vss 0.008764f
C5877 w_4660_n6791.n1469 vss 0.008764f
C5878 w_4660_n6791.n1470 vss 0.011051f
C5879 w_4660_n6791.n1471 vss 0.030484f
C5880 w_4660_n6791.n1472 vss 0.011051f
C5881 w_4660_n6791.n1473 vss 0.059288f
C5882 w_4660_n6791.n1474 vss 0.011051f
C5883 w_4660_n6791.n1475 vss 0.05336f
C5884 w_4660_n6791.n1476 vss 0.011051f
C5885 w_4660_n6791.n1477 vss 0.008764f
C5886 w_4660_n6791.n1478 vss 0.008764f
C5887 w_4660_n6791.n1479 vss 0.008764f
C5888 w_4660_n6791.n1480 vss 0.061865f
C5889 w_4660_n6791.n1481 vss 0.009022f
C5890 w_4660_n6791.n1482 vss 0.008764f
C5891 w_4660_n6791.n1483 vss 0.008764f
C5892 w_4660_n6791.n1484 vss 0.061865f
C5893 w_4660_n6791.n1485 vss 0.008764f
C5894 w_4660_n6791.n1486 vss 0.008764f
C5895 w_4660_n6791.n1487 vss 0.008764f
C5896 w_4660_n6791.n1488 vss 0.061865f
C5897 w_4660_n6791.n1489 vss 0.009022f
C5898 w_4660_n6791.n1490 vss 0.008764f
C5899 w_4660_n6791.n1491 vss 0.008764f
C5900 w_4660_n6791.n1492 vss 0.061865f
C5901 w_4660_n6791.n1493 vss 0.008764f
C5902 w_4660_n6791.n1494 vss 0.008764f
C5903 w_4660_n6791.n1495 vss 0.008764f
C5904 w_4660_n6791.n1496 vss 0.009022f
C5905 w_4660_n6791.n1497 vss 0.061865f
C5906 w_4660_n6791.n1498 vss 0.008764f
C5907 w_4660_n6791.n1499 vss 0.008764f
C5908 w_4660_n6791.n1500 vss 0.008764f
C5909 w_4660_n6791.n1501 vss 0.061865f
C5910 w_4660_n6791.n1502 vss 0.009022f
C5911 w_4660_n6791.n1503 vss 0.009022f
C5912 w_4660_n6791.n1504 vss 0.009022f
C5913 w_4660_n6791.n1505 vss 0.061865f
C5914 w_4660_n6791.n1506 vss 0.008764f
C5915 w_4660_n6791.n1507 vss 0.008764f
C5916 w_4660_n6791.n1508 vss 0.008764f
C5917 w_4660_n6791.n1509 vss 0.061865f
C5918 w_4660_n6791.n1510 vss 0.009022f
C5919 w_4660_n6791.n1511 vss 0.009022f
C5920 w_4660_n6791.n1512 vss 0.009022f
C5921 w_4660_n6791.n1513 vss 0.061865f
C5922 w_4660_n6791.n1514 vss 0.008764f
C5923 w_4660_n6791.n1515 vss 0.008764f
C5924 w_4660_n6791.n1516 vss 0.008764f
C5925 w_4660_n6791.n1517 vss 0.061865f
C5926 w_4660_n6791.n1518 vss 0.007454f
C5927 w_4660_n6791.n1519 vss 0.189961f
C5928 w_4660_n6791.n1520 vss 0.425158f
C5929 w_4660_n6791.n1521 vss 0.008764f
C5930 w_4660_n6791.n1522 vss 0.011345f
C5931 w_4660_n6791.n1523 vss 0.032221f
C5932 w_4660_n6791.n1524 vss 0.008764f
C5933 w_4660_n6791.n1525 vss 0.008764f
C5934 w_4660_n6791.n1526 vss 0.056388f
C5935 w_4660_n6791.n1527 vss 0.008764f
C5936 w_4660_n6791.n1528 vss 0.032221f
C5937 w_4660_n6791.n1529 vss 0.008764f
C5938 w_4660_n6791.n1530 vss 0.008764f
C5939 w_4660_n6791.n1531 vss 0.064443f
C5940 w_4660_n6791.n1532 vss 0.008764f
C5941 w_4660_n6791.n1533 vss 0.008764f
C5942 w_4660_n6791.n1534 vss 0.008764f
C5943 w_4660_n6791.n1535 vss 0.008764f
C5944 w_4660_n6791.n1536 vss 0.008764f
C5945 w_4660_n6791.n1537 vss 0.008764f
C5946 w_4660_n6791.n1538 vss 0.064443f
C5947 w_4660_n6791.n1539 vss 0.008764f
C5948 w_4660_n6791.n1540 vss 0.008764f
C5949 w_4660_n6791.n1541 vss 0.008764f
C5950 w_4660_n6791.n1542 vss 0.032221f
C5951 w_4660_n6791.n1543 vss 0.008764f
C5952 w_4660_n6791.n1544 vss 0.008764f
C5953 w_4660_n6791.n1545 vss 0.008764f
C5954 w_4660_n6791.n1546 vss 0.051017f
C5955 w_4660_n6791.n1547 vss 0.008764f
C5956 w_4660_n6791.n1548 vss 0.032221f
C5957 w_4660_n6791.n1549 vss 0.008764f
C5958 w_4660_n6791.n1550 vss 0.008764f
C5959 w_4660_n6791.n1551 vss 0.064443f
C5960 w_4660_n6791.n1552 vss 0.008764f
C5961 w_4660_n6791.n1553 vss 0.008764f
C5962 w_4660_n6791.n1554 vss 0.008764f
C5963 w_4660_n6791.n1555 vss 0.008764f
C5964 w_4660_n6791.n1556 vss 0.032221f
C5965 w_4660_n6791.n1557 vss 0.008764f
C5966 w_4660_n6791.n1558 vss 0.008764f
C5967 w_4660_n6791.n1559 vss 0.008764f
C5968 w_4660_n6791.n1560 vss 0.064443f
C5969 w_4660_n6791.n1561 vss 0.008764f
C5970 w_4660_n6791.n1562 vss 0.008764f
C5971 w_4660_n6791.n1563 vss 0.008764f
C5972 w_4660_n6791.n1564 vss 0.032221f
C5973 w_4660_n6791.n1565 vss 0.008764f
C5974 w_4660_n6791.n1566 vss 0.008764f
C5975 w_4660_n6791.n1567 vss 0.008764f
C5976 w_4660_n6791.n1568 vss 0.008764f
C5977 w_4660_n6791.n1569 vss 0.045647f
C5978 w_4660_n6791.n1570 vss 0.008764f
C5979 w_4660_n6791.n1571 vss 0.032221f
C5980 w_4660_n6791.n1572 vss 0.008764f
C5981 w_4660_n6791.n1573 vss 0.008764f
C5982 w_4660_n6791.n1574 vss 0.064443f
C5983 w_4660_n6791.n1575 vss 0.008764f
C5984 w_4660_n6791.n1576 vss 0.008764f
C5985 w_4660_n6791.n1577 vss 0.008764f
C5986 w_4660_n6791.n1578 vss 0.008764f
C5987 w_4660_n6791.n1579 vss 0.032221f
C5988 w_4660_n6791.n1580 vss 0.008764f
C5989 w_4660_n6791.n1581 vss 0.008764f
C5990 w_4660_n6791.n1582 vss 0.008764f
C5991 w_4660_n6791.n1583 vss 0.008764f
C5992 w_4660_n6791.n1584 vss 0.008764f
C5993 w_4660_n6791.n1585 vss 0.008764f
C5994 w_4660_n6791.n1586 vss 0.064443f
C5995 w_4660_n6791.n1587 vss 0.008764f
C5996 w_4660_n6791.n1588 vss 0.008764f
C5997 w_4660_n6791.n1589 vss 0.008764f
C5998 w_4660_n6791.n1590 vss 0.008764f
C5999 w_4660_n6791.n1591 vss 0.040277f
C6000 w_4660_n6791.n1592 vss 0.008764f
C6001 w_4660_n6791.n1593 vss 0.032221f
C6002 w_4660_n6791.n1594 vss 0.008764f
C6003 w_4660_n6791.n1595 vss 0.008764f
C6004 w_4660_n6791.n1596 vss 0.064443f
C6005 w_4660_n6791.n1597 vss 0.008764f
C6006 w_4660_n6791.n1598 vss 0.008764f
C6007 w_4660_n6791.n1599 vss 0.008764f
C6008 w_4660_n6791.n1600 vss 0.032221f
C6009 w_4660_n6791.n1601 vss 0.008764f
C6010 w_4660_n6791.n1602 vss 0.008764f
C6011 w_4660_n6791.n1603 vss 0.008764f
C6012 w_4660_n6791.n1604 vss 0.058178f
C6013 w_4660_n6791.n1605 vss 0.004382f
C6014 w_4660_n6791.n1606 vss 0.00633f
C6015 w_4660_n6791.t140 vss 0.031147f
C6016 w_4660_n6791.t161 vss 0.031147f
C6017 w_4660_n6791.n1607 vss 0.07032f
C6018 w_4660_n6791.t100 vss 0.031147f
C6019 w_4660_n6791.t464 vss 0.031147f
C6020 w_4660_n6791.n1608 vss 0.069153f
C6021 w_4660_n6791.t430 vss 0.031147f
C6022 w_4660_n6791.t156 vss 0.031147f
C6023 w_4660_n6791.n1609 vss 0.07032f
C6024 w_4660_n6791.t68 vss 0.031147f
C6025 w_4660_n6791.t478 vss 0.031147f
C6026 w_4660_n6791.n1610 vss 0.069153f
C6027 w_4660_n6791.t87 vss 0.031147f
C6028 w_4660_n6791.t393 vss 0.031147f
C6029 w_4660_n6791.n1611 vss 0.07032f
C6030 w_4660_n6791.t117 vss 0.031147f
C6031 w_4660_n6791.t38 vss 0.031147f
C6032 w_4660_n6791.n1612 vss 0.069153f
C6033 w_4660_n6791.t475 vss 0.031147f
C6034 w_4660_n6791.t128 vss 0.031147f
C6035 w_4660_n6791.n1613 vss 0.07032f
C6036 w_4660_n6791.t400 vss 0.031147f
C6037 w_4660_n6791.t147 vss 0.031147f
C6038 w_4660_n6791.n1614 vss 0.069153f
C6039 w_4660_n6791.t120 vss 0.031147f
C6040 w_4660_n6791.t31 vss 0.031147f
C6041 w_4660_n6791.n1615 vss 0.07032f
C6042 w_4660_n6791.t48 vss 0.031147f
C6043 w_4660_n6791.t392 vss 0.031147f
C6044 w_4660_n6791.n1616 vss 0.069153f
C6045 w_4660_n6791.t416 vss 0.031147f
C6046 w_4660_n6791.t127 vss 0.031147f
C6047 w_4660_n6791.n1617 vss 0.07032f
C6048 w_4660_n6791.t4 vss 0.031147f
C6049 w_4660_n6791.t71 vss 0.031147f
C6050 w_4660_n6791.n1618 vss 0.069153f
C6051 w_4660_n6791.t418 vss 0.031147f
C6052 w_4660_n6791.t66 vss 0.031147f
C6053 w_4660_n6791.n1619 vss 0.07032f
C6054 w_4660_n6791.t8 vss 0.031147f
C6055 w_4660_n6791.t34 vss 0.031147f
C6056 w_4660_n6791.n1620 vss 0.069153f
C6057 w_4660_n6791.t477 vss 0.031147f
C6058 w_4660_n6791.t479 vss 0.031147f
C6059 w_4660_n6791.n1621 vss 0.07032f
C6060 w_4660_n6791.t426 vss 0.031147f
C6061 w_4660_n6791.t95 vss 0.031147f
C6062 w_4660_n6791.n1622 vss 0.069153f
C6063 w_4660_n6791.t119 vss 0.031147f
C6064 w_4660_n6791.t61 vss 0.031147f
C6065 w_4660_n6791.n1623 vss 0.07032f
C6066 w_4660_n6791.t173 vss 0.031147f
C6067 w_4660_n6791.t101 vss 0.031147f
C6068 w_4660_n6791.n1624 vss 0.069153f
C6069 w_4660_n6791.t397 vss 0.031147f
C6070 w_4660_n6791.t155 vss 0.031147f
C6071 w_4660_n6791.n1625 vss 0.07032f
C6072 w_4660_n6791.t422 vss 0.031147f
C6073 w_4660_n6791.t154 vss 0.031147f
C6074 w_4660_n6791.n1626 vss 0.069153f
C6075 w_4660_n6791.t465 vss 0.031147f
C6076 w_4660_n6791.t413 vss 0.031147f
C6077 w_4660_n6791.n1627 vss 0.07032f
C6078 w_4660_n6791.t26 vss 0.031147f
C6079 w_4660_n6791.t167 vss 0.031147f
C6080 w_4660_n6791.n1628 vss 0.069153f
C6081 w_4660_n6791.t417 vss 0.031147f
C6082 w_4660_n6791.t405 vss 0.031147f
C6083 w_4660_n6791.n1629 vss 0.07032f
C6084 w_4660_n6791.t18 vss 0.031147f
C6085 w_4660_n6791.t396 vss 0.031147f
C6086 w_4660_n6791.n1630 vss 0.069153f
C6087 w_4660_n6791.n1631 vss 0.90734f
C6088 w_4660_n6791.n1632 vss 0.90734f
C6089 w_4660_n6791.n1633 vss 0.90734f
C6090 w_4660_n6791.n1634 vss 0.90734f
C6091 w_4660_n6791.n1635 vss 0.90734f
C6092 w_4660_n6791.n1636 vss 0.90734f
C6093 w_4660_n6791.n1637 vss 0.90734f
C6094 w_4660_n6791.n1638 vss 0.90734f
C6095 w_4660_n6791.n1639 vss 0.90734f
C6096 w_4660_n6791.n1640 vss 0.90734f
C6097 w_4660_n6791.n1641 vss 0.90734f
C6098 w_4660_n6791.t44 vss 0.031147f
C6099 w_4660_n6791.t174 vss 0.031147f
C6100 w_4660_n6791.n1642 vss 0.07032f
C6101 w_4660_n6791.t403 vss 0.031147f
C6102 w_4660_n6791.t164 vss 0.031147f
C6103 w_4660_n6791.n1643 vss 0.069153f
C6104 w_4660_n6791.t49 vss 0.031147f
C6105 w_4660_n6791.t451 vss 0.031147f
C6106 w_4660_n6791.n1644 vss 0.07032f
C6107 w_4660_n6791.t85 vss 0.031147f
C6108 w_4660_n6791.t157 vss 0.031147f
C6109 w_4660_n6791.n1645 vss 0.069153f
C6110 w_4660_n6791.t443 vss 0.031147f
C6111 w_4660_n6791.t90 vss 0.031147f
C6112 w_4660_n6791.n1646 vss 0.07032f
C6113 w_4660_n6791.t169 vss 0.031147f
C6114 w_4660_n6791.t114 vss 0.031147f
C6115 w_4660_n6791.n1647 vss 0.069153f
C6116 w_4660_n6791.t408 vss 0.031147f
C6117 w_4660_n6791.t36 vss 0.031147f
C6118 w_4660_n6791.n1648 vss 0.07032f
C6119 w_4660_n6791.t126 vss 0.031147f
C6120 w_4660_n6791.t150 vss 0.031147f
C6121 w_4660_n6791.n1649 vss 0.069153f
C6122 w_4660_n6791.t407 vss 0.031147f
C6123 w_4660_n6791.t391 vss 0.031147f
C6124 w_4660_n6791.n1650 vss 0.07032f
C6125 w_4660_n6791.t73 vss 0.031147f
C6126 w_4660_n6791.t99 vss 0.031147f
C6127 w_4660_n6791.n1651 vss 0.069153f
C6128 w_4660_n6791.t16 vss 0.031147f
C6129 w_4660_n6791.t441 vss 0.031147f
C6130 w_4660_n6791.n1652 vss 0.07032f
C6131 w_4660_n6791.t453 vss 0.031147f
C6132 w_4660_n6791.t406 vss 0.031147f
C6133 w_4660_n6791.n1653 vss 0.069153f
C6134 w_4660_n6791.t179 vss 0.031147f
C6135 w_4660_n6791.t74 vss 0.031147f
C6136 w_4660_n6791.n1654 vss 0.07032f
C6137 w_4660_n6791.t133 vss 0.031147f
C6138 w_4660_n6791.t54 vss 0.031147f
C6139 w_4660_n6791.n1655 vss 0.069153f
C6140 w_4660_n6791.t176 vss 0.031147f
C6141 w_4660_n6791.t76 vss 0.031147f
C6142 w_4660_n6791.n1656 vss 0.07032f
C6143 w_4660_n6791.t24 vss 0.031147f
C6144 w_4660_n6791.t104 vss 0.031147f
C6145 w_4660_n6791.n1657 vss 0.069153f
C6146 w_4660_n6791.t9 vss 0.031147f
C6147 w_4660_n6791.t428 vss 0.031147f
C6148 w_4660_n6791.n1658 vss 0.07032f
C6149 w_4660_n6791.t438 vss 0.031147f
C6150 w_4660_n6791.t75 vss 0.031147f
C6151 w_4660_n6791.n1659 vss 0.069153f
C6152 w_4660_n6791.t135 vss 0.031147f
C6153 w_4660_n6791.t466 vss 0.031147f
C6154 w_4660_n6791.n1660 vss 0.07032f
C6155 w_4660_n6791.t46 vss 0.031147f
C6156 w_4660_n6791.t177 vss 0.031147f
C6157 w_4660_n6791.n1661 vss 0.069153f
C6158 w_4660_n6791.n1662 vss 0.90734f
C6159 w_4660_n6791.n1663 vss 0.90734f
C6160 w_4660_n6791.n1664 vss 0.90734f
C6161 w_4660_n6791.n1665 vss 0.90734f
C6162 w_4660_n6791.n1666 vss 0.90734f
C6163 w_4660_n6791.n1667 vss 0.90734f
C6164 w_4660_n6791.n1668 vss 0.90734f
C6165 w_4660_n6791.n1669 vss 0.90734f
C6166 w_4660_n6791.n1670 vss 0.90734f
C6167 w_4660_n6791.n1671 vss 0.90734f
C6168 w_4660_n6791.n1672 vss 0.90734f
C6169 w_4660_n6791.n1673 vss 0.032221f
C6170 w_4660_n6791.n1674 vss 0.008764f
C6171 w_4660_n6791.n1675 vss 0.008764f
C6172 w_4660_n6791.n1676 vss 0.064443f
C6173 w_4660_n6791.n1677 vss 0.008764f
C6174 w_4660_n6791.n1678 vss 0.00633f
C6175 w_4660_n6791.n1679 vss 0.008764f
C6176 w_4660_n6791.n1680 vss 0.038487f
C6177 w_4660_n6791.n1681 vss 0.008764f
C6178 w_4660_n6791.n1682 vss 0.008764f
C6179 w_4660_n6791.n1683 vss 0.008764f
C6180 w_4660_n6791.n1684 vss 0.064443f
C6181 w_4660_n6791.n1685 vss 0.047437f
C6182 w_4660_n6791.n1686 vss 0.008764f
C6183 w_4660_n6791.n1687 vss 0.008764f
C6184 w_4660_n6791.n1688 vss 0.049227f
C6185 w_4660_n6791.n1689 vss 0.008764f
C6186 w_4660_n6791.n1690 vss 0.008764f
C6187 w_4660_n6791.n1691 vss 0.008764f
C6188 w_4660_n6791.n1692 vss 0.056388f
C6189 w_4660_n6791.n1693 vss 0.008764f
C6190 w_4660_n6791.n1694 vss 0.008764f
C6191 w_4660_n6791.n1695 vss 0.008764f
C6192 w_4660_n6791.n1696 vss 0.064443f
C6193 w_4660_n6791.n1697 vss 0.008764f
C6194 w_4660_n6791.n1698 vss 0.008764f
C6195 w_4660_n6791.n1699 vss 0.008764f
C6196 w_4660_n6791.n1700 vss 0.008764f
C6197 w_4660_n6791.n1701 vss 0.008764f
C6198 w_4660_n6791.n1702 vss 0.008764f
C6199 w_4660_n6791.n1703 vss 0.064443f
C6200 w_4660_n6791.n1704 vss 0.042067f
C6201 w_4660_n6791.n1705 vss 0.008764f
C6202 w_4660_n6791.n1706 vss 0.008764f
C6203 w_4660_n6791.n1707 vss 0.054598f
C6204 w_4660_n6791.n1708 vss 0.008764f
C6205 w_4660_n6791.n1709 vss 0.008764f
C6206 w_4660_n6791.n1710 vss 0.008764f
C6207 w_4660_n6791.n1711 vss 0.051017f
C6208 w_4660_n6791.n1712 vss 0.008764f
C6209 w_4660_n6791.n1713 vss 0.008764f
C6210 w_4660_n6791.n1714 vss 0.008764f
C6211 w_4660_n6791.n1715 vss 0.064443f
C6212 w_4660_n6791.n1716 vss 0.059968f
C6213 w_4660_n6791.n1717 vss 0.008764f
C6214 w_4660_n6791.n1718 vss 0.008764f
C6215 w_4660_n6791.n1719 vss 0.036697f
C6216 w_4660_n6791.n1720 vss 0.008764f
C6217 w_4660_n6791.n1721 vss 0.008764f
C6218 w_4660_n6791.n1722 vss 0.008764f
C6219 w_4660_n6791.n1723 vss 0.064443f
C6220 w_4660_n6791.n1724 vss 0.036697f
C6221 w_4660_n6791.n1725 vss 0.008764f
C6222 w_4660_n6791.n1726 vss 0.008764f
C6223 w_4660_n6791.n1727 vss 0.059968f
C6224 w_4660_n6791.n1728 vss 0.008764f
C6225 w_4660_n6791.n1729 vss 0.008764f
C6226 w_4660_n6791.n1730 vss 0.008764f
C6227 w_4660_n6791.n1731 vss 0.045647f
C6228 w_4660_n6791.n1732 vss 0.008764f
C6229 w_4660_n6791.n1733 vss 0.008764f
C6230 w_4660_n6791.n1734 vss 0.008764f
C6231 w_4660_n6791.n1735 vss 0.064443f
C6232 w_4660_n6791.n1736 vss 0.054598f
C6233 w_4660_n6791.n1737 vss 0.008764f
C6234 w_4660_n6791.n1738 vss 0.008764f
C6235 w_4660_n6791.n1739 vss 0.042067f
C6236 w_4660_n6791.n1740 vss 0.008764f
C6237 w_4660_n6791.n1741 vss 0.008764f
C6238 w_4660_n6791.n1742 vss 0.008764f
C6239 w_4660_n6791.n1743 vss 0.063548f
C6240 w_4660_n6791.n1744 vss 0.008764f
C6241 w_4660_n6791.n1745 vss 0.008764f
C6242 w_4660_n6791.n1746 vss 0.008764f
C6243 w_4660_n6791.n1747 vss 0.064443f
C6244 w_4660_n6791.n1748 vss 0.008764f
C6245 w_4660_n6791.n1749 vss 0.008764f
C6246 w_4660_n6791.n1750 vss 0.008764f
C6247 w_4660_n6791.n1751 vss 0.040277f
C6248 w_4660_n6791.n1752 vss 0.008764f
C6249 w_4660_n6791.n1753 vss 0.008764f
C6250 w_4660_n6791.n1754 vss 0.008764f
C6251 w_4660_n6791.n1755 vss 0.064443f
C6252 w_4660_n6791.n1756 vss 0.049227f
C6253 w_4660_n6791.n1757 vss 0.011345f
C6254 w_4660_n6791.n1758 vss 0.072327f
C6255 w_4660_n6791.n1759 vss 0.063914f
C6256 w_4660_n6791.n1760 vss 0.298677f
C6257 w_4660_n6791.n1761 vss 0.48173f
C6258 w_4660_n6791.n1762 vss 4.17527f
C6259 w_4660_n6791.n1763 vss 0.48173f
C6260 w_4660_n6791.n1764 vss 0.115121f
C6261 w_4660_n6791.n1765 vss 0.063914f
C6262 w_4660_n6791.n1766 vss 0.008764f
C6263 w_4660_n6791.n1767 vss 0.008764f
C6264 w_4660_n6791.n1768 vss 0.008764f
C6265 w_4660_n6791.n1769 vss 0.032221f
C6266 w_4660_n6791.n1770 vss 0.008764f
C6267 w_4660_n6791.n1771 vss 0.008764f
C6268 w_4660_n6791.n1772 vss 0.008764f
C6269 w_4660_n6791.n1773 vss 0.008764f
C6270 w_4660_n6791.n1774 vss 0.008764f
C6271 w_4660_n6791.n1775 vss 0.008764f
C6272 w_4660_n6791.n1776 vss 0.008764f
C6273 w_4660_n6791.n1777 vss 0.008764f
C6274 w_4660_n6791.n1778 vss 0.008764f
C6275 w_4660_n6791.n1779 vss 0.008764f
C6276 w_4660_n6791.n1780 vss 0.008764f
C6277 w_4660_n6791.n1781 vss 0.042067f
C6278 w_4660_n6791.n1782 vss 0.008764f
C6279 w_4660_n6791.n1783 vss 0.032221f
C6280 w_4660_n6791.n1784 vss 0.008764f
C6281 w_4660_n6791.n1785 vss 0.008764f
C6282 w_4660_n6791.n1786 vss 0.064443f
C6283 w_4660_n6791.n1787 vss 0.008764f
C6284 w_4660_n6791.n1788 vss 0.008764f
C6285 w_4660_n6791.n1789 vss 0.008764f
C6286 w_4660_n6791.n1790 vss 0.008764f
C6287 w_4660_n6791.n1791 vss 0.032221f
C6288 w_4660_n6791.n1792 vss 0.008764f
C6289 w_4660_n6791.n1793 vss 0.008764f
C6290 w_4660_n6791.n1794 vss 0.008764f
C6291 w_4660_n6791.n1795 vss 0.059968f
C6292 w_4660_n6791.n1796 vss 0.008764f
C6293 w_4660_n6791.n1797 vss 0.032221f
C6294 w_4660_n6791.n1798 vss 0.008764f
C6295 w_4660_n6791.n1799 vss 0.008764f
C6296 w_4660_n6791.n1800 vss 0.064443f
C6297 w_4660_n6791.n1801 vss 0.008764f
C6298 w_4660_n6791.n1802 vss 0.008764f
C6299 w_4660_n6791.n1803 vss 0.008764f
C6300 w_4660_n6791.n1804 vss 0.008764f
C6301 w_4660_n6791.n1805 vss 0.036697f
C6302 w_4660_n6791.n1806 vss 0.008764f
C6303 w_4660_n6791.n1807 vss 0.032221f
C6304 w_4660_n6791.n1808 vss 0.008764f
C6305 w_4660_n6791.n1809 vss 0.008764f
C6306 w_4660_n6791.n1810 vss 0.064443f
C6307 w_4660_n6791.n1811 vss 0.008764f
C6308 w_4660_n6791.n1812 vss 0.008764f
C6309 w_4660_n6791.n1813 vss 0.008764f
C6310 w_4660_n6791.n1814 vss 0.032221f
C6311 w_4660_n6791.n1815 vss 0.008764f
C6312 w_4660_n6791.n1816 vss 0.008764f
C6313 w_4660_n6791.n1817 vss 0.008764f
C6314 w_4660_n6791.n1818 vss 0.054598f
C6315 w_4660_n6791.n1819 vss 0.008764f
C6316 w_4660_n6791.n1820 vss 0.032221f
C6317 w_4660_n6791.n1821 vss 0.008764f
C6318 w_4660_n6791.n1822 vss 0.008764f
C6319 w_4660_n6791.n1823 vss 0.064443f
C6320 w_4660_n6791.n1824 vss 0.008764f
C6321 w_4660_n6791.n1825 vss 0.008764f
C6322 w_4660_n6791.n1826 vss 0.008764f
C6323 w_4660_n6791.n1827 vss 0.008764f
C6324 w_4660_n6791.n1828 vss 0.008764f
C6325 w_4660_n6791.n1829 vss 0.008764f
C6326 w_4660_n6791.n1830 vss 0.064443f
C6327 w_4660_n6791.n1831 vss 0.008764f
C6328 w_4660_n6791.n1832 vss 0.008764f
C6329 w_4660_n6791.n1833 vss 0.008764f
C6330 w_4660_n6791.n1834 vss 0.032221f
C6331 w_4660_n6791.n1835 vss 0.008764f
C6332 w_4660_n6791.n1836 vss 0.008764f
C6333 w_4660_n6791.n1837 vss 0.008764f
C6334 w_4660_n6791.n1838 vss 0.008764f
C6335 w_4660_n6791.n1839 vss 0.049227f
C6336 w_4660_n6791.n1840 vss 0.008764f
C6337 w_4660_n6791.n1841 vss 0.032221f
C6338 w_4660_n6791.n1842 vss 0.008764f
C6339 w_4660_n6791.n1843 vss 0.008764f
C6340 w_4660_n6791.n1844 vss 0.064443f
C6341 w_4660_n6791.n1845 vss 0.008764f
C6342 w_4660_n6791.n1846 vss 0.008764f
C6343 w_4660_n6791.n1847 vss 0.008764f
C6344 w_4660_n6791.n1848 vss 0.008764f
C6345 w_4660_n6791.n1849 vss 0.032221f
C6346 w_4660_n6791.n1850 vss 0.008764f
C6347 w_4660_n6791.n1851 vss 0.008764f
C6348 w_4660_n6791.n1852 vss 0.00633f
C6349 w_4660_n6791.n1853 vss 0.064443f
C6350 w_4660_n6791.n1854 vss 0.008764f
C6351 w_4660_n6791.n1855 vss 0.006817f
C6352 w_4660_n6791.n1856 vss 0.008764f
C6353 w_4660_n6791.n1857 vss 0.032221f
C6354 w_4660_n6791.n1858 vss 0.008764f
C6355 w_4660_n6791.n1859 vss 0.008764f
C6356 w_4660_n6791.n1860 vss 0.008764f
C6357 w_4660_n6791.n1861 vss 0.008764f
C6358 w_4660_n6791.n1862 vss 0.043857f
C6359 w_4660_n6791.n1863 vss 0.008764f
C6360 w_4660_n6791.n1864 vss 0.032221f
C6361 w_4660_n6791.n1865 vss 0.008764f
C6362 w_4660_n6791.n1866 vss 0.008764f
C6363 w_4660_n6791.n1867 vss 0.064443f
C6364 w_4660_n6791.n1868 vss 0.008764f
C6365 w_4660_n6791.n1869 vss 0.008764f
C6366 w_4660_n6791.n1870 vss 0.008764f
C6367 w_4660_n6791.n1871 vss 0.008764f
C6368 w_4660_n6791.n1872 vss 0.032221f
C6369 w_4660_n6791.n1873 vss 0.008764f
C6370 w_4660_n6791.n1874 vss 0.008764f
C6371 w_4660_n6791.n1875 vss 0.008764f
C6372 w_4660_n6791.n1876 vss 0.061758f
C6373 w_4660_n6791.n1877 vss 0.008764f
C6374 w_4660_n6791.n1878 vss 0.008764f
C6375 w_4660_n6791.n1879 vss 0.008764f
C6376 w_4660_n6791.n1880 vss 0.064443f
C6377 w_4660_n6791.n1881 vss 0.008764f
C6378 w_4660_n6791.n1882 vss 0.008764f
C6379 w_4660_n6791.n1883 vss 0.008764f
C6380 w_4660_n6791.n1884 vss 0.008764f
C6381 w_4660_n6791.n1885 vss 0.038487f
C6382 w_4660_n6791.n1886 vss 0.008764f
C6383 w_4660_n6791.n1887 vss 0.032221f
C6384 w_4660_n6791.n1888 vss 0.008764f
C6385 w_4660_n6791.n1889 vss 0.008764f
C6386 w_4660_n6791.n1890 vss 0.064443f
C6387 w_4660_n6791.n1891 vss 0.008764f
C6388 w_4660_n6791.n1892 vss 0.008764f
C6389 w_4660_n6791.n1893 vss 0.008764f
C6390 w_4660_n6791.n1894 vss 0.032221f
C6391 w_4660_n6791.n1895 vss 0.008764f
C6392 w_4660_n6791.n1896 vss 0.008764f
C6393 w_4660_n6791.n1897 vss 0.008764f
C6394 w_4660_n6791.n1898 vss 0.056388f
C6395 w_4660_n6791.n1899 vss 0.008764f
C6396 w_4660_n6791.n1900 vss 0.032221f
C6397 w_4660_n6791.n1901 vss 0.008764f
C6398 w_4660_n6791.n1902 vss 0.008764f
C6399 w_4660_n6791.n1903 vss 0.064443f
C6400 w_4660_n6791.n1904 vss 0.008764f
C6401 w_4660_n6791.n1905 vss 0.008764f
C6402 w_4660_n6791.n1906 vss 0.008764f
C6403 w_4660_n6791.n1907 vss 0.008764f
C6404 w_4660_n6791.n1908 vss 0.008764f
C6405 w_4660_n6791.n1909 vss 0.008764f
C6406 w_4660_n6791.n1910 vss 0.064443f
C6407 w_4660_n6791.n1911 vss 0.008764f
C6408 w_4660_n6791.n1912 vss 0.008764f
C6409 w_4660_n6791.n1913 vss 0.008764f
C6410 w_4660_n6791.n1914 vss 0.032221f
C6411 w_4660_n6791.n1915 vss 0.008764f
C6412 w_4660_n6791.n1916 vss 0.008764f
C6413 w_4660_n6791.n1917 vss 0.008764f
C6414 w_4660_n6791.n1918 vss 0.051017f
C6415 w_4660_n6791.n1919 vss 0.008764f
C6416 w_4660_n6791.n1920 vss 0.008764f
C6417 w_4660_n6791.t341 vss 0.031147f
C6418 w_4660_n6791.t312 vss 0.031147f
C6419 w_4660_n6791.n1921 vss 0.069153f
C6420 w_4660_n6791.n1922 vss 0.049976f
C6421 w_4660_n6791.n1923 vss 0.081778f
C6422 w_4660_n6791.t353 vss 0.031147f
C6423 w_4660_n6791.t380 vss 0.031147f
C6424 w_4660_n6791.n1924 vss 0.069153f
C6425 w_4660_n6791.n1925 vss 0.092379f
C6426 w_4660_n6791.n1926 vss 0.081778f
C6427 w_4660_n6791.t264 vss 0.031147f
C6428 w_4660_n6791.t386 vss 0.031147f
C6429 w_4660_n6791.n1927 vss 0.069153f
C6430 w_4660_n6791.n1928 vss 0.05149f
C6431 w_4660_n6791.n1929 vss 0.081778f
C6432 w_4660_n6791.t340 vss 0.031147f
C6433 w_4660_n6791.t370 vss 0.031147f
C6434 w_4660_n6791.n1930 vss 0.069153f
C6435 w_4660_n6791.n1931 vss 0.379156f
C6436 w_4660_n6791.n1932 vss 0.081778f
C6437 w_4660_n6791.t203 vss 0.031147f
C6438 w_4660_n6791.t378 vss 0.031147f
C6439 w_4660_n6791.n1933 vss 0.069153f
C6440 w_4660_n6791.n1934 vss 0.37966f
C6441 w_4660_n6791.t276 vss 0.031147f
C6442 w_4660_n6791.t236 vss 0.031147f
C6443 w_4660_n6791.n1935 vss 0.069153f
C6444 w_4660_n6791.n1936 vss 0.074711f
C6445 w_4660_n6791.t330 vss 0.031147f
C6446 w_4660_n6791.t347 vss 0.031147f
C6447 w_4660_n6791.n1937 vss 0.069153f
C6448 w_4660_n6791.n1938 vss 0.081778f
C6449 w_4660_n6791.t124 vss 0.031147f
C6450 w_4660_n6791.t457 vss 0.031147f
C6451 w_4660_n6791.n1939 vss 0.070394f
C6452 w_4660_n6791.n1940 vss 0.65226f
C6453 w_4660_n6791.t196 vss 0.031147f
C6454 w_4660_n6791.t367 vss 0.031147f
C6455 w_4660_n6791.n1941 vss 0.069153f
C6456 w_4660_n6791.n1942 vss 0.081778f
C6457 w_4660_n6791.t467 vss 0.031147f
C6458 w_4660_n6791.t474 vss 0.031147f
C6459 w_4660_n6791.n1943 vss 0.070394f
C6460 w_4660_n6791.n1944 vss 0.651755f
C6461 w_4660_n6791.t258 vss 0.031147f
C6462 w_4660_n6791.t224 vss 0.031147f
C6463 w_4660_n6791.n1945 vss 0.069153f
C6464 w_4660_n6791.n1946 vss 0.081778f
C6465 w_4660_n6791.t472 vss 0.031147f
C6466 w_4660_n6791.t21 vss 0.031147f
C6467 w_4660_n6791.n1947 vss 0.070394f
C6468 w_4660_n6791.n1948 vss 0.65226f
C6469 w_4660_n6791.t272 vss 0.031147f
C6470 w_4660_n6791.t232 vss 0.031147f
C6471 w_4660_n6791.n1949 vss 0.069153f
C6472 w_4660_n6791.n1950 vss 0.081778f
C6473 w_4660_n6791.t129 vss 0.031147f
C6474 w_4660_n6791.t19 vss 0.031147f
C6475 w_4660_n6791.n1951 vss 0.070394f
C6476 w_4660_n6791.n1952 vss 0.65226f
C6477 w_4660_n6791.t192 vss 0.031147f
C6478 w_4660_n6791.t354 vss 0.031147f
C6479 w_4660_n6791.n1953 vss 0.069153f
C6480 w_4660_n6791.n1954 vss 0.081273f
C6481 w_4660_n6791.t56 vss 0.031147f
C6482 w_4660_n6791.t414 vss 0.031147f
C6483 w_4660_n6791.n1955 vss 0.070394f
C6484 w_4660_n6791.n1956 vss 0.65226f
C6485 w_4660_n6791.t250 vss 0.031147f
C6486 w_4660_n6791.t208 vss 0.031147f
C6487 w_4660_n6791.n1957 vss 0.069153f
C6488 w_4660_n6791.n1958 vss 0.081778f
C6489 w_4660_n6791.t460 vss 0.12136f
C6490 w_4660_n6791.n1959 vss 0.663588f
C6491 w_4660_n6791.t263 vss 0.031147f
C6492 w_4660_n6791.t223 vss 0.031147f
C6493 w_4660_n6791.n1960 vss 0.069153f
C6494 w_4660_n6791.n1961 vss 0.081273f
C6495 w_4660_n6791.n1962 vss 0.063101f
C6496 w_4660_n6791.t322 vss 0.031147f
C6497 w_4660_n6791.t300 vss 0.031147f
C6498 w_4660_n6791.n1963 vss 0.069153f
C6499 w_4660_n6791.n1964 vss 0.048966f
C6500 w_4660_n6791.t459 vss 0.031147f
C6501 w_4660_n6791.t184 vss 0.031147f
C6502 w_4660_n6791.n1965 vss 0.070394f
C6503 w_4660_n6791.n1966 vss 0.65226f
C6504 w_4660_n6791.n1967 vss 0.045432f
C6505 w_4660_n6791.t69 vss 0.031147f
C6506 w_4660_n6791.t10 vss 0.031147f
C6507 w_4660_n6791.n1968 vss 0.070394f
C6508 w_4660_n6791.n1969 vss 0.65226f
C6509 w_4660_n6791.t316 vss 0.031147f
C6510 w_4660_n6791.t283 vss 0.031147f
C6511 w_4660_n6791.n1970 vss 0.069153f
C6512 w_4660_n6791.n1971 vss 0.42055f
C6513 w_4660_n6791.t461 vss 0.031147f
C6514 w_4660_n6791.t58 vss 0.031147f
C6515 w_4660_n6791.n1972 vss 0.070394f
C6516 w_4660_n6791.n1973 vss 0.65226f
C6517 w_4660_n6791.t328 vss 0.031147f
C6518 w_4660_n6791.t345 vss 0.031147f
C6519 w_4660_n6791.n1974 vss 0.069153f
C6520 w_4660_n6791.n1975 vss 0.37966f
C6521 w_4660_n6791.n1976 vss 0.047956f
C6522 w_4660_n6791.t247 vss 0.031147f
C6523 w_4660_n6791.t364 vss 0.031147f
C6524 w_4660_n6791.n1977 vss 0.069153f
C6525 w_4660_n6791.n1978 vss 0.37966f
C6526 w_4660_n6791.t315 vss 0.031147f
C6527 w_4660_n6791.t280 vss 0.031147f
C6528 w_4660_n6791.n1979 vss 0.069153f
C6529 w_4660_n6791.n1980 vss 0.37966f
C6530 w_4660_n6791.t326 vss 0.031147f
C6531 w_4660_n6791.t296 vss 0.031147f
C6532 w_4660_n6791.n1981 vss 0.069153f
C6533 w_4660_n6791.n1982 vss 0.379156f
C6534 w_4660_n6791.t468 vss 0.12136f
C6535 w_4660_n6791.n1983 vss 0.081778f
C6536 w_4660_n6791.n1984 vss 0.054014f
C6537 w_4660_n6791.n1985 vss 0.078749f
C6538 w_4660_n6791.t440 vss 0.031147f
C6539 w_4660_n6791.t20 vss 0.031147f
C6540 w_4660_n6791.n1986 vss 0.070394f
C6541 w_4660_n6791.n1987 vss 0.080769f
C6542 w_4660_n6791.n1988 vss 0.068149f
C6543 w_4660_n6791.n1989 vss 0.081778f
C6544 w_4660_n6791.n1990 vss 0.050985f
C6545 w_4660_n6791.n1991 vss 0.081778f
C6546 w_4660_n6791.t470 vss 0.031147f
C6547 w_4660_n6791.t452 vss 0.031147f
C6548 w_4660_n6791.n1992 vss 0.070394f
C6549 w_4660_n6791.n1993 vss 0.07774f
C6550 w_4660_n6791.n1994 vss 0.071682f
C6551 w_4660_n6791.n1995 vss 0.081778f
C6552 w_4660_n6791.n1996 vss 0.047452f
C6553 w_4660_n6791.n1997 vss 0.081778f
C6554 w_4660_n6791.t125 vss 0.031147f
C6555 w_4660_n6791.t146 vss 0.031147f
C6556 w_4660_n6791.n1998 vss 0.070394f
C6557 w_4660_n6791.n1999 vss 0.651755f
C6558 w_4660_n6791.n2000 vss 0.074206f
C6559 w_4660_n6791.n2001 vss 0.074711f
C6560 w_4660_n6791.n2002 vss 0.081273f
C6561 w_4660_n6791.n2003 vss 0.044423f
C6562 w_4660_n6791.n2004 vss 0.081778f
C6563 w_4660_n6791.n2005 vss 0.071177f
C6564 w_4660_n6791.n2006 vss 0.078245f
C6565 w_4660_n6791.n2007 vss 0.081778f
C6566 w_4660_n6791.n2008 vss 0.05149f
C6567 w_4660_n6791.n2009 vss 0.081778f
C6568 w_4660_n6791.n2010 vss 0.067644f
C6569 w_4660_n6791.n2011 vss 0.081778f
C6570 w_4660_n6791.t256 vss 0.031147f
C6571 w_4660_n6791.t214 vss 0.031147f
C6572 w_4660_n6791.n2012 vss 0.069153f
C6573 w_4660_n6791.n2013 vss 0.38067f
C6574 w_4660_n6791.n2014 vss 0.078245f
C6575 w_4660_n6791.n2015 vss 0.056033f
C6576 w_4660_n6791.n2016 vss 0.082788f
C6577 w_4660_n6791.n2017 vss 0.063101f
C6578 w_4660_n6791.n2018 vss 0.081778f
C6579 w_4660_n6791.t191 vss 0.031147f
C6580 w_4660_n6791.t355 vss 0.031147f
C6581 w_4660_n6791.n2019 vss 0.069153f
C6582 w_4660_n6791.n2020 vss 0.37966f
C6583 w_4660_n6791.n2021 vss 0.073701f
C6584 w_4660_n6791.n2022 vss 0.059567f
C6585 w_4660_n6791.n2023 vss 0.081778f
C6586 w_4660_n6791.t82 vss 0.031147f
C6587 w_4660_n6791.t433 vss 0.031147f
C6588 w_4660_n6791.n2024 vss 0.070394f
C6589 w_4660_n6791.n2025 vss 0.65226f
C6590 w_4660_n6791.n2026 vss 0.059567f
C6591 w_4660_n6791.n2027 vss 0.081778f
C6592 w_4660_n6791.n2028 vss 0.070168f
C6593 w_4660_n6791.n2029 vss 0.37966f
C6594 w_4660_n6791.n2030 vss 0.051995f
C6595 w_4660_n6791.n2031 vss 0.081273f
C6596 w_4660_n6791.n2032 vss 0.081273f
C6597 w_4660_n6791.n2033 vss 0.071177f
C6598 w_4660_n6791.n2034 vss 0.067139f
C6599 w_4660_n6791.n2035 vss 0.37966f
C6600 w_4660_n6791.n2036 vss 0.055528f
C6601 w_4660_n6791.n2037 vss 0.05149f
C6602 w_4660_n6791.n2038 vss 0.081778f
C6603 w_4660_n6791.n2039 vss 0.067644f
C6604 w_4660_n6791.n2040 vss 0.063605f
C6605 w_4660_n6791.n2041 vss 0.37966f
C6606 w_4660_n6791.n2042 vss 0.059062f
C6607 w_4660_n6791.n2043 vss 0.055024f
C6608 w_4660_n6791.n2044 vss 0.081273f
C6609 w_4660_n6791.n2045 vss 0.06411f
C6610 w_4660_n6791.n2046 vss 0.060072f
C6611 w_4660_n6791.n2047 vss 0.37966f
C6612 w_4660_n6791.n2048 vss 0.062091f
C6613 w_4660_n6791.n2049 vss 0.058052f
C6614 w_4660_n6791.n2050 vss 0.081778f
C6615 w_4660_n6791.n2051 vss 0.061081f
C6616 w_4660_n6791.n2052 vss 0.057043f
C6617 w_4660_n6791.n2053 vss 0.37966f
C6618 w_4660_n6791.n2054 vss 0.065624f
C6619 w_4660_n6791.n2055 vss 0.061586f
C6620 w_4660_n6791.n2056 vss 0.081778f
C6621 w_4660_n6791.n2057 vss 0.057548f
C6622 w_4660_n6791.n2058 vss 0.053509f
C6623 w_4660_n6791.n2059 vss 0.379156f
C6624 w_4660_n6791.n2060 vss 0.068653f
C6625 w_4660_n6791.n2061 vss 0.064615f
C6626 w_4660_n6791.n2062 vss 0.081778f
C6627 w_4660_n6791.n2063 vss 0.054519f
C6628 w_4660_n6791.n2064 vss 0.05048f
C6629 w_4660_n6791.n2065 vss 0.37966f
C6630 w_4660_n6791.n2066 vss 0.072187f
C6631 w_4660_n6791.n2067 vss 0.068149f
C6632 w_4660_n6791.n2068 vss 0.081778f
C6633 w_4660_n6791.t473 vss 0.031147f
C6634 w_4660_n6791.t57 vss 0.031147f
C6635 w_4660_n6791.n2069 vss 0.070394f
C6636 w_4660_n6791.n2070 vss 0.65226f
C6637 w_4660_n6791.n2071 vss 0.050985f
C6638 w_4660_n6791.n2072 vss 0.046947f
C6639 w_4660_n6791.n2073 vss 0.37966f
C6640 w_4660_n6791.n2074 vss 0.078749f
C6641 w_4660_n6791.n2075 vss 0.084302f
C6642 w_4660_n6791.n2076 vss 0.084807f
C6643 w_4660_n6791.t97 vss 0.031147f
C6644 w_4660_n6791.t22 vss 0.031147f
C6645 w_4660_n6791.n2077 vss 0.070394f
C6646 w_4660_n6791.n2078 vss 0.081778f
C6647 w_4660_n6791.n2079 vss 0.07774f
C6648 w_4660_n6791.n2080 vss 0.081778f
C6649 w_4660_n6791.n2081 vss 0.081778f
C6650 w_4660_n6791.n2082 vss 0.044928f
C6651 w_4660_n6791.n2083 vss 0.081778f
C6652 w_4660_n6791.n2084 vss 0.074206f
C6653 w_4660_n6791.n2085 vss 0.081273f
C6654 w_4660_n6791.n2086 vss 0.081273f
C6655 w_4660_n6791.n2087 vss 0.047956f
C6656 w_4660_n6791.n2088 vss 0.081778f
C6657 w_4660_n6791.t332 vss 0.031147f
C6658 w_4660_n6791.t303 vss 0.031147f
C6659 w_4660_n6791.n2089 vss 0.069153f
C6660 w_4660_n6791.n2090 vss 0.37966f
C6661 w_4660_n6791.n2091 vss 0.071177f
C6662 w_4660_n6791.n2092 vss 0.081778f
C6663 w_4660_n6791.n2093 vss 0.081778f
C6664 w_4660_n6791.n2094 vss 0.081778f
C6665 w_4660_n6791.n2095 vss 0.081778f
C6666 w_4660_n6791.n2096 vss 0.067644f
C6667 w_4660_n6791.n2097 vss 0.37966f
C6668 w_4660_n6791.n2098 vss 0.065624f
C6669 w_4660_n6791.n2099 vss 0.092379f
C6670 w_4660_n6791.n2100 vss 0.092379f
C6671 w_4660_n6791.n2101 vss 0.081778f
C6672 w_4660_n6791.n2102 vss 0.053509f
C6673 w_4660_n6791.n2103 vss 0.37966f
C6674 w_4660_n6791.n2104 vss 0.069158f
C6675 w_4660_n6791.n2105 vss 0.081778f
C6676 w_4660_n6791.n2106 vss 0.081778f
C6677 w_4660_n6791.n2107 vss 0.081778f
C6678 w_4660_n6791.n2108 vss 0.092379f
C6679 w_4660_n6791.n2109 vss 0.081778f
C6680 w_4660_n6791.n2110 vss 0.072692f
C6681 w_4660_n6791.n2111 vss 0.37966f
C6682 w_4660_n6791.n2112 vss 0.032221f
C6683 w_4660_n6791.n2113 vss 0.008764f
C6684 w_4660_n6791.n2114 vss 0.008764f
C6685 w_4660_n6791.n2115 vss 0.008764f
C6686 w_4660_n6791.n2116 vss 0.008764f
C6687 w_4660_n6791.n2117 vss 0.064443f
C6688 w_4660_n6791.n2118 vss 0.008764f
C6689 w_4660_n6791.n2119 vss 0.008764f
C6690 w_4660_n6791.n2120 vss 0.008764f
C6691 w_4660_n6791.n2121 vss 0.045647f
C6692 w_4660_n6791.n2122 vss 0.008764f
C6693 w_4660_n6791.n2123 vss 0.008764f
C6694 w_4660_n6791.n2124 vss 0.008764f
C6695 w_4660_n6791.n2125 vss 0.064443f
C6696 w_4660_n6791.n2126 vss 0.054598f
C6697 w_4660_n6791.n2127 vss 0.008764f
C6698 w_4660_n6791.n2128 vss 0.008764f
C6699 w_4660_n6791.n2129 vss 0.042067f
C6700 w_4660_n6791.n2130 vss 0.008764f
C6701 w_4660_n6791.n2131 vss 0.008764f
C6702 w_4660_n6791.n2132 vss 0.008764f
C6703 w_4660_n6791.n2133 vss 0.063548f
C6704 w_4660_n6791.n2134 vss 0.008764f
C6705 w_4660_n6791.n2135 vss 0.008764f
C6706 w_4660_n6791.n2136 vss 0.008764f
C6707 w_4660_n6791.n2137 vss 0.064443f
C6708 w_4660_n6791.n2138 vss 0.008764f
C6709 w_4660_n6791.n2139 vss 0.008764f
C6710 w_4660_n6791.n2140 vss 0.008764f
C6711 w_4660_n6791.n2141 vss 0.040277f
C6712 w_4660_n6791.n2142 vss 0.008764f
C6713 w_4660_n6791.n2143 vss 0.008764f
C6714 w_4660_n6791.n2144 vss 0.008764f
C6715 w_4660_n6791.n2145 vss 0.064443f
C6716 w_4660_n6791.n2146 vss 0.049227f
C6717 w_4660_n6791.n2147 vss 0.008764f
C6718 w_4660_n6791.n2148 vss 0.008764f
C6719 w_4660_n6791.n2149 vss 0.047437f
C6720 w_4660_n6791.n2150 vss 0.008764f
C6721 w_4660_n6791.n2151 vss 0.008764f
C6722 w_4660_n6791.n2152 vss 0.008764f
C6723 w_4660_n6791.n2153 vss 0.058178f
C6724 w_4660_n6791.n2154 vss 0.008764f
C6725 w_4660_n6791.n2155 vss 0.008764f
C6726 w_4660_n6791.n2156 vss 0.008764f
C6727 w_4660_n6791.n2157 vss 0.064443f
C6728 w_4660_n6791.n2158 vss 0.008764f
C6729 w_4660_n6791.n2159 vss 0.008764f
C6730 w_4660_n6791.n2160 vss 0.008764f
C6731 w_4660_n6791.n2161 vss 0.034907f
C6732 w_4660_n6791.n2162 vss 0.008764f
C6733 w_4660_n6791.n2163 vss 0.008764f
C6734 w_4660_n6791.n2164 vss 0.008764f
C6735 w_4660_n6791.n2165 vss 0.064443f
C6736 w_4660_n6791.n2166 vss 0.043857f
C6737 w_4660_n6791.n2167 vss 0.008764f
C6738 w_4660_n6791.n2168 vss 0.008764f
C6739 w_4660_n6791.n2169 vss 0.052807f
C6740 w_4660_n6791.n2170 vss 0.008764f
C6741 w_4660_n6791.n2171 vss 0.008764f
C6742 w_4660_n6791.n2172 vss 0.008764f
C6743 w_4660_n6791.n2173 vss 0.052807f
C6744 w_4660_n6791.n2174 vss 0.008764f
C6745 w_4660_n6791.n2175 vss 0.008764f
C6746 w_4660_n6791.n2176 vss 0.008764f
C6747 w_4660_n6791.n2177 vss 0.064443f
C6748 w_4660_n6791.n2178 vss 0.061758f
C6749 w_4660_n6791.n2179 vss 0.008764f
C6750 w_4660_n6791.n2180 vss 0.008764f
C6751 w_4660_n6791.n2181 vss 0.034907f
C6752 w_4660_n6791.n2182 vss 0.008764f
C6753 w_4660_n6791.n2183 vss 0.006817f
C6754 w_4660_n6791.n2184 vss 0.004382f
C6755 w_4660_n6791.n2185 vss 0.00633f
C6756 w_4660_n6791.n2186 vss 0.064443f
C6757 w_4660_n6791.n2187 vss 0.038487f
C6758 w_4660_n6791.n2188 vss 0.008764f
C6759 w_4660_n6791.n2189 vss 0.008764f
C6760 w_4660_n6791.n2190 vss 0.058178f
C6761 w_4660_n6791.n2191 vss 0.008764f
C6762 w_4660_n6791.n2192 vss 0.008764f
C6763 w_4660_n6791.n2193 vss 0.008764f
C6764 w_4660_n6791.n2194 vss 0.047437f
C6765 w_4660_n6791.n2195 vss 0.008764f
C6766 w_4660_n6791.n2196 vss 0.008764f
C6767 w_4660_n6791.n2197 vss 0.008764f
C6768 w_4660_n6791.n2198 vss 0.064443f
C6769 w_4660_n6791.n2199 vss 0.056388f
C6770 w_4660_n6791.n2200 vss 0.008764f
C6771 w_4660_n6791.n2201 vss 0.008764f
C6772 w_4660_n6791.n2202 vss 0.040277f
C6773 w_4660_n6791.n2203 vss 0.008764f
C6774 w_4660_n6791.n2204 vss 0.008764f
C6775 w_4660_n6791.n2205 vss 0.008764f
C6776 w_4660_n6791.n2206 vss 0.064443f
C6777 w_4660_n6791.n2207 vss 0.008764f
C6778 w_4660_n6791.n2208 vss 0.008764f
C6779 w_4660_n6791.n2209 vss 0.063548f
C6780 w_4660_n6791.n2210 vss 0.008764f
C6781 w_4660_n6791.n2211 vss 0.008764f
C6782 w_4660_n6791.n2212 vss 0.008764f
C6783 w_4660_n6791.n2213 vss 0.042067f
C6784 w_4660_n6791.n2214 vss 0.008764f
C6785 w_4660_n6791.n2215 vss 0.008764f
C6786 w_4660_n6791.n2216 vss 0.008764f
C6787 w_4660_n6791.n2217 vss 0.064443f
C6788 w_4660_n6791.n2218 vss 0.051017f
C6789 w_4660_n6791.n2219 vss 0.008764f
C6790 w_4660_n6791.n2220 vss 0.008764f
C6791 w_4660_n6791.n2221 vss 0.045647f
C6792 w_4660_n6791.n2222 vss 0.008764f
C6793 w_4660_n6791.n2223 vss 0.008764f
C6794 w_4660_n6791.n2224 vss 0.008764f
C6795 w_4660_n6791.n2225 vss 0.059968f
C6796 w_4660_n6791.n2226 vss 0.008764f
C6797 w_4660_n6791.n2227 vss 0.008764f
C6798 w_4660_n6791.n2228 vss 0.008764f
C6799 w_4660_n6791.n2229 vss 0.064443f
C6800 w_4660_n6791.n2230 vss 0.008764f
C6801 w_4660_n6791.n2231 vss 0.008764f
C6802 w_4660_n6791.n2232 vss 0.008764f
C6803 w_4660_n6791.n2233 vss 0.036697f
C6804 w_4660_n6791.n2234 vss 0.008764f
C6805 w_4660_n6791.n2235 vss 0.008764f
C6806 w_4660_n6791.n2236 vss 0.008764f
C6807 w_4660_n6791.n2237 vss 0.064443f
C6808 w_4660_n6791.n2238 vss 0.045647f
C6809 w_4660_n6791.n2239 vss 0.008764f
C6810 w_4660_n6791.n2240 vss 0.008764f
C6811 w_4660_n6791.n2241 vss 0.051017f
C6812 w_4660_n6791.n2242 vss 0.008764f
C6813 w_4660_n6791.n2243 vss 0.008764f
C6814 w_4660_n6791.n2244 vss 0.008764f
C6815 w_4660_n6791.n2245 vss 0.054598f
C6816 w_4660_n6791.n2246 vss 0.008764f
C6817 w_4660_n6791.n2247 vss 0.008764f
C6818 w_4660_n6791.n2248 vss 0.008764f
C6819 w_4660_n6791.n2249 vss 0.064443f
C6820 w_4660_n6791.n2250 vss 0.063548f
C6821 w_4660_n6791.n2251 vss 0.008764f
C6822 w_4660_n6791.n2252 vss 0.008764f
C6823 w_4660_n6791.n2253 vss 0.008764f
C6824 w_4660_n6791.n2254 vss 0.008764f
C6825 w_4660_n6791.n2255 vss 0.008764f
C6826 w_4660_n6791.n2256 vss 0.064443f
C6827 w_4660_n6791.n2257 vss 0.040277f
C6828 w_4660_n6791.n2258 vss 0.008764f
C6829 w_4660_n6791.n2259 vss 0.008764f
C6830 w_4660_n6791.n2260 vss 0.056388f
C6831 w_4660_n6791.n2261 vss 0.008764f
C6832 w_4660_n6791.n2262 vss 0.008764f
C6833 w_4660_n6791.n2263 vss 0.008764f
C6834 w_4660_n6791.n2264 vss 0.049227f
C6835 w_4660_n6791.n2265 vss 0.032221f
C6836 w_4660_n6791.n2266 vss 0.390843f
C6837 w_4660_n6791.n2267 vss 0.057548f
C6838 w_4660_n6791.n2268 vss 0.081778f
C6839 w_4660_n6791.n2269 vss 0.081778f
C6840 w_4660_n6791.n2271 vss 0.242907f
C6841 w_4660_n6791.n2272 vss 0.100456f
C6842 w_4660_n6791.n2273 vss 2.70648f
C6843 w_4660_n6791.n2274 vss 5.443491f
C6844 w_4660_n6791.n2275 vss 5.70848f
C6845 w_4660_n6791.n2276 vss 6.04988f
C6846 w_4660_n6791.n2277 vss 3.00823f
C6847 w_4660_n6791.n2278 vss 0.056388f
C6848 w_4660_n6791.n2279 vss 0.008764f
C6849 w_4660_n6791.n2280 vss 0.008764f
C6850 w_4660_n6791.n2281 vss 0.008764f
C6851 w_4660_n6791.n2282 vss 0.064443f
C6852 w_4660_n6791.n2283 vss 0.01035f
C6853 w_4660_n6791.n2284 vss 0.049227f
C6854 w_4660_n6791.n2285 vss 0.032221f
C6855 w_4660_n6791.n2286 vss 0.073874f
C6856 w_4660_n6791.n2287 vss 0.5592f
C6857 w_4660_n6791.n2288 vss 0.011345f
C6858 w_4660_n6791.n2289 vss 0.008764f
C6859 w_4660_n6791.n2290 vss 0.008764f
C6860 w_4660_n6791.n2291 vss 0.064443f
C6861 w_4660_n6791.n2292 vss 0.008764f
C6862 w_4660_n6791.n2293 vss 0.008764f
C6863 w_4660_n6791.n2294 vss 0.008764f
C6864 w_4660_n6791.n2295 vss 0.008764f
C6865 w_4660_n6791.n2296 vss 0.040277f
C6866 w_4660_n6791.n2297 vss 0.032221f
C6867 w_4660_n6791.n2298 vss 0.549171f
C6868 w_4660_n6791.t398 vss 0.031147f
C6869 w_4660_n6791.t432 vss 0.031147f
C6870 w_4660_n6791.n2299 vss 0.069153f
C6871 w_4660_n6791.n2300 vss 0.549171f
C6872 w_4660_n6791.n2301 vss 0.549171f
C6873 w_4660_n6791.n2302 vss 0.008764f
C6874 w_4660_n6791.n2303 vss 0.008764f
C6875 w_4660_n6791.n2304 vss 0.008764f
C6876 w_4660_n6791.n2305 vss 0.064443f
C6877 w_4660_n6791.n2306 vss 0.042067f
C6878 w_4660_n6791.n2307 vss 0.008764f
C6879 w_4660_n6791.n2308 vss 0.008764f
C6880 w_4660_n6791.n2309 vss 0.054598f
C6881 w_4660_n6791.n2310 vss 0.008764f
C6882 w_4660_n6791.n2311 vss 0.008764f
C6883 w_4660_n6791.n2312 vss 0.008764f
C6884 w_4660_n6791.n2313 vss 0.051017f
C6885 w_4660_n6791.n2314 vss 0.008764f
C6886 w_4660_n6791.n2315 vss 0.008764f
C6887 w_4660_n6791.n2316 vss 0.008764f
C6888 w_4660_n6791.n2317 vss 0.008764f
C6889 w_4660_n6791.n2318 vss 0.064443f
C6890 w_4660_n6791.n2319 vss 0.008764f
C6891 w_4660_n6791.n2320 vss 0.008764f
C6892 w_4660_n6791.n2321 vss 0.008764f
C6893 w_4660_n6791.n2322 vss 0.008764f
C6894 w_4660_n6791.n2323 vss 0.036697f
C6895 w_4660_n6791.n2324 vss 0.032221f
C6896 w_4660_n6791.n2325 vss 0.549171f
C6897 w_4660_n6791.t81 vss 0.031147f
C6898 w_4660_n6791.t431 vss 0.031147f
C6899 w_4660_n6791.n2326 vss 0.069153f
C6900 w_4660_n6791.n2327 vss 0.549171f
C6901 w_4660_n6791.n2328 vss 0.549171f
C6902 w_4660_n6791.n2329 vss 0.032221f
C6903 w_4660_n6791.n2330 vss 0.036697f
C6904 w_4660_n6791.n2331 vss 0.008764f
C6905 w_4660_n6791.n2332 vss 0.008764f
C6906 w_4660_n6791.n2333 vss 0.008764f
C6907 w_4660_n6791.n2334 vss 0.064443f
C6908 w_4660_n6791.n2335 vss 0.045647f
C6909 w_4660_n6791.n2336 vss 0.008764f
C6910 w_4660_n6791.n2337 vss 0.008764f
C6911 w_4660_n6791.n2338 vss 0.051017f
C6912 w_4660_n6791.n2339 vss 0.008764f
C6913 w_4660_n6791.n2340 vss 0.008764f
C6914 w_4660_n6791.n2341 vss 0.008764f
C6915 w_4660_n6791.n2342 vss 0.054598f
C6916 w_4660_n6791.n2343 vss 0.008764f
C6917 w_4660_n6791.n2344 vss 0.008764f
C6918 w_4660_n6791.n2345 vss 0.008764f
C6919 w_4660_n6791.n2346 vss 0.008764f
C6920 w_4660_n6791.n2347 vss 0.064443f
C6921 w_4660_n6791.n2348 vss 0.008764f
C6922 w_4660_n6791.n2349 vss 0.008764f
C6923 w_4660_n6791.n2350 vss 0.008764f
C6924 w_4660_n6791.n2351 vss 0.008764f
C6925 w_4660_n6791.n2352 vss 0.549171f
C6926 w_4660_n6791.t91 vss 0.031147f
C6927 w_4660_n6791.t89 vss 0.031147f
C6928 w_4660_n6791.n2353 vss 0.069153f
C6929 w_4660_n6791.t162 vss 0.031147f
C6930 w_4660_n6791.t160 vss 0.031147f
C6931 w_4660_n6791.n2354 vss 0.069153f
C6932 w_4660_n6791.n2355 vss 0.549171f
C6933 w_4660_n6791.n2356 vss 0.549171f
C6934 w_4660_n6791.n2357 vss 0.549171f
C6935 w_4660_n6791.n2358 vss 0.032221f
C6936 w_4660_n6791.n2359 vss 0.040277f
C6937 w_4660_n6791.n2360 vss 0.008764f
C6938 w_4660_n6791.n2361 vss 0.008764f
C6939 w_4660_n6791.n2362 vss 0.008764f
C6940 w_4660_n6791.n2363 vss 0.064443f
C6941 w_4660_n6791.n2364 vss 0.049227f
C6942 w_4660_n6791.n2365 vss 0.008764f
C6943 w_4660_n6791.n2366 vss 0.008764f
C6944 w_4660_n6791.n2367 vss 0.047437f
C6945 w_4660_n6791.n2368 vss 0.008764f
C6946 w_4660_n6791.n2369 vss 0.008764f
C6947 w_4660_n6791.n2370 vss 0.008764f
C6948 w_4660_n6791.n2371 vss 0.058178f
C6949 w_4660_n6791.n2372 vss 0.008764f
C6950 w_4660_n6791.n2373 vss 0.008764f
C6951 w_4660_n6791.n2374 vss 0.00633f
C6952 w_4660_n6791.n2375 vss 0.064443f
C6953 w_4660_n6791.n2376 vss 0.00633f
C6954 w_4660_n6791.n2377 vss 0.004382f
C6955 w_4660_n6791.n2378 vss 0.006817f
C6956 w_4660_n6791.n2379 vss 0.008764f
C6957 w_4660_n6791.n2380 vss 0.034907f
C6958 w_4660_n6791.n2381 vss 0.008764f
C6959 w_4660_n6791.n2382 vss 0.008764f
C6960 w_4660_n6791.n2383 vss 0.008764f
C6961 w_4660_n6791.n2384 vss 0.008764f
C6962 w_4660_n6791.n2385 vss 0.064443f
C6963 w_4660_n6791.n2386 vss 0.008764f
C6964 w_4660_n6791.n2387 vss 0.008764f
C6965 w_4660_n6791.n2388 vss 0.008764f
C6966 w_4660_n6791.n2389 vss 0.052807f
C6967 w_4660_n6791.n2390 vss 0.032221f
C6968 w_4660_n6791.n2391 vss 0.549171f
C6969 w_4660_n6791.t1 vss 0.031147f
C6970 w_4660_n6791.t448 vss 0.031147f
C6971 w_4660_n6791.n2392 vss 0.069153f
C6972 w_4660_n6791.t412 vss 0.031147f
C6973 w_4660_n6791.t411 vss 0.031147f
C6974 w_4660_n6791.n2393 vss 0.069153f
C6975 w_4660_n6791.n2394 vss 0.549171f
C6976 w_4660_n6791.n2395 vss 0.549171f
C6977 w_4660_n6791.n2396 vss 0.549171f
C6978 w_4660_n6791.n2397 vss 0.032221f
C6979 w_4660_n6791.n2398 vss 0.052807f
C6980 w_4660_n6791.n2399 vss 0.008764f
C6981 w_4660_n6791.n2400 vss 0.008764f
C6982 w_4660_n6791.n2401 vss 0.008764f
C6983 w_4660_n6791.n2402 vss 0.064443f
C6984 w_4660_n6791.n2403 vss 0.061758f
C6985 w_4660_n6791.n2404 vss 0.008764f
C6986 w_4660_n6791.n2405 vss 0.008764f
C6987 w_4660_n6791.n2406 vss 0.008764f
C6988 w_4660_n6791.n2407 vss 0.034907f
C6989 w_4660_n6791.n2408 vss 0.008764f
C6990 w_4660_n6791.n2409 vss 0.008764f
C6991 w_4660_n6791.n2410 vss 0.008764f
C6992 w_4660_n6791.n2411 vss 0.064443f
C6993 w_4660_n6791.n2412 vss 0.038487f
C6994 w_4660_n6791.n2413 vss 0.008764f
C6995 w_4660_n6791.n2414 vss 0.008764f
C6996 w_4660_n6791.n2415 vss 0.058178f
C6997 w_4660_n6791.n2416 vss 0.008764f
C6998 w_4660_n6791.n2417 vss 0.008764f
C6999 w_4660_n6791.n2418 vss 0.008764f
C7000 w_4660_n6791.n2419 vss 0.047437f
C7001 w_4660_n6791.n2420 vss 0.008764f
C7002 w_4660_n6791.n2421 vss 0.008764f
C7003 w_4660_n6791.n2422 vss 0.008764f
C7004 w_4660_n6791.n2423 vss 0.008764f
C7005 w_4660_n6791.n2424 vss 0.064443f
C7006 w_4660_n6791.n2425 vss 0.008764f
C7007 w_4660_n6791.n2426 vss 0.008764f
C7008 w_4660_n6791.n2427 vss 0.008764f
C7009 w_4660_n6791.n2428 vss 0.008764f
C7010 w_4660_n6791.n2429 vss 0.040277f
C7011 w_4660_n6791.n2430 vss 0.032221f
C7012 w_4660_n6791.n2431 vss 0.549171f
C7013 w_4660_n6791.t6 vss 0.031147f
C7014 w_4660_n6791.t455 vss 0.031147f
C7015 w_4660_n6791.n2432 vss 0.069153f
C7016 w_4660_n6791.n2433 vss 0.549171f
C7017 w_4660_n6791.n2434 vss 0.549171f
C7018 w_4660_n6791.n2435 vss 0.008764f
C7019 w_4660_n6791.n2436 vss 0.008764f
C7020 w_4660_n6791.n2437 vss 0.008764f
C7021 w_4660_n6791.n2438 vss 0.064443f
C7022 w_4660_n6791.n2439 vss 0.042067f
C7023 w_4660_n6791.n2440 vss 0.008764f
C7024 w_4660_n6791.n2441 vss 0.008764f
C7025 w_4660_n6791.n2442 vss 0.054598f
C7026 w_4660_n6791.n2443 vss 0.008764f
C7027 w_4660_n6791.n2444 vss 0.008764f
C7028 w_4660_n6791.n2445 vss 0.008764f
C7029 w_4660_n6791.n2446 vss 0.051017f
C7030 w_4660_n6791.n2447 vss 0.008764f
C7031 w_4660_n6791.n2448 vss 0.008764f
C7032 w_4660_n6791.n2449 vss 0.008764f
C7033 w_4660_n6791.n2450 vss 0.008764f
C7034 w_4660_n6791.n2451 vss 0.064443f
C7035 w_4660_n6791.n2452 vss 0.008764f
C7036 w_4660_n6791.n2453 vss 0.008764f
C7037 w_4660_n6791.n2454 vss 0.008764f
C7038 w_4660_n6791.n2455 vss 0.008764f
C7039 w_4660_n6791.n2456 vss 0.036697f
C7040 w_4660_n6791.n2457 vss 0.032221f
C7041 w_4660_n6791.n2458 vss 0.549171f
C7042 w_4660_n6791.t425 vss 0.120265f
C7043 w_4660_n6791.n2459 vss 0.514524f
C7044 w_4660_n6791.n2460 vss 0.549171f
C7045 w_4660_n6791.n2461 vss 0.032221f
C7046 w_4660_n6791.n2462 vss 0.036697f
C7047 w_4660_n6791.n2463 vss 0.008764f
C7048 w_4660_n6791.n2464 vss 0.008764f
C7049 w_4660_n6791.n2465 vss 0.008764f
C7050 w_4660_n6791.n2466 vss 0.064443f
C7051 w_4660_n6791.n2467 vss 0.045647f
C7052 w_4660_n6791.n2468 vss 0.010661f
C7053 w_4660_n6791.n2469 vss 0.102211f
C7054 w_4660_n6791.n2470 vss 0.014816f
C7055 w_4660_n6791.n2471 vss 0.015057f
C7056 w_4660_n6791.n2472 vss 0.009022f
C7057 w_4660_n6791.n2473 vss 0.061865f
C7058 w_4660_n6791.n2474 vss 0.008912f
C7059 w_4660_n6791.n2475 vss 0.011198f
C7060 w_4660_n6791.n2476 vss 0.008764f
C7061 w_4660_n6791.n2477 vss 0.061865f
C7062 w_4660_n6791.n2478 vss 0.009022f
C7063 w_4660_n6791.n2479 vss 0.009022f
C7064 w_4660_n6791.n2480 vss 0.009022f
C7065 w_4660_n6791.n2481 vss 0.061865f
C7066 w_4660_n6791.n2482 vss 0.008764f
C7067 w_4660_n6791.n2483 vss 0.008764f
C7068 w_4660_n6791.n2484 vss 0.008764f
C7069 w_4660_n6791.n2485 vss 0.061865f
C7070 w_4660_n6791.n2486 vss 0.009022f
C7071 w_4660_n6791.n2487 vss 0.009022f
C7072 w_4660_n6791.n2488 vss 0.009022f
C7073 w_4660_n6791.n2489 vss 0.061865f
C7074 w_4660_n6791.n2490 vss 0.008764f
C7075 w_4660_n6791.n2491 vss 0.008764f
C7076 w_4660_n6791.n2492 vss 0.008764f
C7077 w_4660_n6791.n2493 vss 0.061865f
C7078 w_4660_n6791.n2494 vss 0.004948f
C7079 w_4660_n6791.n2495 vss 0.009022f
C7080 w_4660_n6791.n2496 vss 0.009022f
C7081 w_4660_n6791.n2497 vss 0.061865f
C7082 w_4660_n6791.n2498 vss 0.008764f
C7083 w_4660_n6791.n2499 vss 0.008764f
C7084 w_4660_n6791.n2500 vss 0.008764f
C7085 w_4660_n6791.n2501 vss 0.061865f
C7086 w_4660_n6791.n2502 vss 0.009022f
C7087 w_4660_n6791.n2503 vss 0.009022f
C7088 w_4660_n6791.n2504 vss 0.009022f
C7089 w_4660_n6791.n2505 vss 0.061865f
C7090 w_4660_n6791.n2506 vss 0.008764f
C7091 w_4660_n6791.n2507 vss 0.008764f
C7092 w_4660_n6791.n2508 vss 0.008764f
C7093 w_4660_n6791.n2509 vss 0.061865f
C7094 w_4660_n6791.n2510 vss 0.009022f
C7095 w_4660_n6791.n2511 vss 0.009022f
C7096 w_4660_n6791.n2512 vss 0.009022f
C7097 w_4660_n6791.n2513 vss 0.061865f
C7098 w_4660_n6791.n2514 vss 0.008764f
C7099 w_4660_n6791.n2515 vss 0.008764f
C7100 w_4660_n6791.n2516 vss 0.008764f
C7101 w_4660_n6791.n2517 vss 0.061865f
C7102 w_4660_n6791.n2518 vss 0.005324f
C7103 w_4660_n6791.n2519 vss 0.189923f
C7104 w_4660_n6791.n2520 vss 0.425158f
C7105 w_4660_n6791.n2521 vss 0.479417f
C7106 w_4660_n6791.n2522 vss -2.62744f
C7107 w_4660_n6791.n2523 vss -0.361891f
C7108 w_4660_n6791.n2524 vss 0.006817f
C7109 w_4660_n6791.n2525 vss 0.008764f
C7110 w_4660_n6791.n2526 vss 0.034907f
C7111 w_4660_n6791.n2527 vss 0.008764f
C7112 w_4660_n6791.n2528 vss 0.008764f
C7113 w_4660_n6791.n2529 vss 0.061758f
C7114 w_4660_n6791.n2530 vss 0.008764f
C7115 w_4660_n6791.n2531 vss 0.008764f
C7116 w_4660_n6791.n2532 vss 0.008764f
C7117 w_4660_n6791.n2533 vss 0.043857f
C7118 w_4660_n6791.n2534 vss 0.008764f
C7119 w_4660_n6791.n2535 vss 0.008764f
C7120 w_4660_n6791.n2536 vss 0.052807f
C7121 w_4660_n6791.n2537 vss 0.008764f
C7122 w_4660_n6791.n2538 vss 0.008764f
C7123 w_4660_n6791.n2539 vss 0.008764f
C7124 w_4660_n6791.n2540 vss 0.052807f
C7125 w_4660_n6791.n2541 vss 0.008764f
C7126 w_4660_n6791.n2542 vss 0.008764f
C7127 w_4660_n6791.n2543 vss 0.043857f
C7128 w_4660_n6791.n2544 vss 0.008764f
C7129 w_4660_n6791.n2545 vss 0.008764f
C7130 w_4660_n6791.n2546 vss 0.008764f
C7131 w_4660_n6791.n2547 vss 0.061758f
C7132 w_4660_n6791.n2548 vss 0.008764f
C7133 w_4660_n6791.n2549 vss 0.008764f
C7134 w_4660_n6791.n2550 vss 0.008764f
C7135 w_4660_n6791.n2551 vss 0.064443f
C7136 w_4660_n6791.n2552 vss 0.008764f
C7137 w_4660_n6791.n2553 vss 0.008764f
C7138 w_4660_n6791.n2554 vss 0.008764f
C7139 w_4660_n6791.n2555 vss 0.038487f
C7140 w_4660_n6791.n2556 vss 0.008764f
C7141 w_4660_n6791.n2557 vss 0.008764f
C7142 w_4660_n6791.n2558 vss 0.058178f
C7143 w_4660_n6791.n2559 vss 0.008764f
C7144 w_4660_n6791.n2560 vss 0.008764f
C7145 w_4660_n6791.n2561 vss 0.008764f
C7146 w_4660_n6791.n2562 vss 0.047437f
C7147 w_4660_n6791.n2563 vss 0.008764f
C7148 w_4660_n6791.n2564 vss 0.008764f
C7149 w_4660_n6791.n2565 vss 0.049227f
C7150 w_4660_n6791.n2566 vss 0.008764f
C7151 w_4660_n6791.n2567 vss 0.008764f
C7152 w_4660_n6791.n2568 vss 0.008764f
C7153 w_4660_n6791.n2569 vss 0.056388f
C7154 w_4660_n6791.n2570 vss 0.008764f
C7155 w_4660_n6791.n2571 vss 0.008764f
C7156 w_4660_n6791.n2572 vss 0.008764f
C7157 w_4660_n6791.n2573 vss 0.064443f
C7158 w_4660_n6791.n2574 vss 0.008764f
C7159 w_4660_n6791.n2575 vss 0.008764f
C7160 w_4660_n6791.n2576 vss 0.008764f
C7161 w_4660_n6791.n2577 vss 0.008764f
C7162 w_4660_n6791.n2578 vss 0.008764f
C7163 w_4660_n6791.n2579 vss 0.063548f
C7164 w_4660_n6791.n2580 vss 0.008764f
C7165 w_4660_n6791.n2581 vss 0.008764f
C7166 w_4660_n6791.n2582 vss 0.008764f
C7167 w_4660_n6791.n2583 vss 0.042067f
C7168 w_4660_n6791.n2584 vss 0.008764f
C7169 w_4660_n6791.n2585 vss 0.008764f
C7170 w_4660_n6791.n2586 vss 0.054598f
C7171 w_4660_n6791.n2587 vss 0.008764f
C7172 w_4660_n6791.n2588 vss 0.008764f
C7173 w_4660_n6791.n2589 vss 0.008764f
C7174 w_4660_n6791.n2590 vss 0.051017f
C7175 w_4660_n6791.n2591 vss 0.008764f
C7176 w_4660_n6791.n2592 vss 0.008764f
C7177 w_4660_n6791.n2593 vss 0.045647f
C7178 w_4660_n6791.n2594 vss 0.008764f
C7179 w_4660_n6791.n2595 vss 0.008764f
C7180 w_4660_n6791.n2596 vss 0.008764f
C7181 w_4660_n6791.n2597 vss 0.059968f
C7182 w_4660_n6791.n2598 vss 0.008764f
C7183 w_4660_n6791.n2599 vss 0.008764f
C7184 w_4660_n6791.n2600 vss 0.036697f
C7185 w_4660_n6791.n2601 vss 0.008764f
C7186 w_4660_n6791.n2602 vss 0.008764f
C7187 w_4660_n6791.n2603 vss 0.008764f
C7188 w_4660_n6791.n2604 vss 0.008764f
C7189 w_4660_n6791.n2605 vss 0.064443f
C7190 w_4660_n6791.n2606 vss 0.008764f
C7191 w_4660_n6791.n2607 vss 0.008764f
C7192 w_4660_n6791.n2608 vss 0.008764f
C7193 w_4660_n6791.n2609 vss 0.008764f
C7194 w_4660_n6791.n2610 vss 0.008764f
C7195 w_4660_n6791.n2611 vss 0.059968f
C7196 w_4660_n6791.n2612 vss 0.032221f
C7197 w_4660_n6791.n2613 vss 0.90734f
C7198 w_4660_n6791.n2614 vss 0.884154f
C7199 w_4660_n6791.n2615 vss 0.032221f
C7200 w_4660_n6791.n2616 vss 0.051465f
C7201 w_4660_n6791.n2617 vss 0.008825f
C7202 w_4660_n6791.n2618 vss 0.008825f
C7203 w_4660_n6791.n2619 vss 0.003287f
C7204 w_4660_n6791.n2620 vss 0.013195f
C7205 w_4660_n6791.n2621 vss 0.001438f
C7206 w_4660_n6791.n2622 vss 0.010797f
C7207 w_4660_n6791.n2623 vss 0.008582f
C7208 w_4660_n6791.n2624 vss 0.009022f
C7209 w_4660_n6791.n2625 vss 0.061865f
C7210 w_4660_n6791.n2626 vss 0.008764f
C7211 w_4660_n6791.n2627 vss 0.008764f
C7212 w_4660_n6791.n2628 vss 0.008764f
C7213 w_4660_n6791.n2629 vss 0.061865f
C7214 w_4660_n6791.n2630 vss 0.009022f
C7215 w_4660_n6791.n2631 vss 0.009022f
C7216 w_4660_n6791.n2632 vss 0.009022f
C7217 w_4660_n6791.n2633 vss 0.061865f
C7218 w_4660_n6791.n2634 vss 0.008764f
C7219 w_4660_n6791.n2635 vss 0.008764f
C7220 w_4660_n6791.n2636 vss 0.008764f
C7221 w_4660_n6791.n2637 vss 0.061865f
C7222 w_4660_n6791.n2638 vss 0.009022f
C7223 w_4660_n6791.n2639 vss 0.009022f
C7224 w_4660_n6791.n2640 vss 0.009022f
C7225 w_4660_n6791.n2641 vss 0.061865f
C7226 w_4660_n6791.n2642 vss 0.008764f
C7227 w_4660_n6791.n2643 vss 0.008764f
C7228 w_4660_n6791.n2644 vss 0.008764f
C7229 w_4660_n6791.n2645 vss 0.061865f
C7230 w_4660_n6791.n2646 vss 0.006201f
C7231 w_4660_n6791.n2647 vss 0.004507f
C7232 w_4660_n6791.n2648 vss 0.48173f
C7233 w_4660_n6791.n2649 vss 4.17527f
C7234 w_4660_n6791.n2650 vss 0.48173f
C7235 w_4660_n6791.n2651 vss 0.004507f
C7236 w_4660_n6791.n2652 vss 0.007579f
C7237 w_4660_n6791.n2653 vss 0.061865f
C7238 w_4660_n6791.n2654 vss 0.008764f
C7239 w_4660_n6791.n2655 vss 0.008764f
C7240 w_4660_n6791.n2656 vss 0.008764f
C7241 w_4660_n6791.n2657 vss 0.061865f
C7242 w_4660_n6791.n2658 vss 0.009022f
C7243 w_4660_n6791.n2659 vss 0.009022f
C7244 w_4660_n6791.n2660 vss 0.009022f
C7245 w_4660_n6791.n2661 vss 0.061865f
C7246 w_4660_n6791.n2662 vss 0.008764f
C7247 w_4660_n6791.n2663 vss 0.008764f
C7248 w_4660_n6791.n2664 vss 0.008764f
C7249 w_4660_n6791.n2665 vss 0.061865f
C7250 w_4660_n6791.n2666 vss 0.009022f
C7251 w_4660_n6791.n2667 vss 0.009022f
C7252 w_4660_n6791.n2668 vss 0.009022f
C7253 w_4660_n6791.n2669 vss 0.061865f
C7254 w_4660_n6791.n2670 vss 0.008764f
C7255 w_4660_n6791.n2671 vss 0.008764f
C7256 w_4660_n6791.n2672 vss 0.008764f
C7257 w_4660_n6791.n2673 vss 0.061865f
C7258 w_4660_n6791.n2674 vss 0.051499f
C7259 w_4660_n6791.n2675 vss 0.007203f
C7260 w_4660_n6791.n2676 vss 0.007858f
C7261 w_4660_n6791.n2677 vss 0.004325f
C7262 w_4660_n6791.n2678 vss 0.044892f
C7263 w_4660_n6791.n2679 vss 0.008764f
C7264 w_4660_n6791.n2680 vss 0.008764f
C7265 w_4660_n6791.n2681 vss 0.008764f
C7266 w_4660_n6791.n2682 vss 0.010263f
C7267 w_4660_n6791.n2683 vss 0.045647f
C7268 w_4660_n6791.n2684 vss 0.008764f
C7269 w_4660_n6791.n2685 vss 0.008764f
C7270 w_4660_n6791.n2686 vss 0.008764f
C7271 w_4660_n6791.n2687 vss 0.059968f
C7272 w_4660_n6791.n2688 vss 0.008764f
C7273 w_4660_n6791.n2689 vss 0.008764f
C7274 w_4660_n6791.n2690 vss 0.008764f
C7275 w_4660_n6791.n2691 vss 0.064443f
C7276 w_4660_n6791.n2692 vss 0.008764f
C7277 w_4660_n6791.n2693 vss 0.008764f
C7278 w_4660_n6791.n2694 vss 0.008764f
C7279 w_4660_n6791.n2695 vss 0.036697f
C7280 w_4660_n6791.n2696 vss 0.032221f
C7281 w_4660_n6791.n2697 vss 0.390261f
C7282 w_4660_n6791.n2698 vss 0.045937f
C7283 w_4660_n6791.n2699 vss 0.081778f
C7284 w_4660_n6791.n2700 vss 0.081778f
C7285 w_4660_n6791.n2701 vss 0.383942f
C7286 w_4660_n6791.n2702 vss 0.082195f
C7287 w_4660_n6791.n2703 vss 0.46332f
C7288 w_4660_n6791.n2704 vss 0.069153f
C7289 w_4660_n6791.t388 vss 0.031147f
C7290 vbn.n0 vss 0.384278f
C7291 vbn.n1 vss 0.384278f
C7292 vbn.n2 vss 0.384278f
C7293 vbn.n3 vss 0.384278f
C7294 vbn.n4 vss 0.384278f
C7295 vbn.n5 vss 24.1002f
C7296 vbn.n7 vss 2.46247f
C7297 vbn.n9 vss 2.46247f
C7298 vbn.n11 vss 2.46247f
C7299 vbn.n13 vss 2.46247f
C7300 vbn.n14 vss 1.4833f
C7301 vbn.n15 vss 1.64165f
C7302 vbn.n16 vss 1.64165f
C7303 vbn.n17 vss 1.64165f
C7304 vbn.n18 vss 1.64165f
C7305 vbn.n19 vss 1.64165f
C7306 vbn.n20 vss 1.64165f
C7307 vbn.n22 vss 1.64165f
C7308 vbn.n23 vss 1.64165f
C7309 vbn.n24 vss 1.64165f
C7310 vbn.n26 vss 1.4833f
C7311 vbn.n27 vss 1.64141f
C7312 vbn.n28 vss 1.64165f
C7313 vbn.n29 vss 1.64116f
C7314 vbn.n30 vss 1.64141f
C7315 vbn.n31 vss 1.64165f
C7316 vbn.n32 vss 1.64165f
C7317 vbn.n34 vss 1.64165f
C7318 vbn.n35 vss 1.64165f
C7319 vbn.n36 vss 1.64165f
C7320 vbn.n38 vss 1.4833f
C7321 vbn.n39 vss 1.64165f
C7322 vbn.n40 vss 1.64165f
C7323 vbn.n41 vss 1.64165f
C7324 vbn.n42 vss 1.64165f
C7325 vbn.n43 vss 1.64165f
C7326 vbn.n44 vss 1.64165f
C7327 vbn.n46 vss 1.64165f
C7328 vbn.n47 vss 1.64165f
C7329 vbn.n48 vss 1.64165f
C7330 vbn.n50 vss 1.4833f
C7331 vbn.n51 vss 1.64141f
C7332 vbn.n52 vss 1.64165f
C7333 vbn.n53 vss 1.64116f
C7334 vbn.n54 vss 1.64141f
C7335 vbn.n55 vss 1.64165f
C7336 vbn.n56 vss 1.64165f
C7337 vbn.n58 vss 1.64165f
C7338 vbn.n59 vss 1.64165f
C7339 vbn.n60 vss 1.64165f
C7340 vbn.n62 vss 17.8336f
C7341 vbn.n63 vss 32.658802f
C7342 vbn.n64 vss 1.48338f
C7343 vbn.n65 vss 1.48338f
C7344 vbn.n66 vss 1.48338f
C7345 vbn.n67 vss 1.48338f
C7346 vbn.t277 vss 0.098636f
C7347 vbn.t283 vss 0.098636f
C7348 vbn.n68 vss 0.098173f
C7349 vbn.t275 vss 0.098636f
C7350 vbn.t282 vss 0.098636f
C7351 vbn.n69 vss 0.097984f
C7352 vbn.n70 vss 0.282123f
C7353 vbn.t273 vss 0.098636f
C7354 vbn.t281 vss 0.098636f
C7355 vbn.n71 vss 0.097984f
C7356 vbn.n72 vss 0.132261f
C7357 vbn.t270 vss 0.098636f
C7358 vbn.t280 vss 0.098636f
C7359 vbn.n73 vss 0.097984f
C7360 vbn.n74 vss 0.132261f
C7361 vbn.t263 vss 0.098636f
C7362 vbn.t272 vss 0.098636f
C7363 vbn.n75 vss 0.097984f
C7364 vbn.n76 vss 0.132261f
C7365 vbn.t288 vss 0.098636f
C7366 vbn.t267 vss 0.098636f
C7367 vbn.n77 vss 0.097984f
C7368 vbn.n78 vss 0.132261f
C7369 vbn.t287 vss 0.098636f
C7370 vbn.t265 vss 0.098636f
C7371 vbn.n79 vss 0.097984f
C7372 vbn.n80 vss 0.132261f
C7373 vbn.t286 vss 0.098636f
C7374 vbn.t262 vss 0.098636f
C7375 vbn.n81 vss 0.097984f
C7376 vbn.n82 vss 0.132261f
C7377 vbn.t284 vss 0.098636f
C7378 vbn.t260 vss 0.098636f
C7379 vbn.n83 vss 0.097984f
C7380 vbn.n84 vss 0.132261f
C7381 vbn.t279 vss 0.098636f
C7382 vbn.t285 vss 0.098636f
C7383 vbn.n85 vss 0.097984f
C7384 vbn.n86 vss 0.132261f
C7385 vbn.t268 vss 0.098636f
C7386 vbn.t278 vss 0.098636f
C7387 vbn.n87 vss 0.097984f
C7388 vbn.n88 vss 0.132261f
C7389 vbn.t266 vss 0.098636f
C7390 vbn.t276 vss 0.098636f
C7391 vbn.n89 vss 0.097984f
C7392 vbn.n90 vss 0.132261f
C7393 vbn.t264 vss 0.098636f
C7394 vbn.t274 vss 0.098636f
C7395 vbn.n91 vss 0.097984f
C7396 vbn.n92 vss 0.132261f
C7397 vbn.t261 vss 0.098636f
C7398 vbn.t271 vss 0.098636f
C7399 vbn.n93 vss 0.097984f
C7400 vbn.n94 vss 0.132261f
C7401 vbn.t289 vss 0.098636f
C7402 vbn.t269 vss 0.098636f
C7403 vbn.n95 vss 0.097984f
C7404 vbn.n96 vss 0.185948f
C7405 vbn.n97 vss 0.175755f
C7406 vbn.t11 vss 0.031767f
C7407 vbn.t17 vss 0.031767f
C7408 vbn.n98 vss 0.071954f
C7409 vbn.t16 vss 0.098636f
C7410 vbn.t58 vss 0.098636f
C7411 vbn.n99 vss 0.097984f
C7412 vbn.n100 vss 0.113519f
C7413 vbn.t7 vss 0.11586f
C7414 vbn.n101 vss 0.443563f
C7415 vbn.t55 vss 0.11586f
C7416 vbn.n102 vss 0.443475f
C7417 vbn.t13 vss 0.031767f
C7418 vbn.t19 vss 0.031767f
C7419 vbn.n103 vss 0.071954f
C7420 vbn.n104 vss 0.384278f
C7421 vbn.t39 vss 0.031767f
C7422 vbn.t49 vss 0.031767f
C7423 vbn.n105 vss 0.071954f
C7424 vbn.n106 vss 0.384278f
C7425 vbn.t9 vss 0.031767f
C7426 vbn.t15 vss 0.031767f
C7427 vbn.n107 vss 0.071954f
C7428 vbn.n108 vss 0.384278f
C7429 vbn.t29 vss 0.031767f
C7430 vbn.t21 vss 0.031767f
C7431 vbn.n109 vss 0.071954f
C7432 vbn.n110 vss 0.384278f
C7433 vbn.t53 vss 0.031767f
C7434 vbn.t5 vss 0.031767f
C7435 vbn.n111 vss 0.071954f
C7436 vbn.n112 vss 0.384278f
C7437 vbn.t43 vss 0.031767f
C7438 vbn.t47 vss 0.031767f
C7439 vbn.n113 vss 0.071954f
C7440 vbn.t42 vss 0.098636f
C7441 vbn.t24 vss 0.098636f
C7442 vbn.n114 vss 0.097984f
C7443 vbn.n115 vss 0.113519f
C7444 vbn.t51 vss 0.031767f
C7445 vbn.t1 vss 0.031767f
C7446 vbn.n116 vss 0.071954f
C7447 vbn.t3 vss 0.031767f
C7448 vbn.t23 vss 0.031767f
C7449 vbn.n117 vss 0.071954f
C7450 vbn.t27 vss 0.031767f
C7451 vbn.t35 vss 0.031767f
C7452 vbn.n118 vss 0.071954f
C7453 vbn.t120 vss 0.031767f
C7454 vbn.t213 vss 0.031767f
C7455 vbn.n119 vss 0.068563f
C7456 vbn.t257 vss 0.031767f
C7457 vbn.t75 vss 0.031767f
C7458 vbn.n120 vss 0.068475f
C7459 vbn.t92 vss 0.031767f
C7460 vbn.t200 vss 0.031767f
C7461 vbn.n121 vss 0.068475f
C7462 vbn.t217 vss 0.031767f
C7463 vbn.t133 vss 0.031767f
C7464 vbn.n122 vss 0.068475f
C7465 vbn.t123 vss 0.031767f
C7466 vbn.t115 vss 0.031767f
C7467 vbn.n123 vss 0.068475f
C7468 vbn.t111 vss 0.031767f
C7469 vbn.t247 vss 0.031767f
C7470 vbn.n124 vss 0.068475f
C7471 vbn.t128 vss 0.031767f
C7472 vbn.t186 vss 0.031767f
C7473 vbn.n125 vss 0.068475f
C7474 vbn.t164 vss 0.031767f
C7475 vbn.t227 vss 0.031767f
C7476 vbn.n126 vss 0.068475f
C7477 vbn.t121 vss 0.031767f
C7478 vbn.t114 vss 0.031767f
C7479 vbn.n127 vss 0.068475f
C7480 vbn.t156 vss 0.031767f
C7481 vbn.t245 vss 0.031767f
C7482 vbn.n128 vss 0.068475f
C7483 vbn.t214 vss 0.031767f
C7484 vbn.t77 vss 0.031767f
C7485 vbn.n129 vss 0.068475f
C7486 vbn.t249 vss 0.031767f
C7487 vbn.t256 vss 0.031767f
C7488 vbn.n130 vss 0.068646f
C7489 vbn.t208 vss 0.031767f
C7490 vbn.t104 vss 0.031767f
C7491 vbn.n131 vss 0.068475f
C7492 vbn.t73 vss 0.031767f
C7493 vbn.t91 vss 0.031767f
C7494 vbn.n132 vss 0.068475f
C7495 vbn.t234 vss 0.031767f
C7496 vbn.t210 vss 0.031767f
C7497 vbn.n133 vss 0.068475f
C7498 vbn.t212 vss 0.031767f
C7499 vbn.t105 vss 0.031767f
C7500 vbn.n134 vss 0.068475f
C7501 vbn.t99 vss 0.031767f
C7502 vbn.t232 vss 0.031767f
C7503 vbn.n135 vss 0.068475f
C7504 vbn.t94 vss 0.031767f
C7505 vbn.t84 vss 0.031767f
C7506 vbn.n136 vss 0.068475f
C7507 vbn.t87 vss 0.031767f
C7508 vbn.t64 vss 0.031767f
C7509 vbn.n137 vss 0.068475f
C7510 vbn.t189 vss 0.031767f
C7511 vbn.t185 vss 0.031767f
C7512 vbn.n138 vss 0.068475f
C7513 vbn.t144 vss 0.031767f
C7514 vbn.t135 vss 0.031767f
C7515 vbn.n139 vss 0.068475f
C7516 vbn.t182 vss 0.031767f
C7517 vbn.t85 vss 0.031767f
C7518 vbn.n140 vss 0.068475f
C7519 vbn.t86 vss 0.031767f
C7520 vbn.t242 vss 0.031767f
C7521 vbn.n141 vss 0.068475f
C7522 vbn.t127 vss 0.031767f
C7523 vbn.t196 vss 0.031767f
C7524 vbn.n142 vss 0.068475f
C7525 vbn.t145 vss 0.031767f
C7526 vbn.t221 vss 0.031767f
C7527 vbn.n143 vss 0.068475f
C7528 vbn.t224 vss 0.031767f
C7529 vbn.t103 vss 0.031767f
C7530 vbn.n144 vss 0.068563f
C7531 vbn.t226 vss 0.031767f
C7532 vbn.t151 vss 0.031767f
C7533 vbn.n145 vss 0.068475f
C7534 vbn.t177 vss 0.031767f
C7535 vbn.t109 vss 0.031767f
C7536 vbn.n146 vss 0.068475f
C7537 vbn.t173 vss 0.031767f
C7538 vbn.t229 vss 0.031767f
C7539 vbn.n147 vss 0.068475f
C7540 vbn.t149 vss 0.031767f
C7541 vbn.t241 vss 0.031767f
C7542 vbn.n148 vss 0.068475f
C7543 vbn.t236 vss 0.031767f
C7544 vbn.t130 vss 0.031767f
C7545 vbn.n149 vss 0.068475f
C7546 vbn.t66 vss 0.031767f
C7547 vbn.t238 vss 0.031767f
C7548 vbn.n150 vss 0.068475f
C7549 vbn.t246 vss 0.031767f
C7550 vbn.t199 vss 0.031767f
C7551 vbn.n151 vss 0.068475f
C7552 vbn.t167 vss 0.031767f
C7553 vbn.t170 vss 0.031767f
C7554 vbn.n152 vss 0.068475f
C7555 vbn.t143 vss 0.031767f
C7556 vbn.t155 vss 0.031767f
C7557 vbn.n153 vss 0.068475f
C7558 vbn.t134 vss 0.031767f
C7559 vbn.t166 vss 0.031767f
C7560 vbn.n154 vss 0.068475f
C7561 vbn.t74 vss 0.031767f
C7562 vbn.t132 vss 0.031767f
C7563 vbn.n155 vss 0.068646f
C7564 vbn.t206 vss 0.031767f
C7565 vbn.t122 vss 0.031767f
C7566 vbn.n156 vss 0.068475f
C7567 vbn.t258 vss 0.031767f
C7568 vbn.t78 vss 0.031767f
C7569 vbn.n157 vss 0.068475f
C7570 vbn.t131 vss 0.031767f
C7571 vbn.t154 vss 0.031767f
C7572 vbn.n158 vss 0.068475f
C7573 vbn.t174 vss 0.031767f
C7574 vbn.t223 vss 0.031767f
C7575 vbn.n159 vss 0.068475f
C7576 vbn.t162 vss 0.031767f
C7577 vbn.t63 vss 0.031767f
C7578 vbn.n160 vss 0.068475f
C7579 vbn.t231 vss 0.031767f
C7580 vbn.t218 vss 0.031767f
C7581 vbn.n161 vss 0.068475f
C7582 vbn.t116 vss 0.031767f
C7583 vbn.t71 vss 0.031767f
C7584 vbn.n162 vss 0.068475f
C7585 vbn.t159 vss 0.031767f
C7586 vbn.t207 vss 0.031767f
C7587 vbn.n163 vss 0.068475f
C7588 vbn.t139 vss 0.031767f
C7589 vbn.t259 vss 0.031767f
C7590 vbn.n164 vss 0.068475f
C7591 vbn.t89 vss 0.031767f
C7592 vbn.t255 vss 0.031767f
C7593 vbn.n165 vss 0.068475f
C7594 vbn.t183 vss 0.031767f
C7595 vbn.t184 vss 0.031767f
C7596 vbn.n166 vss 0.068475f
C7597 vbn.t219 vss 0.031767f
C7598 vbn.t98 vss 0.031767f
C7599 vbn.n167 vss 0.068475f
C7600 vbn.t233 vss 0.031767f
C7601 vbn.t204 vss 0.031767f
C7602 vbn.n168 vss 0.068475f
C7603 vbn.t136 vss 0.031767f
C7604 vbn.t230 vss 0.031767f
C7605 vbn.n169 vss 0.068563f
C7606 vbn.t150 vss 0.031767f
C7607 vbn.t117 vss 0.031767f
C7608 vbn.n170 vss 0.068475f
C7609 vbn.t220 vss 0.031767f
C7610 vbn.t202 vss 0.031767f
C7611 vbn.n171 vss 0.068475f
C7612 vbn.t168 vss 0.031767f
C7613 vbn.t197 vss 0.031767f
C7614 vbn.n172 vss 0.068475f
C7615 vbn.t209 vss 0.031767f
C7616 vbn.t169 vss 0.031767f
C7617 vbn.n173 vss 0.068475f
C7618 vbn.t228 vss 0.031767f
C7619 vbn.t180 vss 0.031767f
C7620 vbn.n174 vss 0.068475f
C7621 vbn.t175 vss 0.031767f
C7622 vbn.t93 vss 0.031767f
C7623 vbn.n175 vss 0.068475f
C7624 vbn.t76 vss 0.031767f
C7625 vbn.t72 vss 0.031767f
C7626 vbn.n176 vss 0.068475f
C7627 vbn.t100 vss 0.031767f
C7628 vbn.t152 vss 0.031767f
C7629 vbn.n177 vss 0.068475f
C7630 vbn.t193 vss 0.031767f
C7631 vbn.t110 vss 0.031767f
C7632 vbn.n178 vss 0.068475f
C7633 vbn.t124 vss 0.031767f
C7634 vbn.t201 vss 0.031767f
C7635 vbn.n179 vss 0.068475f
C7636 vbn.t141 vss 0.031767f
C7637 vbn.t147 vss 0.031767f
C7638 vbn.n180 vss 0.068646f
C7639 vbn.t187 vss 0.031767f
C7640 vbn.t160 vss 0.031767f
C7641 vbn.n181 vss 0.068475f
C7642 vbn.t235 vss 0.031767f
C7643 vbn.t237 vss 0.031767f
C7644 vbn.n182 vss 0.068475f
C7645 vbn.t161 vss 0.031767f
C7646 vbn.t81 vss 0.031767f
C7647 vbn.n183 vss 0.068475f
C7648 vbn.t106 vss 0.031767f
C7649 vbn.t61 vss 0.031767f
C7650 vbn.n184 vss 0.068475f
C7651 vbn.t65 vss 0.031767f
C7652 vbn.t253 vss 0.031767f
C7653 vbn.n185 vss 0.068475f
C7654 vbn.t243 vss 0.031767f
C7655 vbn.t82 vss 0.031767f
C7656 vbn.n186 vss 0.068475f
C7657 vbn.t69 vss 0.031767f
C7658 vbn.t79 vss 0.031767f
C7659 vbn.n187 vss 0.068475f
C7660 vbn.t203 vss 0.031767f
C7661 vbn.t129 vss 0.031767f
C7662 vbn.n188 vss 0.068475f
C7663 vbn.t108 vss 0.031767f
C7664 vbn.t251 vss 0.031767f
C7665 vbn.n189 vss 0.068475f
C7666 vbn.t216 vss 0.031767f
C7667 vbn.t67 vss 0.031767f
C7668 vbn.n190 vss 0.068475f
C7669 vbn.t163 vss 0.031767f
C7670 vbn.t178 vss 0.031767f
C7671 vbn.n191 vss 0.068475f
C7672 vbn.t138 vss 0.031767f
C7673 vbn.t190 vss 0.031767f
C7674 vbn.n192 vss 0.068475f
C7675 vbn.t248 vss 0.031767f
C7676 vbn.t88 vss 0.031767f
C7677 vbn.n193 vss 0.068475f
C7678 vbn.t137 vss 0.031767f
C7679 vbn.t195 vss 0.031767f
C7680 vbn.n194 vss 0.068563f
C7681 vbn.t113 vss 0.031767f
C7682 vbn.t118 vss 0.031767f
C7683 vbn.n195 vss 0.068475f
C7684 vbn.t165 vss 0.031767f
C7685 vbn.t240 vss 0.031767f
C7686 vbn.n196 vss 0.068475f
C7687 vbn.t225 vss 0.031767f
C7688 vbn.t198 vss 0.031767f
C7689 vbn.n197 vss 0.068475f
C7690 vbn.t211 vss 0.031767f
C7691 vbn.t171 vss 0.031767f
C7692 vbn.n198 vss 0.068475f
C7693 vbn.t179 vss 0.031767f
C7694 vbn.t181 vss 0.031767f
C7695 vbn.n199 vss 0.068475f
C7696 vbn.t176 vss 0.031767f
C7697 vbn.t96 vss 0.031767f
C7698 vbn.n200 vss 0.068475f
C7699 vbn.t70 vss 0.031767f
C7700 vbn.t97 vss 0.031767f
C7701 vbn.n201 vss 0.068475f
C7702 vbn.t146 vss 0.031767f
C7703 vbn.t153 vss 0.031767f
C7704 vbn.n202 vss 0.068475f
C7705 vbn.t194 vss 0.031767f
C7706 vbn.t112 vss 0.031767f
C7707 vbn.n203 vss 0.068475f
C7708 vbn.t126 vss 0.031767f
C7709 vbn.t239 vss 0.031767f
C7710 vbn.n204 vss 0.068475f
C7711 vbn.t142 vss 0.031767f
C7712 vbn.t148 vss 0.031767f
C7713 vbn.n205 vss 0.068646f
C7714 vbn.t188 vss 0.031767f
C7715 vbn.t192 vss 0.031767f
C7716 vbn.n206 vss 0.068475f
C7717 vbn.t157 vss 0.031767f
C7718 vbn.t172 vss 0.031767f
C7719 vbn.n207 vss 0.068475f
C7720 vbn.t101 vss 0.031767f
C7721 vbn.t90 vss 0.031767f
C7722 vbn.n208 vss 0.068475f
C7723 vbn.t60 vss 0.031767f
C7724 vbn.t62 vss 0.031767f
C7725 vbn.n209 vss 0.068475f
C7726 vbn.t254 vss 0.031767f
C7727 vbn.t215 vss 0.031767f
C7728 vbn.n210 vss 0.068475f
C7729 vbn.t244 vss 0.031767f
C7730 vbn.t83 vss 0.031767f
C7731 vbn.n211 vss 0.068475f
C7732 vbn.t125 vss 0.031767f
C7733 vbn.t80 vss 0.031767f
C7734 vbn.n212 vss 0.068475f
C7735 vbn.t205 vss 0.031767f
C7736 vbn.t107 vss 0.031767f
C7737 vbn.n213 vss 0.068475f
C7738 vbn.t222 vss 0.031767f
C7739 vbn.t252 vss 0.031767f
C7740 vbn.n214 vss 0.068475f
C7741 vbn.t119 vss 0.031767f
C7742 vbn.t68 vss 0.031767f
C7743 vbn.n215 vss 0.068475f
C7744 vbn.t102 vss 0.031767f
C7745 vbn.t95 vss 0.031767f
C7746 vbn.n216 vss 0.068475f
C7747 vbn.t140 vss 0.031767f
C7748 vbn.t191 vss 0.031767f
C7749 vbn.n217 vss 0.068475f
C7750 vbn.t250 vss 0.031767f
C7751 vbn.t158 vss 0.031767f
C7752 vbn.n218 vss 0.068475f
C7753 vbn.t31 vss 0.031767f
C7754 vbn.t37 vss 0.031767f
C7755 vbn.n219 vss 0.071954f
C7756 vbn.t30 vss 0.098636f
C7757 vbn.t12 vss 0.098636f
C7758 vbn.n220 vss 0.097984f
C7759 vbn.n221 vss 0.113519f
C7760 vbn.t36 vss 0.098636f
C7761 vbn.t18 vss 0.098636f
C7762 vbn.n222 vss 0.097984f
C7763 vbn.n223 vss 0.113519f
C7764 vbn.n224 vss 0.103327f
C7765 vbn.n225 vss 0.384278f
C7766 vbn.t45 vss 0.031767f
C7767 vbn.t41 vss 0.031767f
C7768 vbn.n226 vss 0.071954f
C7769 vbn.n227 vss 0.384278f
C7770 vbn.t40 vss 0.098636f
C7771 vbn.t20 vss 0.098636f
C7772 vbn.n228 vss 0.098044f
C7773 vbn.n229 vss 0.197726f
C7774 vbn.t44 vss 0.098636f
C7775 vbn.t28 vss 0.098636f
C7776 vbn.n230 vss 0.097984f
C7777 vbn.n231 vss 0.113519f
C7778 vbn.t34 vss 0.098636f
C7779 vbn.t14 vss 0.098636f
C7780 vbn.n232 vss 0.097984f
C7781 vbn.n233 vss 0.113519f
C7782 vbn.n234 vss 0.103327f
C7783 vbn.t26 vss 0.098636f
C7784 vbn.t8 vss 0.098636f
C7785 vbn.n235 vss 0.097984f
C7786 vbn.n236 vss 0.113519f
C7787 vbn.t22 vss 0.098636f
C7788 vbn.t4 vss 0.098636f
C7789 vbn.n237 vss 0.097984f
C7790 vbn.n238 vss 0.113519f
C7791 vbn.n239 vss 0.103327f
C7792 vbn.t2 vss 0.098636f
C7793 vbn.t52 vss 0.098636f
C7794 vbn.n240 vss 0.097984f
C7795 vbn.n241 vss 0.113519f
C7796 vbn.t0 vss 0.098636f
C7797 vbn.t48 vss 0.098636f
C7798 vbn.n242 vss 0.097984f
C7799 vbn.n243 vss 0.113519f
C7800 vbn.n244 vss 0.103327f
C7801 vbn.t50 vss 0.098636f
C7802 vbn.t38 vss 0.098636f
C7803 vbn.n245 vss 0.097984f
C7804 vbn.n246 vss 0.113519f
C7805 vbn.t46 vss 0.098636f
C7806 vbn.t32 vss 0.098636f
C7807 vbn.n247 vss 0.097984f
C7808 vbn.n248 vss 0.113519f
C7809 vbn.n249 vss 0.103327f
C7810 vbn.t25 vss 0.031767f
C7811 vbn.t33 vss 0.031767f
C7812 vbn.n250 vss 0.071954f
C7813 vbn.n251 vss 0.384278f
C7814 vbn.t57 vss 0.031767f
C7815 vbn.t59 vss 0.031767f
C7816 vbn.n252 vss 0.071954f
C7817 vbn.n253 vss 0.384278f
C7818 vbn.n254 vss 0.103327f
C7819 vbn.t10 vss 0.098636f
C7820 vbn.t56 vss 0.098636f
C7821 vbn.n255 vss 0.097984f
C7822 vbn.n256 vss 0.113519f
C7823 vbn.t6 vss 0.098636f
C7824 vbn.t54 vss 0.098636f
C7825 vbn.n257 vss 0.097984f
C7826 vbn.n258 vss 0.113519f
C7827 vin_n.t39 vss 0.128597f
C7828 vin_n.t114 vss 0.128597f
C7829 vin_n.n0 vss 0.126803f
C7830 vin_n.t62 vss 0.128597f
C7831 vin_n.t36 vss 0.128597f
C7832 vin_n.n1 vss 0.126618f
C7833 vin_n.n2 vss 0.303932f
C7834 vin_n.t92 vss 0.128597f
C7835 vin_n.t94 vss 0.128597f
C7836 vin_n.n3 vss 0.126618f
C7837 vin_n.n4 vss 0.163639f
C7838 vin_n.t73 vss 0.128597f
C7839 vin_n.t9 vss 0.128597f
C7840 vin_n.n5 vss 0.126618f
C7841 vin_n.n6 vss 0.163639f
C7842 vin_n.t107 vss 0.128597f
C7843 vin_n.t75 vss 0.128597f
C7844 vin_n.n7 vss 0.126618f
C7845 vin_n.n8 vss 0.163639f
C7846 vin_n.t140 vss 0.128597f
C7847 vin_n.t146 vss 0.128597f
C7848 vin_n.n9 vss 0.126618f
C7849 vin_n.n10 vss 0.163639f
C7850 vin_n.t24 vss 0.128597f
C7851 vin_n.t37 vss 0.128597f
C7852 vin_n.n11 vss 0.126618f
C7853 vin_n.n12 vss 0.163639f
C7854 vin_n.t60 vss 0.128597f
C7855 vin_n.t97 vss 0.128597f
C7856 vin_n.n13 vss 0.126618f
C7857 vin_n.n14 vss 0.163639f
C7858 vin_n.t43 vss 0.128597f
C7859 vin_n.t11 vss 0.128597f
C7860 vin_n.n15 vss 0.126618f
C7861 vin_n.n16 vss 0.163639f
C7862 vin_n.t72 vss 0.128597f
C7863 vin_n.t78 vss 0.128597f
C7864 vin_n.n17 vss 0.126618f
C7865 vin_n.n18 vss 0.163639f
C7866 vin_n.t104 vss 0.128597f
C7867 vin_n.t152 vss 0.128597f
C7868 vin_n.n19 vss 0.126618f
C7869 vin_n.n20 vss 0.163639f
C7870 vin_n.t131 vss 0.128597f
C7871 vin_n.t67 vss 0.128597f
C7872 vin_n.n21 vss 0.126618f
C7873 vin_n.n22 vss 0.163639f
C7874 vin_n.t172 vss 0.128597f
C7875 vin_n.t132 vss 0.128597f
C7876 vin_n.n23 vss 0.126618f
C7877 vin_n.n24 vss 0.163639f
C7878 vin_n.t195 vss 0.128597f
C7879 vin_n.t193 vss 0.128597f
C7880 vin_n.n25 vss 0.126618f
C7881 vin_n.n26 vss 0.163639f
C7882 vin_n.t33 vss 0.128597f
C7883 vin_n.t46 vss 0.128597f
C7884 vin_n.n27 vss 0.126618f
C7885 vin_n.n28 vss 0.163639f
C7886 vin_n.t66 vss 0.128597f
C7887 vin_n.t109 vss 0.128597f
C7888 vin_n.n29 vss 0.126618f
C7889 vin_n.n30 vss 0.163639f
C7890 vin_n.t88 vss 0.128597f
C7891 vin_n.t30 vss 0.128597f
C7892 vin_n.n31 vss 0.126618f
C7893 vin_n.n32 vss 0.163639f
C7894 vin_n.t124 vss 0.128597f
C7895 vin_n.t93 vss 0.128597f
C7896 vin_n.n33 vss 0.126618f
C7897 vin_n.n34 vss 0.163639f
C7898 vin_n.t163 vss 0.128597f
C7899 vin_n.t168 vss 0.128597f
C7900 vin_n.n35 vss 0.126618f
C7901 vin_n.n36 vss 0.163639f
C7902 vin_n.t137 vss 0.128597f
C7903 vin_n.t74 vss 0.128597f
C7904 vin_n.n37 vss 0.126618f
C7905 vin_n.n38 vss 0.163639f
C7906 vin_n.t178 vss 0.128597f
C7907 vin_n.t142 vss 0.128597f
C7908 vin_n.n39 vss 0.126618f
C7909 vin_n.n40 vss 0.163639f
C7910 vin_n.t194 vss 0.128597f
C7911 vin_n.t63 vss 0.128597f
C7912 vin_n.n41 vss 0.126618f
C7913 vin_n.n42 vss 0.163639f
C7914 vin_n.t34 vss 0.128597f
C7915 vin_n.t126 vss 0.128597f
C7916 vin_n.n43 vss 0.126618f
C7917 vin_n.n44 vss 0.163639f
C7918 vin_n.t115 vss 0.128597f
C7919 vin_n.t125 vss 0.128597f
C7920 vin_n.n45 vss 0.126618f
C7921 vin_n.n46 vss 0.163639f
C7922 vin_n.t154 vss 0.128597f
C7923 vin_n.t192 vss 0.128597f
C7924 vin_n.n47 vss 0.126618f
C7925 vin_n.n48 vss 0.163639f
C7926 vin_n.t129 vss 0.128597f
C7927 vin_n.t105 vss 0.128597f
C7928 vin_n.n49 vss 0.126618f
C7929 vin_n.n50 vss 0.163639f
C7930 vin_n.t162 vss 0.128597f
C7931 vin_n.t25 vss 0.128597f
C7932 vin_n.n51 vss 0.126618f
C7933 vin_n.n52 vss 0.163639f
C7934 vin_n.t190 vss 0.128597f
C7935 vin_n.t90 vss 0.128597f
C7936 vin_n.n53 vss 0.126618f
C7937 vin_n.n54 vss 0.163639f
C7938 vin_n.t21 vss 0.128597f
C7939 vin_n.t164 vss 0.128597f
C7940 vin_n.n55 vss 0.126618f
C7941 vin_n.n56 vss 0.163639f
C7942 vin_n.t58 vss 0.128597f
C7943 vin_n.t22 vss 0.128597f
C7944 vin_n.n57 vss 0.126618f
C7945 vin_n.n58 vss 0.163639f
C7946 vin_n.t41 vss 0.128597f
C7947 vin_n.t138 vss 0.128597f
C7948 vin_n.n59 vss 0.126618f
C7949 vin_n.n60 vss 0.163639f
C7950 vin_n.t111 vss 0.128597f
C7951 vin_n.t188 vss 0.128597f
C7952 vin_n.n61 vss 0.126618f
C7953 vin_n.n62 vss 0.163639f
C7954 vin_n.t150 vss 0.128597f
C7955 vin_n.t57 vss 0.128597f
C7956 vin_n.n63 vss 0.126618f
C7957 vin_n.n64 vss 0.163639f
C7958 vin_n.t183 vss 0.128597f
C7959 vin_n.t122 vss 0.128597f
C7960 vin_n.n65 vss 0.126618f
C7961 vin_n.n66 vss 0.163639f
C7962 vin_n.t10 vss 0.128597f
C7963 vin_n.t187 vss 0.128597f
C7964 vin_n.n67 vss 0.126618f
C7965 vin_n.n68 vss 0.163639f
C7966 vin_n.t48 vss 0.128597f
C7967 vin_n.t54 vss 0.128597f
C7968 vin_n.n69 vss 0.126618f
C7969 vin_n.n70 vss 0.163639f
C7970 vin_n.t18 vss 0.128597f
C7971 vin_n.t16 vss 0.128597f
C7972 vin_n.n71 vss 0.126618f
C7973 vin_n.n72 vss 0.163639f
C7974 vin_n.t56 vss 0.128597f
C7975 vin_n.t83 vss 0.128597f
C7976 vin_n.n73 vss 0.126618f
C7977 vin_n.n74 vss 0.163639f
C7978 vin_n.t85 vss 0.128597f
C7979 vin_n.t161 vss 0.128597f
C7980 vin_n.n75 vss 0.126618f
C7981 vin_n.n76 vss 0.163639f
C7982 vin_n.t123 vss 0.128597f
C7983 vin_n.t14 vss 0.128597f
C7984 vin_n.n77 vss 0.126618f
C7985 vin_n.n78 vss 0.163639f
C7986 vin_n.t2 vss 0.128597f
C7987 vin_n.t12 vss 0.128597f
C7988 vin_n.n79 vss 0.126618f
C7989 vin_n.n80 vss 0.163639f
C7990 vin_n.t35 vss 0.128597f
C7991 vin_n.t134 vss 0.128597f
C7992 vin_n.n81 vss 0.126618f
C7993 vin_n.n82 vss 0.163639f
C7994 vin_n.t8 vss 0.128597f
C7995 vin_n.t52 vss 0.128597f
C7996 vin_n.n83 vss 0.126618f
C7997 vin_n.n84 vss 0.163639f
C7998 vin_n.t47 vss 0.128597f
C7999 vin_n.t116 vss 0.128597f
C8000 vin_n.n85 vss 0.126618f
C8001 vin_n.n86 vss 0.163639f
C8002 vin_n.t76 vss 0.128597f
C8003 vin_n.t184 vss 0.128597f
C8004 vin_n.n87 vss 0.126618f
C8005 vin_n.n88 vss 0.163639f
C8006 vin_n.t113 vss 0.128597f
C8007 vin_n.t50 vss 0.128597f
C8008 vin_n.n89 vss 0.126618f
C8009 vin_n.n90 vss 0.163639f
C8010 vin_n.t139 vss 0.128597f
C8011 vin_n.t175 vss 0.128597f
C8012 vin_n.n91 vss 0.126618f
C8013 vin_n.n92 vss 0.163639f
C8014 vin_n.t121 vss 0.128597f
C8015 vin_n.t80 vss 0.128597f
C8016 vin_n.n93 vss 0.126618f
C8017 vin_n.n94 vss 0.163639f
C8018 vin_n.t0 vss 0.128597f
C8019 vin_n.t77 vss 0.128597f
C8020 vin_n.n95 vss 0.126618f
C8021 vin_n.n96 vss 0.163639f
C8022 vin_n.t42 vss 0.128597f
C8023 vin_n.t147 vss 0.128597f
C8024 vin_n.n97 vss 0.126618f
C8025 vin_n.n98 vss 0.730131f
C8026 vin_n.t166 vss 0.128597f
C8027 vin_n.t165 vss 0.128597f
C8028 vin_n.n99 vss 0.126803f
C8029 vin_n.t101 vss 0.128597f
C8030 vin_n.t100 vss 0.128597f
C8031 vin_n.n100 vss 0.126618f
C8032 vin_n.n101 vss 0.303932f
C8033 vin_n.t96 vss 0.128597f
C8034 vin_n.t95 vss 0.128597f
C8035 vin_n.n102 vss 0.126618f
C8036 vin_n.n103 vss 0.163639f
C8037 vin_n.t29 vss 0.128597f
C8038 vin_n.t28 vss 0.128597f
C8039 vin_n.n104 vss 0.126618f
C8040 vin_n.n105 vss 0.163639f
C8041 vin_n.t23 vss 0.128597f
C8042 vin_n.t20 vss 0.128597f
C8043 vin_n.n106 vss 0.126618f
C8044 vin_n.n107 vss 0.163639f
C8045 vin_n.t15 vss 0.128597f
C8046 vin_n.t13 vss 0.128597f
C8047 vin_n.n108 vss 0.126618f
C8048 vin_n.n109 vss 0.163639f
C8049 vin_n.t153 vss 0.128597f
C8050 vin_n.t149 vss 0.128597f
C8051 vin_n.n110 vss 0.126618f
C8052 vin_n.n111 vss 0.163639f
C8053 vin_n.t143 vss 0.128597f
C8054 vin_n.t141 vss 0.128597f
C8055 vin_n.n112 vss 0.126618f
C8056 vin_n.n113 vss 0.163639f
C8057 vin_n.t71 vss 0.128597f
C8058 vin_n.t70 vss 0.128597f
C8059 vin_n.n114 vss 0.126618f
C8060 vin_n.n115 vss 0.163639f
C8061 vin_n.t69 vss 0.128597f
C8062 vin_n.t68 vss 0.128597f
C8063 vin_n.n116 vss 0.126618f
C8064 vin_n.n117 vss 0.163639f
C8065 vin_n.t65 vss 0.128597f
C8066 vin_n.t64 vss 0.128597f
C8067 vin_n.n118 vss 0.126618f
C8068 vin_n.n119 vss 0.163639f
C8069 vin_n.t5 vss 0.128597f
C8070 vin_n.t4 vss 0.128597f
C8071 vin_n.n120 vss 0.126618f
C8072 vin_n.n121 vss 0.163639f
C8073 vin_n.t199 vss 0.128597f
C8074 vin_n.t198 vss 0.128597f
C8075 vin_n.n122 vss 0.126618f
C8076 vin_n.n123 vss 0.163639f
C8077 vin_n.t197 vss 0.128597f
C8078 vin_n.t196 vss 0.128597f
C8079 vin_n.n124 vss 0.126618f
C8080 vin_n.n125 vss 0.163639f
C8081 vin_n.t158 vss 0.128597f
C8082 vin_n.t156 vss 0.128597f
C8083 vin_n.n126 vss 0.126618f
C8084 vin_n.n127 vss 0.163639f
C8085 vin_n.t145 vss 0.128597f
C8086 vin_n.t144 vss 0.128597f
C8087 vin_n.n128 vss 0.126618f
C8088 vin_n.n129 vss 0.163639f
C8089 vin_n.t91 vss 0.128597f
C8090 vin_n.t89 vss 0.128597f
C8091 vin_n.n130 vss 0.126618f
C8092 vin_n.n131 vss 0.163639f
C8093 vin_n.t84 vss 0.128597f
C8094 vin_n.t82 vss 0.128597f
C8095 vin_n.n132 vss 0.126618f
C8096 vin_n.n133 vss 0.163639f
C8097 vin_n.t81 vss 0.128597f
C8098 vin_n.t79 vss 0.128597f
C8099 vin_n.n134 vss 0.126618f
C8100 vin_n.n135 vss 0.163639f
C8101 vin_n.t7 vss 0.128597f
C8102 vin_n.t6 vss 0.128597f
C8103 vin_n.n136 vss 0.126618f
C8104 vin_n.n137 vss 0.163639f
C8105 vin_n.t3 vss 0.128597f
C8106 vin_n.t1 vss 0.128597f
C8107 vin_n.n138 vss 0.126618f
C8108 vin_n.n139 vss 0.163639f
C8109 vin_n.t160 vss 0.128597f
C8110 vin_n.t159 vss 0.128597f
C8111 vin_n.n140 vss 0.126618f
C8112 vin_n.n141 vss 0.163639f
C8113 vin_n.t151 vss 0.128597f
C8114 vin_n.t148 vss 0.128597f
C8115 vin_n.n142 vss 0.126618f
C8116 vin_n.n143 vss 0.163639f
C8117 vin_n.t174 vss 0.128597f
C8118 vin_n.t171 vss 0.128597f
C8119 vin_n.n144 vss 0.126618f
C8120 vin_n.n145 vss 0.163639f
C8121 vin_n.t169 vss 0.128597f
C8122 vin_n.t167 vss 0.128597f
C8123 vin_n.n146 vss 0.126618f
C8124 vin_n.n147 vss 0.163639f
C8125 vin_n.t87 vss 0.128597f
C8126 vin_n.t86 vss 0.128597f
C8127 vin_n.n148 vss 0.126618f
C8128 vin_n.n149 vss 0.163639f
C8129 vin_n.t40 vss 0.128597f
C8130 vin_n.t38 vss 0.128597f
C8131 vin_n.n150 vss 0.126618f
C8132 vin_n.n151 vss 0.163639f
C8133 vin_n.t32 vss 0.128597f
C8134 vin_n.t31 vss 0.128597f
C8135 vin_n.n152 vss 0.126618f
C8136 vin_n.n153 vss 0.163639f
C8137 vin_n.t27 vss 0.128597f
C8138 vin_n.t26 vss 0.128597f
C8139 vin_n.n154 vss 0.126618f
C8140 vin_n.n155 vss 0.163639f
C8141 vin_n.t19 vss 0.128597f
C8142 vin_n.t17 vss 0.128597f
C8143 vin_n.n156 vss 0.126618f
C8144 vin_n.n157 vss 0.163639f
C8145 vin_n.t157 vss 0.128597f
C8146 vin_n.t155 vss 0.128597f
C8147 vin_n.n158 vss 0.126618f
C8148 vin_n.n159 vss 0.163639f
C8149 vin_n.t120 vss 0.128597f
C8150 vin_n.t118 vss 0.128597f
C8151 vin_n.n160 vss 0.126618f
C8152 vin_n.n161 vss 0.163639f
C8153 vin_n.t112 vss 0.128597f
C8154 vin_n.t110 vss 0.128597f
C8155 vin_n.n162 vss 0.126618f
C8156 vin_n.n163 vss 0.163639f
C8157 vin_n.t108 vss 0.128597f
C8158 vin_n.t106 vss 0.128597f
C8159 vin_n.n164 vss 0.126618f
C8160 vin_n.n165 vss 0.163639f
C8161 vin_n.t103 vss 0.128597f
C8162 vin_n.t102 vss 0.128597f
C8163 vin_n.n166 vss 0.126618f
C8164 vin_n.n167 vss 0.163639f
C8165 vin_n.t99 vss 0.128597f
C8166 vin_n.t98 vss 0.128597f
C8167 vin_n.n168 vss 0.126618f
C8168 vin_n.n169 vss 0.163639f
C8169 vin_n.t182 vss 0.128597f
C8170 vin_n.t181 vss 0.128597f
C8171 vin_n.n170 vss 0.126618f
C8172 vin_n.n171 vss 0.163639f
C8173 vin_n.t180 vss 0.128597f
C8174 vin_n.t179 vss 0.128597f
C8175 vin_n.n172 vss 0.126618f
C8176 vin_n.n173 vss 0.163639f
C8177 vin_n.t177 vss 0.128597f
C8178 vin_n.t176 vss 0.128597f
C8179 vin_n.n174 vss 0.126618f
C8180 vin_n.n175 vss 0.163639f
C8181 vin_n.t173 vss 0.128597f
C8182 vin_n.t170 vss 0.128597f
C8183 vin_n.n176 vss 0.126618f
C8184 vin_n.n177 vss 0.163639f
C8185 vin_n.t186 vss 0.128597f
C8186 vin_n.t185 vss 0.128597f
C8187 vin_n.n178 vss 0.126618f
C8188 vin_n.n179 vss 0.163639f
C8189 vin_n.t128 vss 0.128597f
C8190 vin_n.t127 vss 0.128597f
C8191 vin_n.n180 vss 0.126618f
C8192 vin_n.n181 vss 0.163639f
C8193 vin_n.t61 vss 0.128597f
C8194 vin_n.t59 vss 0.128597f
C8195 vin_n.n182 vss 0.126618f
C8196 vin_n.n183 vss 0.163639f
C8197 vin_n.t55 vss 0.128597f
C8198 vin_n.t53 vss 0.128597f
C8199 vin_n.n184 vss 0.126618f
C8200 vin_n.n185 vss 0.163639f
C8201 vin_n.t51 vss 0.128597f
C8202 vin_n.t49 vss 0.128597f
C8203 vin_n.n186 vss 0.126618f
C8204 vin_n.n187 vss 0.163639f
C8205 vin_n.t45 vss 0.128597f
C8206 vin_n.t44 vss 0.128597f
C8207 vin_n.n188 vss 0.126618f
C8208 vin_n.n189 vss 0.163639f
C8209 vin_n.t191 vss 0.128597f
C8210 vin_n.t189 vss 0.128597f
C8211 vin_n.n190 vss 0.126618f
C8212 vin_n.n191 vss 0.163639f
C8213 vin_n.t119 vss 0.128597f
C8214 vin_n.t117 vss 0.128597f
C8215 vin_n.n192 vss 0.126618f
C8216 vin_n.n193 vss 0.163639f
C8217 vin_n.t136 vss 0.128597f
C8218 vin_n.t135 vss 0.128597f
C8219 vin_n.n194 vss 0.126618f
C8220 vin_n.n195 vss 0.163639f
C8221 vin_n.t133 vss 0.128597f
C8222 vin_n.t130 vss 0.128597f
C8223 vin_n.n196 vss 0.126618f
C8224 vin_n.n197 vss 0.729315f
C8225 vin_n.n198 vss 1.98787f
C8226 vout.n0 vss 11.5269f
C8227 vout.t300 vss 18.4756f
C8228 vout.n1 vss 9.562031f
C8229 vout.n2 vss 0.03822f
C8230 vout.n3 vss 0.041846f
C8231 vout.n4 vss 0.07007f
C8232 vout.t64 vss 0.022897f
C8233 vout.t59 vss 0.022897f
C8234 vout.n5 vss 0.08525f
C8235 vout.t71 vss 0.022897f
C8236 vout.t131 vss 0.022897f
C8237 vout.n6 vss 0.064815f
C8238 vout.n7 vss 0.933316f
C8239 vout.n8 vss 0.079405f
C8240 vout.n9 vss 0.07007f
C8241 vout.t119 vss 0.022897f
C8242 vout.t121 vss 0.022897f
C8243 vout.n10 vss 0.08525f
C8244 vout.t67 vss 0.022897f
C8245 vout.t105 vss 0.022897f
C8246 vout.n11 vss 0.064815f
C8247 vout.n12 vss 0.933316f
C8248 vout.n13 vss 0.079405f
C8249 vout.n14 vss 0.415663f
C8250 vout.t185 vss 0.022897f
C8251 vout.t66 vss 0.022897f
C8252 vout.n15 vss 0.08525f
C8253 vout.t146 vss 0.022897f
C8254 vout.t133 vss 0.022897f
C8255 vout.n16 vss 0.064815f
C8256 vout.n17 vss 0.933316f
C8257 vout.t95 vss 0.110787f
C8258 vout.t73 vss 0.09359f
C8259 vout.n18 vss 0.979206f
C8260 vout.n19 vss 0.275322f
C8261 vout.n20 vss 0.147407f
C8262 vout.n21 vss 0.05529f
C8263 vout.n22 vss 0.054195f
C8264 vout.n23 vss 0.07007f
C8265 vout.n24 vss 0.07007f
C8266 vout.n25 vss 0.031203f
C8267 vout.n26 vss 0.056932f
C8268 vout.n27 vss 0.049816f
C8269 vout.n28 vss 0.07007f
C8270 vout.n29 vss 0.07007f
C8271 vout.n30 vss 0.035583f
C8272 vout.n31 vss 0.056932f
C8273 vout.t77 vss 0.022897f
C8274 vout.t195 vss 0.022897f
C8275 vout.n32 vss 0.08525f
C8276 vout.t181 vss 0.022897f
C8277 vout.t175 vss 0.022897f
C8278 vout.n33 vss 0.064815f
C8279 vout.n34 vss 0.933316f
C8280 vout.n35 vss 0.079981f
C8281 vout.n36 vss 0.04566f
C8282 vout.n37 vss 0.07007f
C8283 vout.n38 vss 0.07007f
C8284 vout.n39 vss 0.07007f
C8285 vout.t68 vss 0.022897f
C8286 vout.t111 vss 0.022897f
C8287 vout.n40 vss 0.08525f
C8288 vout.t203 vss 0.022897f
C8289 vout.t74 vss 0.022897f
C8290 vout.n41 vss 0.064815f
C8291 vout.n42 vss 0.933316f
C8292 vout.n43 vss 0.079985f
C8293 vout.t174 vss 0.022897f
C8294 vout.t143 vss 0.022897f
C8295 vout.n44 vss 0.08525f
C8296 vout.t190 vss 0.022897f
C8297 vout.t113 vss 0.022897f
C8298 vout.n45 vss 0.064815f
C8299 vout.n46 vss 0.933316f
C8300 vout.n47 vss 0.079405f
C8301 vout.n48 vss 0.07007f
C8302 vout.t154 vss 0.022897f
C8303 vout.t151 vss 0.022897f
C8304 vout.n49 vss 0.08525f
C8305 vout.t165 vss 0.022897f
C8306 vout.t202 vss 0.022897f
C8307 vout.n50 vss 0.064815f
C8308 vout.n51 vss 0.933316f
C8309 vout.n52 vss 0.079405f
C8310 vout.n53 vss 0.07007f
C8311 vout.t89 vss 0.022897f
C8312 vout.t80 vss 0.022897f
C8313 vout.n54 vss 0.08525f
C8314 vout.t139 vss 0.022897f
C8315 vout.t136 vss 0.022897f
C8316 vout.n55 vss 0.064815f
C8317 vout.n56 vss 0.933316f
C8318 vout.n57 vss 0.056932f
C8319 vout.n58 vss 0.07007f
C8320 vout.t88 vss 0.022897f
C8321 vout.t193 vss 0.022897f
C8322 vout.n59 vss 0.08525f
C8323 vout.t124 vss 0.022897f
C8324 vout.t115 vss 0.022897f
C8325 vout.n60 vss 0.064815f
C8326 vout.n61 vss 0.933316f
C8327 vout.t84 vss 0.022897f
C8328 vout.t180 vss 0.022897f
C8329 vout.n62 vss 0.080802f
C8330 vout.n63 vss 0.526899f
C8331 vout.t125 vss 0.022897f
C8332 vout.t99 vss 0.022897f
C8333 vout.n64 vss 0.08525f
C8334 vout.t135 vss 0.022897f
C8335 vout.t134 vss 0.022897f
C8336 vout.n65 vss 0.064815f
C8337 vout.n66 vss 0.960223f
C8338 vout.t197 vss 0.022897f
C8339 vout.t144 vss 0.022897f
C8340 vout.n67 vss 0.064815f
C8341 vout.n68 vss 0.407409f
C8342 vout.n69 vss 0.124561f
C8343 vout.n70 vss 0.034779f
C8344 vout.n71 vss 0.039962f
C8345 vout.n72 vss 0.07007f
C8346 vout.t102 vss 0.022897f
C8347 vout.t177 vss 0.022897f
C8348 vout.n73 vss 0.064815f
C8349 vout.n74 vss 0.423242f
C8350 vout.t153 vss 0.022897f
C8351 vout.t169 vss 0.022897f
C8352 vout.n75 vss 0.08525f
C8353 vout.t172 vss 0.022897f
C8354 vout.t142 vss 0.022897f
C8355 vout.n76 vss 0.064815f
C8356 vout.n77 vss 1.00039f
C8357 vout.t63 vss 0.022897f
C8358 vout.t128 vss 0.022897f
C8359 vout.n78 vss 0.077621f
C8360 vout.n79 vss 0.517394f
C8361 vout.n80 vss 0.040657f
C8362 vout.n81 vss 0.099536f
C8363 vout.t104 vss 0.022897f
C8364 vout.t147 vss 0.022897f
C8365 vout.n82 vss 0.08525f
C8366 vout.t70 vss 0.022897f
C8367 vout.t168 vss 0.022897f
C8368 vout.n83 vss 0.064815f
C8369 vout.n84 vss 0.933316f
C8370 vout.n85 vss 0.056932f
C8371 vout.n86 vss 0.07007f
C8372 vout.t85 vss 0.022897f
C8373 vout.t194 vss 0.022897f
C8374 vout.n87 vss 0.08525f
C8375 vout.t166 vss 0.022897f
C8376 vout.t201 vss 0.022897f
C8377 vout.n88 vss 0.064815f
C8378 vout.n89 vss 0.933316f
C8379 vout.n90 vss 0.033119f
C8380 vout.n91 vss 0.07007f
C8381 vout.t140 vss 0.022897f
C8382 vout.t90 vss 0.022897f
C8383 vout.n92 vss 0.08525f
C8384 vout.t150 vss 0.022897f
C8385 vout.t78 vss 0.022897f
C8386 vout.n93 vss 0.064815f
C8387 vout.n94 vss 0.933316f
C8388 vout.n95 vss 0.079405f
C8389 vout.t191 vss 0.022897f
C8390 vout.t200 vss 0.022897f
C8391 vout.n96 vss 0.08525f
C8392 vout.t97 vss 0.022897f
C8393 vout.t87 vss 0.022897f
C8394 vout.n97 vss 0.064815f
C8395 vout.n98 vss 0.933316f
C8396 vout.n99 vss 0.079405f
C8397 vout.n100 vss 0.07007f
C8398 vout.t167 vss 0.022897f
C8399 vout.t123 vss 0.022897f
C8400 vout.n101 vss 0.08525f
C8401 vout.t156 vss 0.022897f
C8402 vout.t162 vss 0.022897f
C8403 vout.n102 vss 0.064815f
C8404 vout.n103 vss 0.933316f
C8405 vout.n104 vss 0.039415f
C8406 vout.n105 vss 0.07007f
C8407 vout.n106 vss 1.85155f
C8408 vout.t75 vss 0.022897f
C8409 vout.t206 vss 0.022897f
C8410 vout.n107 vss 0.08525f
C8411 vout.t61 vss 0.022897f
C8412 vout.t152 vss 0.022897f
C8413 vout.n108 vss 0.064815f
C8414 vout.n109 vss 0.933316f
C8415 vout.n110 vss 0.044068f
C8416 vout.n111 vss 0.07007f
C8417 vout.t155 vss 0.022897f
C8418 vout.t183 vss 0.022897f
C8419 vout.n112 vss 0.08525f
C8420 vout.t198 vss 0.022897f
C8421 vout.t176 vss 0.022897f
C8422 vout.n113 vss 0.064815f
C8423 vout.n114 vss 0.933316f
C8424 vout.n115 vss 0.079405f
C8425 vout.t130 vss 0.022897f
C8426 vout.t145 vss 0.022897f
C8427 vout.n116 vss 0.08525f
C8428 vout.t100 vss 0.022897f
C8429 vout.t108 vss 0.022897f
C8430 vout.n117 vss 0.064815f
C8431 vout.n118 vss 0.933316f
C8432 vout.n119 vss 0.079405f
C8433 vout.n120 vss 0.07007f
C8434 vout.t138 vss 0.022897f
C8435 vout.t186 vss 0.022897f
C8436 vout.n121 vss 0.08525f
C8437 vout.t163 vss 0.022897f
C8438 vout.t65 vss 0.022897f
C8439 vout.n122 vss 0.064815f
C8440 vout.n123 vss 0.933316f
C8441 vout.n124 vss 0.079405f
C8442 vout.n125 vss 0.07007f
C8443 vout.t182 vss 0.022897f
C8444 vout.t110 vss 0.022897f
C8445 vout.n126 vss 0.08525f
C8446 vout.t196 vss 0.022897f
C8447 vout.t158 vss 0.022897f
C8448 vout.n127 vss 0.064815f
C8449 vout.n128 vss 0.933316f
C8450 vout.n129 vss 0.079405f
C8451 vout.n130 vss 0.07007f
C8452 vout.t208 vss 0.022897f
C8453 vout.t62 vss 0.022897f
C8454 vout.n131 vss 0.08525f
C8455 vout.t93 vss 0.022897f
C8456 vout.t161 vss 0.022897f
C8457 vout.n132 vss 0.064815f
C8458 vout.n133 vss 0.933316f
C8459 vout.t170 vss 0.022897f
C8460 vout.t106 vss 0.022897f
C8461 vout.n134 vss 0.08525f
C8462 vout.t82 vss 0.022897f
C8463 vout.t149 vss 0.022897f
C8464 vout.n135 vss 0.064815f
C8465 vout.n136 vss 0.95587f
C8466 vout.n137 vss 0.172125f
C8467 vout.t141 vss 0.022897f
C8468 vout.t76 vss 0.022897f
C8469 vout.n138 vss 0.08525f
C8470 vout.t91 vss 0.022897f
C8471 vout.t117 vss 0.022897f
C8472 vout.n139 vss 0.064815f
C8473 vout.n140 vss 0.933316f
C8474 vout.n141 vss 0.056932f
C8475 vout.n142 vss 0.07007f
C8476 vout.t96 vss 0.022897f
C8477 vout.t126 vss 0.022897f
C8478 vout.n143 vss 0.08525f
C8479 vout.t164 vss 0.022897f
C8480 vout.t207 vss 0.022897f
C8481 vout.n144 vss 0.064815f
C8482 vout.n145 vss 0.933316f
C8483 vout.n146 vss 0.046531f
C8484 vout.n147 vss 0.07007f
C8485 vout.t159 vss 0.022897f
C8486 vout.t173 vss 0.022897f
C8487 vout.n148 vss 0.08525f
C8488 vout.t112 vss 0.022897f
C8489 vout.t72 vss 0.022897f
C8490 vout.n149 vss 0.064815f
C8491 vout.n150 vss 0.933316f
C8492 vout.n151 vss 0.079405f
C8493 vout.t129 vss 0.022897f
C8494 vout.t109 vss 0.022897f
C8495 vout.n152 vss 0.08525f
C8496 vout.t120 vss 0.022897f
C8497 vout.t118 vss 0.022897f
C8498 vout.n153 vss 0.064815f
C8499 vout.n154 vss 0.933316f
C8500 vout.n155 vss 0.079405f
C8501 vout.n156 vss 0.07007f
C8502 vout.t199 vss 0.022897f
C8503 vout.t178 vss 0.022897f
C8504 vout.n157 vss 0.08525f
C8505 vout.t103 vss 0.022897f
C8506 vout.t171 vss 0.022897f
C8507 vout.n158 vss 0.064815f
C8508 vout.n159 vss 0.933316f
C8509 vout.n160 vss 0.079405f
C8510 vout.n161 vss 0.07007f
C8511 vout.n162 vss 0.014507f
C8512 vout.t266 vss 0.015265f
C8513 vout.t298 vss 0.015265f
C8514 vout.n163 vss 0.036928f
C8515 vout.t3 vss 0.015265f
C8516 vout.t299 vss 0.015265f
C8517 vout.n164 vss 0.034443f
C8518 vout.n165 vss 0.638656f
C8519 vout.n166 vss 0.064133f
C8520 vout.n167 vss 0.07007f
C8521 vout.t23 vss 0.015265f
C8522 vout.t292 vss 0.015265f
C8523 vout.n168 vss 0.036928f
C8524 vout.t249 vss 0.015265f
C8525 vout.t253 vss 0.015265f
C8526 vout.n169 vss 0.034443f
C8527 vout.n170 vss 0.638656f
C8528 vout.n171 vss 0.056385f
C8529 vout.n172 vss 0.07007f
C8530 vout.t33 vss 0.015265f
C8531 vout.t216 vss 0.015265f
C8532 vout.n173 vss 0.036928f
C8533 vout.t294 vss 0.015265f
C8534 vout.t220 vss 0.015265f
C8535 vout.n174 vss 0.034443f
C8536 vout.n175 vss 0.638656f
C8537 vout.n176 vss 0.064133f
C8538 vout.n177 vss 0.07007f
C8539 vout.t227 vss 0.015265f
C8540 vout.t55 vss 0.015265f
C8541 vout.n178 vss 0.036928f
C8542 vout.t232 vss 0.015265f
C8543 vout.t262 vss 0.015265f
C8544 vout.n179 vss 0.034443f
C8545 vout.n180 vss 0.638656f
C8546 vout.n181 vss 0.05091f
C8547 vout.n182 vss 0.07007f
C8548 vout.t283 vss 0.061675f
C8549 vout.t246 vss 0.059427f
C8550 vout.n183 vss 0.649984f
C8551 vout.n184 vss 0.118714f
C8552 vout.n185 vss 0.096111f
C8553 vout.t286 vss 0.015265f
C8554 vout.t40 vss 0.015265f
C8555 vout.n186 vss 0.036928f
C8556 vout.t239 vss 0.015265f
C8557 vout.t25 vss 0.015265f
C8558 vout.n187 vss 0.034443f
C8559 vout.n188 vss 0.638656f
C8560 vout.t295 vss 0.015265f
C8561 vout.t13 vss 0.015265f
C8562 vout.n189 vss 0.036928f
C8563 vout.t218 vss 0.015265f
C8564 vout.t247 vss 0.015265f
C8565 vout.n190 vss 0.034443f
C8566 vout.n191 vss 0.638656f
C8567 vout.n192 vss 0.064133f
C8568 vout.n193 vss 0.07007f
C8569 vout.t243 vss 0.015265f
C8570 vout.t34 vss 0.015265f
C8571 vout.n194 vss 0.036928f
C8572 vout.t263 vss 0.015265f
C8573 vout.t296 vss 0.015265f
C8574 vout.n195 vss 0.034443f
C8575 vout.n196 vss 0.638656f
C8576 vout.n197 vss 0.054195f
C8577 vout.n198 vss 0.07007f
C8578 vout.t52 vss 0.015265f
C8579 vout.t223 vss 0.015265f
C8580 vout.n199 vss 0.036928f
C8581 vout.t39 vss 0.015265f
C8582 vout.t48 vss 0.015265f
C8583 vout.n200 vss 0.034443f
C8584 vout.n201 vss 0.638656f
C8585 vout.n202 vss 0.064133f
C8586 vout.n203 vss 0.07007f
C8587 vout.t267 vss 0.015265f
C8588 vout.t252 vss 0.015265f
C8589 vout.n204 vss 0.036928f
C8590 vout.t257 vss 0.015265f
C8591 vout.t224 vss 0.015265f
C8592 vout.n205 vss 0.034443f
C8593 vout.n206 vss 0.638656f
C8594 vout.t24 vss 0.015265f
C8595 vout.t53 vss 0.015265f
C8596 vout.n207 vss 0.036928f
C8597 vout.t290 vss 0.015265f
C8598 vout.t215 vss 0.015265f
C8599 vout.n208 vss 0.034443f
C8600 vout.n209 vss 0.638656f
C8601 vout.n210 vss 0.050995f
C8602 vout.n213 vss 0.07007f
C8603 vout.n214 vss 0.07007f
C8604 vout.t291 vss 0.015265f
C8605 vout.t12 vss 0.015265f
C8606 vout.n215 vss 0.036928f
C8607 vout.t30 vss 0.015265f
C8608 vout.t287 vss 0.015265f
C8609 vout.n216 vss 0.034443f
C8610 vout.n217 vss 0.638656f
C8611 vout.n218 vss 0.064133f
C8612 vout.n219 vss 0.07007f
C8613 vout.t0 vss 0.015265f
C8614 vout.t251 vss 0.015265f
C8615 vout.n220 vss 0.036928f
C8616 vout.t256 vss 0.015265f
C8617 vout.t35 vss 0.015265f
C8618 vout.n221 vss 0.034443f
C8619 vout.n222 vss 0.638656f
C8620 vout.n223 vss 0.05091f
C8621 vout.n224 vss 0.07007f
C8622 vout.t14 vss 0.015265f
C8623 vout.t230 vss 0.015265f
C8624 vout.n225 vss 0.036928f
C8625 vout.t16 vss 0.015265f
C8626 vout.t42 vss 0.015265f
C8627 vout.n226 vss 0.034443f
C8628 vout.n227 vss 0.638656f
C8629 vout.n228 vss 0.064133f
C8630 vout.n229 vss 0.07007f
C8631 vout.t297 vss 0.061675f
C8632 vout.t241 vss 0.059427f
C8633 vout.n230 vss 0.649984f
C8634 vout.n231 vss 0.096111f
C8635 vout.t58 vss 0.015265f
C8636 vout.t288 vss 0.015265f
C8637 vout.n232 vss 0.036928f
C8638 vout.t254 vss 0.015265f
C8639 vout.t9 vss 0.015265f
C8640 vout.n233 vss 0.034443f
C8641 vout.n234 vss 0.638656f
C8642 vout.t4 vss 0.015265f
C8643 vout.t47 vss 0.015265f
C8644 vout.n235 vss 0.036928f
C8645 vout.t233 vss 0.015265f
C8646 vout.t276 vss 0.015265f
C8647 vout.n236 vss 0.034443f
C8648 vout.n237 vss 0.638656f
C8649 vout.n238 vss 0.064133f
C8650 vout.n239 vss 0.07007f
C8651 vout.t37 vss 0.015265f
C8652 vout.t277 vss 0.015265f
C8653 vout.n240 vss 0.036928f
C8654 vout.t212 vss 0.015265f
C8655 vout.t240 vss 0.015265f
C8656 vout.n241 vss 0.034443f
C8657 vout.n242 vss 0.638656f
C8658 vout.n243 vss 0.055837f
C8659 vout.n244 vss 0.07007f
C8660 vout.t29 vss 0.015265f
C8661 vout.t51 vss 0.015265f
C8662 vout.n245 vss 0.036928f
C8663 vout.t222 vss 0.015265f
C8664 vout.t5 vss 0.015265f
C8665 vout.n246 vss 0.034443f
C8666 vout.n247 vss 0.638656f
C8667 vout.n248 vss 0.064133f
C8668 vout.n249 vss 0.07007f
C8669 vout.t49 vss 0.015265f
C8670 vout.t228 vss 0.015265f
C8671 vout.n250 vss 0.036928f
C8672 vout.t10 vss 0.015265f
C8673 vout.t282 vss 0.015265f
C8674 vout.n251 vss 0.034443f
C8675 vout.n252 vss 0.638656f
C8676 vout.n253 vss 0.050363f
C8677 vout.n254 vss 0.07007f
C8678 vout.n255 vss 8.44505f
C8679 vout.t248 vss 0.015265f
C8680 vout.t238 vss 0.015265f
C8681 vout.n256 vss 0.036928f
C8682 vout.t1 vss 0.015265f
C8683 vout.t41 vss 0.015265f
C8684 vout.n257 vss 0.034443f
C8685 vout.n258 vss 0.638656f
C8686 vout.n259 vss 0.064133f
C8687 vout.n260 vss 0.07007f
C8688 vout.t274 vss 0.015265f
C8689 vout.t56 vss 0.015265f
C8690 vout.n261 vss 0.036928f
C8691 vout.t45 vss 0.015265f
C8692 vout.t280 vss 0.015265f
C8693 vout.n262 vss 0.034443f
C8694 vout.n263 vss 0.638656f
C8695 vout.n264 vss 0.044889f
C8696 vout.n265 vss 0.07007f
C8697 vout.t8 vss 0.015265f
C8698 vout.t50 vss 0.015265f
C8699 vout.n266 vss 0.036928f
C8700 vout.t38 vss 0.015265f
C8701 vout.t285 vss 0.015265f
C8702 vout.n267 vss 0.034443f
C8703 vout.n268 vss 0.638656f
C8704 vout.n269 vss 0.056932f
C8705 vout.t226 vss 0.061675f
C8706 vout.t214 vss 0.059427f
C8707 vout.n270 vss 0.653128f
C8708 vout.n271 vss 0.183135f
C8709 vout.t46 vss 0.015265f
C8710 vout.t293 vss 0.015265f
C8711 vout.n272 vss 0.036928f
C8712 vout.t225 vss 0.015265f
C8713 vout.t19 vss 0.015265f
C8714 vout.n273 vss 0.034443f
C8715 vout.n274 vss 0.638656f
C8716 vout.n275 vss 0.093557f
C8717 vout.n276 vss 0.031751f
C8718 vout.n277 vss 0.306161f
C8719 vout.n278 vss 0.07007f
C8720 vout.n279 vss 0.07007f
C8721 vout.n280 vss 0.032846f
C8722 vout.n281 vss 0.064133f
C8723 vout.n282 vss 0.052553f
C8724 vout.t231 vss 0.015265f
C8725 vout.t213 vss 0.015265f
C8726 vout.n283 vss 0.036928f
C8727 vout.t271 vss 0.015265f
C8728 vout.t7 vss 0.015265f
C8729 vout.n284 vss 0.034443f
C8730 vout.n285 vss 0.638656f
C8731 vout.n286 vss 0.064133f
C8732 vout.n287 vss 0.040509f
C8733 vout.n288 vss 0.07007f
C8734 vout.n289 vss 0.07007f
C8735 vout.n290 vss 0.07007f
C8736 vout.n291 vss 0.048173f
C8737 vout.n292 vss 0.064133f
C8738 vout.n293 vss 0.037225f
C8739 vout.n294 vss 0.055837f
C8740 vout.n295 vss 0.07007f
C8741 vout.n296 vss 0.07007f
C8742 vout.n297 vss 0.029561f
C8743 vout.n298 vss 0.054469f
C8744 vout.n299 vss 1.51519f
C8745 vout.t258 vss 0.015265f
C8746 vout.t289 vss 0.015265f
C8747 vout.n300 vss 0.036928f
C8748 vout.t272 vss 0.015265f
C8749 vout.t278 vss 0.015265f
C8750 vout.n301 vss 0.034443f
C8751 vout.n302 vss 0.638656f
C8752 vout.n303 vss 0.064133f
C8753 vout.n304 vss 0.009032f
C8754 vout.n305 vss 0.07007f
C8755 vout.n306 vss 0.07007f
C8756 vout.n307 vss 0.07007f
C8757 vout.n308 vss 0.042699f
C8758 vout.n309 vss 0.064133f
C8759 vout.n310 vss 0.042699f
C8760 vout.n311 vss 0.050363f
C8761 vout.n312 vss 0.07007f
C8762 vout.n313 vss 0.07007f
C8763 vout.n314 vss 0.035035f
C8764 vout.n315 vss 0.056932f
C8765 vout.t260 vss 0.015265f
C8766 vout.t18 vss 0.015265f
C8767 vout.n316 vss 0.036928f
C8768 vout.t275 vss 0.015265f
C8769 vout.t234 vss 0.015265f
C8770 vout.n317 vss 0.034443f
C8771 vout.n318 vss 0.638656f
C8772 vout.n319 vss 0.064133f
C8773 vout.n320 vss 0.029561f
C8774 vout.n321 vss 0.07007f
C8775 vout.n322 vss 0.07007f
C8776 vout.n323 vss 0.07007f
C8777 vout.n324 vss 0.037225f
C8778 vout.n325 vss 0.064133f
C8779 vout.n326 vss 0.048173f
C8780 vout.n327 vss 0.044889f
C8781 vout.n328 vss 0.07007f
C8782 vout.n329 vss 0.07007f
C8783 vout.n330 vss 0.040509f
C8784 vout.n331 vss 0.052553f
C8785 vout.n332 vss 0.152762f
C8786 vout.n333 vss 0.427989f
C8787 vout.n334 vss 0.4295f
C8788 vout.n335 vss 0.111321f
C8789 vout.n336 vss 0.037772f
C8790 vout.n337 vss 0.05529f
C8791 vout.n338 vss 0.07007f
C8792 vout.n339 vss 0.07007f
C8793 vout.n340 vss 0.030108f
C8794 vout.n341 vss 0.056932f
C8795 vout.t31 vss 0.015265f
C8796 vout.t235 vss 0.015265f
C8797 vout.n342 vss 0.036928f
C8798 vout.t244 vss 0.015265f
C8799 vout.t237 vss 0.015265f
C8800 vout.n343 vss 0.034443f
C8801 vout.n344 vss 0.638656f
C8802 vout.n345 vss 0.064133f
C8803 vout.n346 vss 0.034488f
C8804 vout.n347 vss 0.07007f
C8805 vout.n348 vss 0.07007f
C8806 vout.n349 vss 0.07007f
C8807 vout.n350 vss 0.042152f
C8808 vout.n351 vss 0.064133f
C8809 vout.n352 vss 0.043246f
C8810 vout.n353 vss 0.049816f
C8811 vout.n354 vss 0.07007f
C8812 vout.n355 vss 0.07007f
C8813 vout.n356 vss 0.035583f
C8814 vout.n357 vss 0.056932f
C8815 vout.n358 vss 0.029013f
C8816 vout.n359 vss 0.07007f
C8817 vout.n360 vss 0.07007f
C8818 vout.t305 vss 18.4756f
C8819 vout.n362 vss 16.2236f
C8820 vout.t302 vss 18.4756f
C8821 vout.n363 vss 16.4113f
C8822 vout.t22 vss 0.015265f
C8823 vout.t2 vss 0.015265f
C8824 vout.n364 vss 0.036928f
C8825 vout.t273 vss 0.015265f
C8826 vout.t229 vss 0.015265f
C8827 vout.n365 vss 0.034443f
C8828 vout.n366 vss 0.639416f
C8829 vout.n367 vss 0.07007f
C8830 vout.n368 vss 0.104977f
C8831 vout.n370 vss 0.07007f
C8832 vout.n371 vss 1.7028f
C8833 vout.n373 vss 0.094157f
C8834 vout.n374 vss 0.057564f
C8835 vout.n375 vss 0.041057f
C8836 vout.n376 vss 0.052005f
C8837 vout.n377 vss 0.07007f
C8838 vout.n378 vss 0.07007f
C8839 vout.n379 vss 0.033393f
C8840 vout.n380 vss 0.056932f
C8841 vout.t209 vss 0.015265f
C8842 vout.t284 vss 0.015265f
C8843 vout.n381 vss 0.036928f
C8844 vout.t54 vss 0.015265f
C8845 vout.t269 vss 0.015265f
C8846 vout.n382 vss 0.034443f
C8847 vout.n383 vss 0.638656f
C8848 vout.n384 vss 0.064133f
C8849 vout.n385 vss 0.031203f
C8850 vout.n386 vss 0.07007f
C8851 vout.n387 vss 0.07007f
C8852 vout.n388 vss 0.07007f
C8853 vout.n389 vss 0.038867f
C8854 vout.n390 vss 0.064133f
C8855 vout.n391 vss 0.046531f
C8856 vout.n392 vss 0.046531f
C8857 vout.n393 vss 0.07007f
C8858 vout.n394 vss 0.07007f
C8859 vout.n395 vss 0.038867f
C8860 vout.n396 vss 0.054195f
C8861 vout.n397 vss 0.151264f
C8862 vout.n398 vss 0.420418f
C8863 vout.n399 vss 0.422374f
C8864 vout.n400 vss 0.07007f
C8865 vout.n401 vss 0.030108f
C8866 vout.n402 vss 0.056932f
C8867 vout.t32 vss 0.015265f
C8868 vout.t279 vss 0.015265f
C8869 vout.n403 vss 0.036928f
C8870 vout.t15 vss 0.015265f
C8871 vout.t20 vss 0.015265f
C8872 vout.n404 vss 0.034443f
C8873 vout.n405 vss 0.638656f
C8874 vout.n406 vss 0.064133f
C8875 vout.n407 vss 0.034488f
C8876 vout.n408 vss 0.07007f
C8877 vout.n409 vss 0.07007f
C8878 vout.n410 vss 0.07007f
C8879 vout.n411 vss 0.042152f
C8880 vout.n412 vss 0.064133f
C8881 vout.n413 vss 0.043246f
C8882 vout.n414 vss 0.049816f
C8883 vout.n415 vss 0.07007f
C8884 vout.n416 vss 0.07007f
C8885 vout.n417 vss 0.035583f
C8886 vout.n418 vss 0.056932f
C8887 vout.t250 vss 0.015265f
C8888 vout.t57 vss 0.015265f
C8889 vout.n419 vss 0.036928f
C8890 vout.t255 vss 0.015265f
C8891 vout.t242 vss 0.015265f
C8892 vout.n420 vss 0.034443f
C8893 vout.n421 vss 0.638656f
C8894 vout.n422 vss 0.064133f
C8895 vout.n423 vss 0.029013f
C8896 vout.n424 vss 0.07007f
C8897 vout.n425 vss 0.07007f
C8898 vout.n426 vss 0.07007f
C8899 vout.n427 vss 0.036677f
C8900 vout.n428 vss 0.064133f
C8901 vout.n429 vss 0.048721f
C8902 vout.t27 vss 0.015265f
C8903 vout.t217 vss 0.015265f
C8904 vout.n430 vss 0.036928f
C8905 vout.t11 vss 0.015265f
C8906 vout.t236 vss 0.015265f
C8907 vout.n431 vss 0.034443f
C8908 vout.n432 vss 0.638656f
C8909 vout.n433 vss 0.064133f
C8910 vout.n434 vss 0.044341f
C8911 vout.n435 vss 0.07007f
C8912 vout.n436 vss 0.07007f
C8913 vout.n437 vss 0.07007f
C8914 vout.t210 vss 0.015265f
C8915 vout.t270 vss 0.015265f
C8916 vout.n438 vss 0.036928f
C8917 vout.t265 vss 0.015265f
C8918 vout.t281 vss 0.015265f
C8919 vout.n439 vss 0.034443f
C8920 vout.n440 vss 0.638656f
C8921 vout.n441 vss 0.064133f
C8922 vout.n442 vss 0.07007f
C8923 vout.t28 vss 0.015265f
C8924 vout.t36 vss 0.015265f
C8925 vout.n443 vss 0.036928f
C8926 vout.t221 vss 0.015265f
C8927 vout.t6 vss 0.015265f
C8928 vout.n444 vss 0.034443f
C8929 vout.n445 vss 0.638656f
C8930 vout.n446 vss 0.046531f
C8931 vout.n447 vss 0.40343f
C8932 vout.t259 vss 0.015265f
C8933 vout.t264 vss 0.015265f
C8934 vout.n448 vss 0.036928f
C8935 vout.t219 vss 0.015265f
C8936 vout.t43 vss 0.015265f
C8937 vout.n449 vss 0.034443f
C8938 vout.n450 vss 0.638656f
C8939 vout.n451 vss 0.064133f
C8940 vout.t17 vss 0.015265f
C8941 vout.t26 vss 0.015265f
C8942 vout.n452 vss 0.036928f
C8943 vout.t21 vss 0.015265f
C8944 vout.t211 vss 0.015265f
C8945 vout.n453 vss 0.034443f
C8946 vout.n454 vss 0.638656f
C8947 vout.t245 vss 0.015265f
C8948 vout.t44 vss 0.015265f
C8949 vout.n455 vss 0.036928f
C8950 vout.t268 vss 0.015265f
C8951 vout.t261 vss 0.015265f
C8952 vout.n456 vss 0.034443f
C8953 vout.n457 vss 0.644509f
C8954 vout.n458 vss 0.208187f
C8955 vout.n459 vss 0.117553f
C8956 vout.n460 vss 0.054195f
C8957 vout.n461 vss 0.038867f
C8958 vout.n462 vss 0.07007f
C8959 vout.n463 vss 0.07007f
C8960 vout.n464 vss 0.07007f
C8961 vout.n465 vss 0.046531f
C8962 vout.n466 vss 0.064133f
C8963 vout.n467 vss 0.038867f
C8964 vout.n468 vss 0.054195f
C8965 vout.n469 vss 0.07007f
C8966 vout.n470 vss 0.07007f
C8967 vout.n471 vss 0.031203f
C8968 vout.n472 vss 0.056932f
C8969 vout.n473 vss 0.033393f
C8970 vout.n474 vss 0.07007f
C8971 vout.n475 vss 0.07007f
C8972 vout.n476 vss 0.050089f
C8973 vout.n477 vss 1.86626f
C8974 vout.t304 vss 18.4756f
C8975 vout.n478 vss 16.2062f
C8976 vout.t301 vss 18.4756f
C8977 vout.n479 vss 16.2236f
C8978 vout.t179 vss 0.022897f
C8979 vout.t114 vss 0.022897f
C8980 vout.n480 vss 0.08525f
C8981 vout.t83 vss 0.022897f
C8982 vout.t69 vss 0.022897f
C8983 vout.n481 vss 0.064815f
C8984 vout.n482 vss 0.933316f
C8985 vout.n483 vss 0.079405f
C8986 vout.n484 vss 0.07007f
C8987 vout.t94 vss 0.022897f
C8988 vout.t188 vss 0.022897f
C8989 vout.n485 vss 0.08525f
C8990 vout.t92 vss 0.022897f
C8991 vout.t79 vss 0.022897f
C8992 vout.n486 vss 0.064815f
C8993 vout.n487 vss 0.933316f
C8994 vout.n488 vss 0.079405f
C8995 vout.n489 vss 0.07007f
C8996 vout.t101 vss 0.022897f
C8997 vout.t122 vss 0.022897f
C8998 vout.n490 vss 0.08525f
C8999 vout.t137 vss 0.022897f
C9000 vout.t148 vss 0.022897f
C9001 vout.n491 vss 0.064815f
C9002 vout.n492 vss 0.933316f
C9003 vout.n493 vss 0.056932f
C9004 vout.t204 vss 0.022897f
C9005 vout.t98 vss 0.022897f
C9006 vout.n494 vss 0.08525f
C9007 vout.t187 vss 0.022897f
C9008 vout.t160 vss 0.022897f
C9009 vout.n495 vss 0.064815f
C9010 vout.n496 vss 0.941375f
C9011 vout.n497 vss 0.294885f
C9012 vout.t157 vss 0.022897f
C9013 vout.t81 vss 0.022897f
C9014 vout.n498 vss 0.08525f
C9015 vout.t189 vss 0.022897f
C9016 vout.t184 vss 0.022897f
C9017 vout.n499 vss 0.064815f
C9018 vout.n500 vss 0.933316f
C9019 vout.n501 vss 0.140696f
C9020 vout.n502 vss 0.048721f
C9021 vout.n503 vss 0.454403f
C9022 vout.n504 vss 0.07007f
C9023 vout.n505 vss 0.07007f
C9024 vout.n506 vss 0.032298f
C9025 vout.n507 vss 0.079405f
C9026 vout.n508 vss 0.0531f
C9027 vout.n509 vss 0.056385f
C9028 vout.n510 vss 0.07007f
C9029 vout.n511 vss 0.07007f
C9030 vout.n512 vss 0.029013f
C9031 vout.n513 vss 0.056932f
C9032 vout.n514 vss 0.052005f
C9033 vout.n515 vss 0.07007f
C9034 vout.n516 vss 0.07007f
C9035 vout.n517 vss 0.031477f
C9036 vout.n518 vss 1.85155f
C9037 vout.n519 vss 0.030382f
C9038 vout.n520 vss 0.047626f
C9039 vout.n521 vss 0.07007f
C9040 vout.n522 vss 0.07007f
C9041 vout.n523 vss 0.037772f
C9042 vout.n524 vss 0.056932f
C9043 vout.n525 vss 0.043246f
C9044 vout.n526 vss 0.07007f
C9045 vout.n527 vss 0.07007f
C9046 vout.n528 vss 0.042152f
C9047 vout.n529 vss 0.056932f
C9048 vout.n530 vss 0.038867f
C9049 vout.n531 vss 0.07007f
C9050 vout.n532 vss 0.07007f
C9051 vout.n533 vss 0.07007f
C9052 vout.n534 vss 0.056932f
C9053 vout.n535 vss 0.034488f
C9054 vout.n536 vss 0.079405f
C9055 vout.n537 vss 0.05091f
C9056 vout.n538 vss 0.07007f
C9057 vout.n539 vss 0.07007f
C9058 vout.n540 vss 0.07007f
C9059 vout.n541 vss 0.030108f
C9060 vout.n542 vss 0.079405f
C9061 vout.n543 vss 0.05529f
C9062 vout.n544 vss 0.054195f
C9063 vout.n545 vss 0.398525f
C9064 vout.n546 vss 0.398525f
C9065 vout.t205 vss 0.022897f
C9066 vout.t132 vss 0.022897f
C9067 vout.n547 vss 0.08525f
C9068 vout.t127 vss 0.022897f
C9069 vout.t116 vss 0.022897f
C9070 vout.n548 vss 0.064815f
C9071 vout.n549 vss 0.933316f
C9072 vout.t107 vss 0.022897f
C9073 vout.t60 vss 0.022897f
C9074 vout.n550 vss 0.08525f
C9075 vout.t192 vss 0.022897f
C9076 vout.t86 vss 0.022897f
C9077 vout.n551 vss 0.064815f
C9078 vout.n552 vss 0.95587f
C9079 vout.n553 vss 0.172946f
C9080 vout.n554 vss 0.055016f
C9081 vout.n555 vss 0.054469f
C9082 vout.n556 vss 0.07007f
C9083 vout.n557 vss 0.07007f
C9084 vout.n558 vss 0.03093f
C9085 vout.n559 vss 0.056932f
C9086 vout.n560 vss 0.050089f
C9087 vout.n561 vss 0.07007f
C9088 vout.n562 vss 0.07007f
C9089 vout.n563 vss 0.035309f
C9090 vout.n564 vss 0.056932f
C9091 vout.n565 vss 0.04571f
C9092 vout.n566 vss 0.07007f
C9093 vout.n567 vss 0.07007f
C9094 vout.n568 vss 0.039688f
C9095 vout.n569 vss 0.056932f
C9096 vout.n570 vss 0.041331f
C9097 vout.n571 vss 0.07007f
C9098 vout.n572 vss 0.07007f
C9099 vout.n573 vss 0.07007f
C9100 vout.n574 vss 0.056932f
C9101 vout.n575 vss 0.036951f
C9102 vout.n576 vss 0.079405f
C9103 vout.n577 vss 0.037499f
C9104 vout.n578 vss 0.07007f
C9105 vout.n579 vss 0.07007f
C9106 vout.n580 vss 0.07007f
C9107 vout.n581 vss 0.032572f
C9108 vout.n582 vss 0.079405f
C9109 vout.n583 vss 0.052827f
C9110 vout.n584 vss 0.056658f
C9111 vout.n585 vss 0.07007f
C9112 vout.n586 vss 0.07007f
C9113 vout.n587 vss 0.02874f
C9114 vout.n588 vss 0.056932f
C9115 vout.n589 vss 0.052279f
C9116 vout.n590 vss 0.07007f
C9117 vout.n591 vss 0.07007f
C9118 vout.n592 vss 0.07007f
C9119 vout.n593 vss 0.056932f
C9120 vout.n594 vss 0.0479f
C9121 vout.n595 vss 0.079405f
C9122 vout.n596 vss 0.037499f
C9123 vout.n597 vss 0.07007f
C9124 vout.n598 vss 0.07007f
C9125 vout.n599 vss 0.07007f
C9126 vout.n600 vss 0.04352f
C9127 vout.n601 vss 0.079405f
C9128 vout.n602 vss 0.041878f
C9129 vout.n603 vss 0.067333f
C9130 vout.n604 vss 0.405936f
C9131 vout.n605 vss 0.405936f
C9132 vout.n606 vss 0.07007f
C9133 vout.n607 vss 0.056932f
C9134 vout.n608 vss 0.033393f
C9135 vout.n609 vss 0.079405f
C9136 vout.n610 vss 0.052005f
C9137 vout.n611 vss 0.07007f
C9138 vout.n612 vss 0.07007f
C9139 vout.n613 vss 0.07007f
C9140 vout.n614 vss 0.029013f
C9141 vout.n615 vss 0.079405f
C9142 vout.n616 vss 0.056385f
C9143 vout.n617 vss 0.0531f
C9144 vout.n618 vss 0.07007f
C9145 vout.n619 vss 0.07007f
C9146 vout.n620 vss 0.032298f
C9147 vout.n621 vss 0.056932f
C9148 vout.n622 vss 0.048721f
C9149 vout.n623 vss 0.07007f
C9150 vout.n624 vss 0.07007f
C9151 vout.n625 vss 0.036677f
C9152 vout.n626 vss 0.056932f
C9153 vout.n627 vss 0.044403f
C9154 vout.n628 vss 0.07007f
C9155 vout.n629 vss 0.07007f
C9156 vout.n630 vss 0.07007f
C9157 vout.n631 vss 0.031524f
C9158 vout.n632 vss 1.87429f
C9159 vout.t303 vss 18.4756f
C9160 vout.n633 vss 7.417911f
C9161 vout.n634 vss 9.746651f
C9162 vout.n635 vss 1.55665f
C9163 voe1.n0 vss 2.59057f
C9164 voe1.n1 vss 3.09556f
C9165 voe1.n2 vss 2.59057f
C9166 voe1.n3 vss 2.59057f
C9167 voe1.n4 vss 1.76958f
C9168 voe1.n5 vss 0.115752p
C9169 voe1.n6 vss 18.7701f
C9170 voe1.t111 vss 0.028328f
C9171 voe1.t358 vss 0.246755f
C9172 voe1.t260 vss 0.246755f
C9173 voe1.n7 vss 0.175385f
C9174 voe1.t263 vss 0.246755f
C9175 voe1.t320 vss 0.246755f
C9176 voe1.n8 vss 0.175158f
C9177 voe1.t366 vss 0.246755f
C9178 voe1.t274 vss 0.246755f
C9179 voe1.n9 vss 0.175158f
C9180 voe1.t275 vss 0.246755f
C9181 voe1.t331 vss 0.246755f
C9182 voe1.n10 vss 0.175158f
C9183 voe1.t363 vss 0.246755f
C9184 voe1.t267 vss 0.246755f
C9185 voe1.n11 vss 0.175158f
C9186 voe1.t270 vss 0.246755f
C9187 voe1.t324 vss 0.246755f
C9188 voe1.n12 vss 0.175158f
C9189 voe1.t372 vss 0.246755f
C9190 voe1.t279 vss 0.246755f
C9191 voe1.n13 vss 0.175158f
C9192 voe1.t282 vss 0.246755f
C9193 voe1.t335 vss 0.246755f
C9194 voe1.n14 vss 0.175158f
C9195 voe1.t380 vss 0.246755f
C9196 voe1.t292 vss 0.246755f
C9197 voe1.n15 vss 0.175158f
C9198 voe1.t306 vss 0.246755f
C9199 voe1.t355 vss 0.246755f
C9200 voe1.n16 vss 0.175158f
C9201 voe1.t356 vss 0.246755f
C9202 voe1.t258 vss 0.246755f
C9203 voe1.n17 vss 0.175158f
C9204 voe1.t332 vss 0.246755f
C9205 voe1.t383 vss 0.246755f
C9206 voe1.n18 vss 0.175158f
C9207 voe1.t385 vss 0.246755f
C9208 voe1.t295 vss 0.246755f
C9209 voe1.n19 vss 0.175158f
C9210 voe1.t345 vss 0.246755f
C9211 voe1.t246 vss 0.246755f
C9212 voe1.n20 vss 0.175158f
C9213 voe1.t360 vss 0.246755f
C9214 voe1.t264 vss 0.246755f
C9215 voe1.n21 vss 0.175158f
C9216 voe1.t317 vss 0.246755f
C9217 voe1.t367 vss 0.246755f
C9218 voe1.n22 vss 0.175158f
C9219 voe1.t368 vss 0.246755f
C9220 voe1.t276 vss 0.246755f
C9221 voe1.n23 vss 0.175158f
C9222 voe1.t329 vss 0.246755f
C9223 voe1.t379 vss 0.246755f
C9224 voe1.n24 vss 0.175158f
C9225 voe1.t250 vss 0.246755f
C9226 voe1.t308 vss 0.246755f
C9227 voe1.n25 vss 0.175158f
C9228 voe1.t319 vss 0.246755f
C9229 voe1.t371 vss 0.246755f
C9230 voe1.n26 vss 0.175158f
C9231 voe1.t374 vss 0.246755f
C9232 voe1.t283 vss 0.246755f
C9233 voe1.n27 vss 0.175158f
C9234 voe1.t330 vss 0.246755f
C9235 voe1.t381 vss 0.246755f
C9236 voe1.n28 vss 0.175158f
C9237 voe1.t382 vss 0.246755f
C9238 voe1.t293 vss 0.246755f
C9239 voe1.n29 vss 0.175158f
C9240 voe1.t344 vss 0.246755f
C9241 voe1.t245 vss 0.246755f
C9242 voe1.n30 vss 0.175158f
C9243 voe1.t316 vss 0.246755f
C9244 voe1.t365 vss 0.246755f
C9245 voe1.n31 vss 0.175158f
C9246 voe1.t272 vss 0.246755f
C9247 voe1.t326 vss 0.246755f
C9248 voe1.n32 vss 0.175158f
C9249 voe1.t328 vss 0.246755f
C9250 voe1.t378 vss 0.246755f
C9251 voe1.n33 vss 0.175158f
C9252 voe1.t286 vss 0.246755f
C9253 voe1.t336 vss 0.246755f
C9254 voe1.n34 vss 0.175158f
C9255 voe1.t339 vss 0.246755f
C9256 voe1.t241 vss 0.246755f
C9257 voe1.n35 vss 0.175158f
C9258 voe1.t256 vss 0.246755f
C9259 voe1.t314 vss 0.246755f
C9260 voe1.n36 vss 0.175158f
C9261 voe1.t315 vss 0.246755f
C9262 voe1.t364 vss 0.246755f
C9263 voe1.n37 vss 0.175158f
C9264 voe1.t290 vss 0.246755f
C9265 voe1.t341 vss 0.246755f
C9266 voe1.n38 vss 0.175158f
C9267 voe1.t343 vss 0.246755f
C9268 voe1.t244 vss 0.246755f
C9269 voe1.n39 vss 0.175158f
C9270 voe1.t301 vss 0.246755f
C9271 voe1.t350 vss 0.246755f
C9272 voe1.n40 vss 0.175158f
C9273 voe1.t361 vss 0.246755f
C9274 voe1.t266 vss 0.246755f
C9275 voe1.n41 vss 0.175158f
C9276 voe1.t269 vss 0.246755f
C9277 voe1.t323 vss 0.246755f
C9278 voe1.n42 vss 0.175158f
C9279 voe1.t370 vss 0.246755f
C9280 voe1.t278 vss 0.246755f
C9281 voe1.n43 vss 0.175158f
C9282 voe1.t281 vss 0.246755f
C9283 voe1.t333 vss 0.246755f
C9284 voe1.n44 vss 0.175158f
C9285 voe1.t252 vss 0.246755f
C9286 voe1.t310 vss 0.246755f
C9287 voe1.n45 vss 0.175158f
C9288 voe1.t273 vss 0.246755f
C9289 voe1.t327 vss 0.246755f
C9290 voe1.n46 vss 0.175158f
C9291 voe1.t376 vss 0.246755f
C9292 voe1.t285 vss 0.246755f
C9293 voe1.n47 vss 0.175158f
C9294 voe1.t288 vss 0.246755f
C9295 voe1.t338 vss 0.246755f
C9296 voe1.n48 vss 0.175158f
C9297 voe1.t384 vss 0.246755f
C9298 voe1.t294 vss 0.246755f
C9299 voe1.n49 vss 0.175158f
C9300 voe1.t297 vss 0.246755f
C9301 voe1.t348 vss 0.246755f
C9302 voe1.n50 vss 0.175158f
C9303 voe1.t359 vss 0.246755f
C9304 voe1.t262 vss 0.246755f
C9305 voe1.n51 vss 0.175158f
C9306 voe1.t291 vss 0.246755f
C9307 voe1.t342 vss 0.246755f
C9308 voe1.n52 vss 0.175158f
C9309 voe1.t240 vss 0.246755f
C9310 voe1.t300 vss 0.246755f
C9311 voe1.n53 vss 0.175158f
C9312 voe1.t303 vss 0.246755f
C9313 voe1.t352 vss 0.246755f
C9314 voe1.n54 vss 0.175158f
C9315 voe1.t249 vss 0.246755f
C9316 voe1.t307 vss 0.246755f
C9317 voe1.n55 vss 0.175158f
C9318 voe1.t271 vss 0.246755f
C9319 voe1.t325 vss 0.246755f
C9320 voe1.n56 vss 0.175158f
C9321 voe1.t373 vss 0.246755f
C9322 voe1.t280 vss 0.246755f
C9323 voe1.n57 vss 0.175158f
C9324 voe1.t305 vss 0.246755f
C9325 voe1.t353 vss 0.246755f
C9326 voe1.n58 vss 0.175158f
C9327 voe1.t254 vss 0.246755f
C9328 voe1.t311 vss 0.246755f
C9329 voe1.n59 vss 0.175158f
C9330 voe1.t313 vss 0.246755f
C9331 voe1.t362 vss 0.246755f
C9332 voe1.n60 vss 0.175158f
C9333 voe1.t377 vss 0.246755f
C9334 voe1.t287 vss 0.246755f
C9335 voe1.n61 vss 0.175158f
C9336 voe1.t289 vss 0.246755f
C9337 voe1.t340 vss 0.246755f
C9338 voe1.n62 vss 0.175158f
C9339 voe1.t237 vss 0.246755f
C9340 voe1.t296 vss 0.246755f
C9341 voe1.n63 vss 0.175158f
C9342 voe1.t299 vss 0.246755f
C9343 voe1.t349 vss 0.246755f
C9344 voe1.n64 vss 0.175158f
C9345 voe1.t265 vss 0.246755f
C9346 voe1.t321 vss 0.246755f
C9347 voe1.n65 vss 0.175158f
C9348 voe1.t337 vss 0.246755f
C9349 voe1.t239 vss 0.246755f
C9350 voe1.n66 vss 0.175158f
C9351 voe1.t242 vss 0.246755f
C9352 voe1.t302 vss 0.246755f
C9353 voe1.n67 vss 0.175158f
C9354 voe1.t347 vss 0.246755f
C9355 voe1.t248 vss 0.246755f
C9356 voe1.n68 vss 0.175158f
C9357 voe1.t251 vss 0.246755f
C9358 voe1.t309 vss 0.246755f
C9359 voe1.n69 vss 0.175158f
C9360 voe1.t354 vss 0.246755f
C9361 voe1.t257 vss 0.246755f
C9362 voe1.n70 vss 0.175158f
C9363 voe1.t375 vss 0.246755f
C9364 voe1.t284 vss 0.246755f
C9365 voe1.n71 vss 0.175158f
C9366 voe1.t351 vss 0.246755f
C9367 voe1.t253 vss 0.246755f
C9368 voe1.n72 vss 0.175158f
C9369 voe1.t255 vss 0.246755f
C9370 voe1.t312 vss 0.246755f
C9371 voe1.n73 vss 0.175158f
C9372 voe1.t357 vss 0.246755f
C9373 voe1.t259 vss 0.246755f
C9374 voe1.n74 vss 0.175158f
C9375 voe1.t261 vss 0.246755f
C9376 voe1.t318 vss 0.246755f
C9377 voe1.n75 vss 0.175158f
C9378 voe1.t334 vss 0.246755f
C9379 voe1.t236 vss 0.246755f
C9380 voe1.n76 vss 0.175158f
C9381 voe1.t238 vss 0.246755f
C9382 voe1.t298 vss 0.246755f
C9383 voe1.n77 vss 0.175158f
C9384 voe1.t346 vss 0.246755f
C9385 voe1.t247 vss 0.246755f
C9386 voe1.n78 vss 0.175158f
C9387 voe1.t268 vss 0.246755f
C9388 voe1.t322 vss 0.246755f
C9389 voe1.n79 vss 0.175158f
C9390 voe1.t369 vss 0.246755f
C9391 voe1.t277 vss 0.246755f
C9392 voe1.n80 vss 0.175158f
C9393 voe1.t243 vss 0.246755f
C9394 voe1.t304 vss 0.246755f
C9395 voe1.n81 vss 0.175158f
C9396 voe1.t12 vss 0.027964f
C9397 voe1.t110 vss 0.027964f
C9398 voe1.t77 vss 0.027964f
C9399 voe1.t78 vss 0.027964f
C9400 voe1.t10 vss 0.037069f
C9401 voe1.t199 vss 0.112663f
C9402 voe1.t222 vss 0.029512f
C9403 voe1.t220 vss 0.029512f
C9404 voe1.n82 vss 0.072673f
C9405 voe1.t29 vss 0.125261f
C9406 voe1.t101 vss 0.029512f
C9407 voe1.t57 vss 0.029512f
C9408 voe1.n83 vss 0.087554f
C9409 voe1.t181 vss 0.029512f
C9410 voe1.t50 vss 0.029512f
C9411 voe1.n84 vss 0.063615f
C9412 voe1.t107 vss 0.029512f
C9413 voe1.t206 vss 0.029512f
C9414 voe1.n85 vss 0.063774f
C9415 voe1.t149 vss 0.029512f
C9416 voe1.t71 vss 0.029512f
C9417 voe1.n86 vss 0.063615f
C9418 voe1.t96 vss 0.029512f
C9419 voe1.t228 vss 0.029512f
C9420 voe1.n87 vss 0.063615f
C9421 voe1.t23 vss 0.029512f
C9422 voe1.t145 vss 0.029512f
C9423 voe1.n88 vss 0.063615f
C9424 voe1.t150 vss 0.029512f
C9425 voe1.t180 vss 0.029512f
C9426 voe1.n89 vss 0.063615f
C9427 voe1.t32 vss 0.029512f
C9428 voe1.t215 vss 0.029512f
C9429 voe1.n90 vss 0.063615f
C9430 voe1.t212 vss 0.029512f
C9431 voe1.t232 vss 0.029512f
C9432 voe1.n91 vss 0.063615f
C9433 voe1.t131 vss 0.029512f
C9434 voe1.t17 vss 0.029512f
C9435 voe1.n92 vss 0.063615f
C9436 voe1.t148 vss 0.029512f
C9437 voe1.t136 vss 0.029512f
C9438 voe1.n93 vss 0.063615f
C9439 voe1.t31 vss 0.029512f
C9440 voe1.t115 vss 0.029512f
C9441 voe1.n94 vss 0.063615f
C9442 voe1.t129 vss 0.029512f
C9443 voe1.t205 vss 0.029512f
C9444 voe1.n95 vss 0.063615f
C9445 voe1.t142 vss 0.029512f
C9446 voe1.t120 vss 0.029512f
C9447 voe1.n96 vss 0.063615f
C9448 voe1.t47 vss 0.029512f
C9449 voe1.t155 vss 0.029512f
C9450 voe1.n97 vss 0.063615f
C9451 voe1.t66 vss 0.029512f
C9452 voe1.t203 vss 0.029512f
C9453 voe1.n98 vss 0.063615f
C9454 voe1.t35 vss 0.029512f
C9455 voe1.t75 vss 0.029512f
C9456 voe1.n99 vss 0.063615f
C9457 voe1.t198 vss 0.029512f
C9458 voe1.t69 vss 0.029512f
C9459 voe1.n100 vss 0.063615f
C9460 voe1.t160 vss 0.029512f
C9461 voe1.t37 vss 0.029512f
C9462 voe1.n101 vss 0.063615f
C9463 voe1.t179 vss 0.029512f
C9464 voe1.t19 vss 0.029512f
C9465 voe1.n102 vss 0.063615f
C9466 voe1.t183 vss 0.029512f
C9467 voe1.t1 vss 0.029512f
C9468 voe1.n103 vss 0.063615f
C9469 voe1.t103 vss 0.029512f
C9470 voe1.t90 vss 0.029512f
C9471 voe1.n104 vss 0.063615f
C9472 voe1.t162 vss 0.029512f
C9473 voe1.t146 vss 0.029512f
C9474 voe1.n105 vss 0.063615f
C9475 voe1.t156 vss 0.029512f
C9476 voe1.t15 vss 0.029512f
C9477 voe1.n106 vss 0.063615f
C9478 voe1.t184 vss 0.029512f
C9479 voe1.t196 vss 0.029512f
C9480 voe1.n107 vss 0.063615f
C9481 voe1.t217 vss 0.029512f
C9482 voe1.t76 vss 0.029512f
C9483 voe1.n108 vss 0.063697f
C9484 voe1.t234 vss 0.029512f
C9485 voe1.t64 vss 0.029512f
C9486 voe1.n109 vss 0.063615f
C9487 voe1.t109 vss 0.029512f
C9488 voe1.t46 vss 0.029512f
C9489 voe1.n110 vss 0.063774f
C9490 voe1.t151 vss 0.029512f
C9491 voe1.t130 vss 0.029512f
C9492 voe1.n111 vss 0.063615f
C9493 voe1.t141 vss 0.029512f
C9494 voe1.t97 vss 0.029512f
C9495 voe1.n112 vss 0.063615f
C9496 voe1.t44 vss 0.029512f
C9497 voe1.t26 vss 0.029512f
C9498 voe1.n113 vss 0.063615f
C9499 voe1.t67 vss 0.029512f
C9500 voe1.t197 vss 0.029512f
C9501 voe1.n114 vss 0.063615f
C9502 voe1.t33 vss 0.029512f
C9503 voe1.t13 vss 0.029512f
C9504 voe1.n115 vss 0.063615f
C9505 voe1.t167 vss 0.029512f
C9506 voe1.t91 vss 0.029512f
C9507 voe1.n116 vss 0.063615f
C9508 voe1.t63 vss 0.029512f
C9509 voe1.t211 vss 0.029512f
C9510 voe1.n117 vss 0.063615f
C9511 voe1.t108 vss 0.029512f
C9512 voe1.t42 vss 0.029512f
C9513 voe1.n118 vss 0.063615f
C9514 voe1.t74 vss 0.029512f
C9515 voe1.t86 vss 0.029512f
C9516 voe1.n119 vss 0.063615f
C9517 voe1.t119 vss 0.029512f
C9518 voe1.t128 vss 0.029512f
C9519 voe1.n120 vss 0.063615f
C9520 voe1.t125 vss 0.029512f
C9521 voe1.t52 vss 0.029512f
C9522 voe1.n121 vss 0.063615f
C9523 voe1.t218 vss 0.029512f
C9524 voe1.t164 vss 0.029512f
C9525 voe1.n122 vss 0.063615f
C9526 voe1.t106 vss 0.029512f
C9527 voe1.t79 vss 0.029512f
C9528 voe1.n123 vss 0.063615f
C9529 voe1.t22 vss 0.029512f
C9530 voe1.t40 vss 0.029512f
C9531 voe1.n124 vss 0.063615f
C9532 voe1.t41 vss 0.029512f
C9533 voe1.t27 vss 0.029512f
C9534 voe1.n125 vss 0.063615f
C9535 voe1.t153 vss 0.029512f
C9536 voe1.t161 vss 0.029512f
C9537 voe1.n126 vss 0.063615f
C9538 voe1.t61 vss 0.029512f
C9539 voe1.t4 vss 0.029512f
C9540 voe1.n127 vss 0.063615f
C9541 voe1.t20 vss 0.029512f
C9542 voe1.t2 vss 0.029512f
C9543 voe1.n128 vss 0.063615f
C9544 voe1.t116 vss 0.029512f
C9545 voe1.t133 vss 0.029512f
C9546 voe1.n129 vss 0.063615f
C9547 voe1.t65 vss 0.029512f
C9548 voe1.t186 vss 0.029512f
C9549 voe1.n130 vss 0.063615f
C9550 voe1.t157 vss 0.029512f
C9551 voe1.t14 vss 0.029512f
C9552 voe1.n131 vss 0.063615f
C9553 voe1.t127 vss 0.029512f
C9554 voe1.t182 vss 0.029512f
C9555 voe1.n132 vss 0.063615f
C9556 voe1.t83 vss 0.029512f
C9557 voe1.t9 vss 0.029512f
C9558 voe1.n133 vss 0.063697f
C9559 voe1.t118 vss 0.029512f
C9560 voe1.t98 vss 0.029512f
C9561 voe1.n134 vss 0.063615f
C9562 voe1.t195 vss 0.029512f
C9563 voe1.t193 vss 0.029512f
C9564 voe1.n135 vss 0.063774f
C9565 voe1.t147 vss 0.029512f
C9566 voe1.t72 vss 0.029512f
C9567 voe1.n136 vss 0.063615f
C9568 voe1.t221 vss 0.029512f
C9569 voe1.t16 vss 0.029512f
C9570 voe1.n137 vss 0.063615f
C9571 voe1.t188 vss 0.029512f
C9572 voe1.t93 vss 0.029512f
C9573 voe1.n138 vss 0.063615f
C9574 voe1.t45 vss 0.029512f
C9575 voe1.t5 vss 0.029512f
C9576 voe1.n139 vss 0.063615f
C9577 voe1.t43 vss 0.029512f
C9578 voe1.t140 vss 0.029512f
C9579 voe1.n140 vss 0.063615f
C9580 voe1.t200 vss 0.029512f
C9581 voe1.t143 vss 0.029512f
C9582 voe1.n141 vss 0.063615f
C9583 voe1.t152 vss 0.029512f
C9584 voe1.t8 vss 0.029512f
C9585 voe1.n142 vss 0.063615f
C9586 voe1.t21 vss 0.029512f
C9587 voe1.t168 vss 0.029512f
C9588 voe1.n143 vss 0.063615f
C9589 voe1.t55 vss 0.029512f
C9590 voe1.t169 vss 0.029512f
C9591 voe1.n144 vss 0.063615f
C9592 voe1.t210 vss 0.029512f
C9593 voe1.t202 vss 0.029512f
C9594 voe1.n145 vss 0.063615f
C9595 voe1.t134 vss 0.029512f
C9596 voe1.t30 vss 0.029512f
C9597 voe1.n146 vss 0.063615f
C9598 voe1.t123 vss 0.029512f
C9599 voe1.t25 vss 0.029512f
C9600 voe1.n147 vss 0.063615f
C9601 voe1.t88 vss 0.029512f
C9602 voe1.t53 vss 0.029512f
C9603 voe1.n148 vss 0.063615f
C9604 voe1.t154 vss 0.029512f
C9605 voe1.t190 vss 0.029512f
C9606 voe1.n149 vss 0.063615f
C9607 voe1.t87 vss 0.029512f
C9608 voe1.t81 vss 0.029512f
C9609 voe1.n150 vss 0.063615f
C9610 voe1.t18 vss 0.029512f
C9611 voe1.t231 vss 0.029512f
C9612 voe1.n151 vss 0.063615f
C9613 voe1.t235 vss 0.029512f
C9614 voe1.t178 vss 0.029512f
C9615 voe1.n152 vss 0.063615f
C9616 voe1.t39 vss 0.029512f
C9617 voe1.t176 vss 0.029512f
C9618 voe1.n153 vss 0.063615f
C9619 voe1.t117 vss 0.029512f
C9620 voe1.t80 vss 0.029512f
C9621 voe1.n154 vss 0.063615f
C9622 voe1.t36 vss 0.029512f
C9623 voe1.t233 vss 0.029512f
C9624 voe1.n155 vss 0.063615f
C9625 voe1.t166 vss 0.029512f
C9626 voe1.t219 vss 0.029512f
C9627 voe1.n156 vss 0.063615f
C9628 voe1.t174 vss 0.029512f
C9629 voe1.t158 vss 0.029512f
C9630 voe1.n157 vss 0.063615f
C9631 voe1.t121 vss 0.029512f
C9632 voe1.t177 vss 0.029512f
C9633 voe1.n158 vss 0.063697f
C9634 voe1.t194 vss 0.029512f
C9635 voe1.t185 vss 0.029512f
C9636 voe1.n159 vss 0.063774f
C9637 voe1.t60 vss 0.029512f
C9638 voe1.t171 vss 0.029512f
C9639 voe1.n160 vss 0.063615f
C9640 voe1.t89 vss 0.029512f
C9641 voe1.t7 vss 0.029512f
C9642 voe1.n161 vss 0.063615f
C9643 voe1.t213 vss 0.029512f
C9644 voe1.t92 vss 0.029512f
C9645 voe1.n162 vss 0.063615f
C9646 voe1.t38 vss 0.029512f
C9647 voe1.t3 vss 0.029512f
C9648 voe1.n163 vss 0.063615f
C9649 voe1.t95 vss 0.029512f
C9650 voe1.t102 vss 0.029512f
C9651 voe1.n164 vss 0.063615f
C9652 voe1.t99 vss 0.029512f
C9653 voe1.t24 vss 0.029512f
C9654 voe1.n165 vss 0.063615f
C9655 voe1.t172 vss 0.029512f
C9656 voe1.t34 vss 0.029512f
C9657 voe1.n166 vss 0.063615f
C9658 voe1.t207 vss 0.029512f
C9659 voe1.t173 vss 0.029512f
C9660 voe1.n167 vss 0.063615f
C9661 voe1.t126 vss 0.029512f
C9662 voe1.t0 vss 0.029512f
C9663 voe1.n168 vss 0.063615f
C9664 voe1.t73 vss 0.029512f
C9665 voe1.t175 vss 0.029512f
C9666 voe1.n169 vss 0.063615f
C9667 voe1.t170 vss 0.029512f
C9668 voe1.t6 vss 0.029512f
C9669 voe1.n170 vss 0.063615f
C9670 voe1.t122 vss 0.029512f
C9671 voe1.t209 vss 0.029512f
C9672 voe1.n171 vss 0.063615f
C9673 voe1.t54 vss 0.029512f
C9674 voe1.t124 vss 0.029512f
C9675 voe1.n172 vss 0.063615f
C9676 voe1.t216 vss 0.029512f
C9677 voe1.t208 vss 0.029512f
C9678 voe1.n173 vss 0.063615f
C9679 voe1.t163 vss 0.029512f
C9680 voe1.t56 vss 0.029512f
C9681 voe1.n174 vss 0.063615f
C9682 voe1.t191 vss 0.029512f
C9683 voe1.t204 vss 0.029512f
C9684 voe1.n175 vss 0.063615f
C9685 voe1.t82 vss 0.029512f
C9686 voe1.t112 vss 0.029512f
C9687 voe1.n176 vss 0.063615f
C9688 voe1.t187 vss 0.029512f
C9689 voe1.t68 vss 0.029512f
C9690 voe1.n177 vss 0.063615f
C9691 voe1.t201 vss 0.029512f
C9692 voe1.t49 vss 0.029512f
C9693 voe1.n178 vss 0.063615f
C9694 voe1.t192 vss 0.029512f
C9695 voe1.t189 vss 0.029512f
C9696 voe1.n179 vss 0.063615f
C9697 voe1.t144 vss 0.029512f
C9698 voe1.t70 vss 0.029512f
C9699 voe1.n180 vss 0.063615f
C9700 voe1.t165 vss 0.029512f
C9701 voe1.t214 vss 0.029512f
C9702 voe1.n181 vss 0.063615f
C9703 voe1.t227 vss 0.029512f
C9704 voe1.t159 vss 0.029512f
C9705 voe1.n182 vss 0.063615f
C9706 voe1.t94 vss 0.029512f
C9707 voe1.t62 vss 0.029512f
C9708 voe1.n183 vss 0.063697f
C9709 voe1.t58 vss 0.029512f
C9710 voe1.t225 vss 0.029512f
C9711 voe1.n184 vss 0.081241f
C9712 voe1.t132 vss 0.029512f
C9713 voe1.t28 vss 0.029512f
C9714 voe1.n185 vss 0.081241f
C9715 voe1.t11 vss 0.029512f
C9716 voe1.t230 vss 0.029512f
C9717 voe1.n186 vss 0.081241f
C9718 voe1.t223 vss 0.029512f
C9719 voe1.t226 vss 0.029512f
C9720 voe1.n187 vss 0.081241f
C9721 voe1.t113 vss 0.029512f
C9722 voe1.t84 vss 0.029512f
C9723 voe1.n188 vss 0.081241f
C9724 voe1.t51 vss 0.029512f
C9725 voe1.t135 vss 0.029512f
C9726 voe1.n189 vss 0.081241f
C9727 voe1.t138 vss 0.029512f
C9728 voe1.t48 vss 0.029512f
C9729 voe1.n190 vss 0.072673f
C9730 voe1.t100 vss 0.029512f
C9731 voe1.t59 vss 0.029512f
C9732 voe1.n191 vss 0.073638f
C9733 voe1.t224 vss 0.029512f
C9734 voe1.t105 vss 0.029512f
C9735 voe1.n192 vss 0.072673f
C9736 voe1.t229 vss 0.029512f
C9737 voe1.t137 vss 0.029512f
C9738 voe1.n193 vss 0.072673f
C9739 voe1.t114 vss 0.029512f
C9740 voe1.t104 vss 0.029512f
C9741 voe1.n194 vss 0.072673f
C9742 voe1.t85 vss 0.029512f
C9743 voe1.t139 vss 0.029512f
C9744 voe1.n195 vss 0.072673f
.ends


magic
tech sky130A
magscale 1 2
timestamp 1702073221
<< error_p >>
rect -29 5475 29 5481
rect -29 5441 -17 5475
rect -29 5435 29 5441
rect -29 2719 29 2725
rect -29 2685 -17 2719
rect -29 2679 29 2685
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -2793 29 -2787
rect -29 -2827 -17 -2793
rect -29 -2833 29 -2827
<< pwell >>
rect -226 -5613 226 5613
<< nmos >>
rect -30 2803 30 5403
rect -30 47 30 2647
rect -30 -2709 30 -109
rect -30 -5465 30 -2865
<< ndiff >>
rect -88 5391 -30 5403
rect -88 2815 -76 5391
rect -42 2815 -30 5391
rect -88 2803 -30 2815
rect 30 5391 88 5403
rect 30 2815 42 5391
rect 76 2815 88 5391
rect 30 2803 88 2815
rect -88 2635 -30 2647
rect -88 59 -76 2635
rect -42 59 -30 2635
rect -88 47 -30 59
rect 30 2635 88 2647
rect 30 59 42 2635
rect 76 59 88 2635
rect 30 47 88 59
rect -88 -121 -30 -109
rect -88 -2697 -76 -121
rect -42 -2697 -30 -121
rect -88 -2709 -30 -2697
rect 30 -121 88 -109
rect 30 -2697 42 -121
rect 76 -2697 88 -121
rect 30 -2709 88 -2697
rect -88 -2877 -30 -2865
rect -88 -5453 -76 -2877
rect -42 -5453 -30 -2877
rect -88 -5465 -30 -5453
rect 30 -2877 88 -2865
rect 30 -5453 42 -2877
rect 76 -5453 88 -2877
rect 30 -5465 88 -5453
<< ndiffc >>
rect -76 2815 -42 5391
rect 42 2815 76 5391
rect -76 59 -42 2635
rect 42 59 76 2635
rect -76 -2697 -42 -121
rect 42 -2697 76 -121
rect -76 -5453 -42 -2877
rect 42 -5453 76 -2877
<< psubdiff >>
rect -190 5543 190 5577
rect -190 -5543 -156 5543
rect 156 -5543 190 5543
rect -190 -5577 -94 -5543
rect 94 -5577 190 -5543
<< psubdiffcont >>
rect -94 -5577 94 -5543
<< poly >>
rect -33 5475 33 5491
rect -33 5441 -17 5475
rect 17 5441 33 5475
rect -33 5425 33 5441
rect -30 5403 30 5425
rect -30 2777 30 2803
rect -33 2719 33 2735
rect -33 2685 -17 2719
rect 17 2685 33 2719
rect -33 2669 33 2685
rect -30 2647 30 2669
rect -30 21 30 47
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -30 -109 30 -87
rect -30 -2735 30 -2709
rect -33 -2793 33 -2777
rect -33 -2827 -17 -2793
rect 17 -2827 33 -2793
rect -33 -2843 33 -2827
rect -30 -2865 30 -2843
rect -30 -5491 30 -5465
<< polycont >>
rect -17 5441 17 5475
rect -17 2685 17 2719
rect -17 -71 17 -37
rect -17 -2827 17 -2793
<< locali >>
rect -33 5441 -17 5475
rect 17 5441 33 5475
rect -76 5391 -42 5407
rect -76 2799 -42 2815
rect 42 5391 76 5407
rect 42 2799 76 2815
rect -33 2685 -17 2719
rect 17 2685 33 2719
rect -76 2635 -42 2651
rect -76 43 -42 59
rect 42 2635 76 2651
rect 42 43 76 59
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -76 -121 -42 -105
rect -76 -2713 -42 -2697
rect 42 -121 76 -105
rect 42 -2713 76 -2697
rect -33 -2827 -17 -2793
rect 17 -2827 33 -2793
rect -76 -2877 -42 -2861
rect -76 -5469 -42 -5453
rect 42 -2877 76 -2861
rect 42 -5469 76 -5453
rect -110 -5577 -94 -5543
rect 94 -5577 110 -5543
<< viali >>
rect -17 5441 17 5475
rect -76 2815 -42 5391
rect 42 3201 76 5005
rect -17 2685 17 2719
rect -76 59 -42 2635
rect 42 445 76 2249
rect -17 -71 17 -37
rect -76 -2697 -42 -121
rect 42 -2311 76 -507
rect -17 -2827 17 -2793
rect -76 -5453 -42 -2877
rect 42 -5067 76 -3263
<< metal1 >>
rect -29 5475 29 5481
rect -29 5441 -17 5475
rect 17 5441 29 5475
rect -29 5435 29 5441
rect -82 5391 -36 5403
rect -82 2815 -76 5391
rect -42 2815 -36 5391
rect 36 5005 82 5017
rect 36 3201 42 5005
rect 76 3201 82 5005
rect 36 3189 82 3201
rect -82 2803 -36 2815
rect -29 2719 29 2725
rect -29 2685 -17 2719
rect 17 2685 29 2719
rect -29 2679 29 2685
rect -82 2635 -36 2647
rect -82 59 -76 2635
rect -42 59 -36 2635
rect 36 2249 82 2261
rect 36 445 42 2249
rect 76 445 82 2249
rect 36 433 82 445
rect -82 47 -36 59
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -82 -121 -36 -109
rect -82 -2697 -76 -121
rect -42 -2697 -36 -121
rect 36 -507 82 -495
rect 36 -2311 42 -507
rect 76 -2311 82 -507
rect 36 -2323 82 -2311
rect -82 -2709 -36 -2697
rect -29 -2793 29 -2787
rect -29 -2827 -17 -2793
rect 17 -2827 29 -2793
rect -29 -2833 29 -2827
rect -82 -2877 -36 -2865
rect -82 -5453 -76 -2877
rect -42 -5453 -36 -2877
rect 36 -3263 82 -3251
rect 36 -5067 42 -3263
rect 76 -5067 82 -3263
rect 36 -5079 82 -5067
rect -82 -5465 -36 -5453
<< properties >>
string FIXED_BBOX -173 -5560 173 5560
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 13 l 0.3 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 70 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

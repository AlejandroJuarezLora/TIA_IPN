magic
tech sky130A
magscale 1 2
timestamp 1701914711
<< pwell >>
rect -451 -1017 451 1017
<< psubdiff >>
rect -415 947 -319 981
rect 319 947 415 981
rect -415 -947 -381 947
rect 381 -947 415 947
rect -415 -981 415 -947
<< psubdiffcont >>
rect -319 947 319 981
<< xpolycontact >>
rect -285 419 285 851
rect -285 -851 285 -419
<< ppolyres >>
rect -285 -419 285 419
<< locali >>
rect -335 947 -319 981
rect 319 947 335 981
<< viali >>
rect -269 436 269 833
rect -269 -833 269 -436
<< metal1 >>
rect -281 833 281 839
rect -281 436 -269 833
rect 269 436 281 833
rect -281 430 281 436
rect -281 -436 281 -430
rect -281 -833 -269 -436
rect 269 -833 281 -436
rect -281 -839 281 -833
<< properties >>
string FIXED_BBOX -398 -964 398 964
string gencell sky130_fd_pr__res_high_po_2p85
string library sky130
string parameters w 2.850 l 4.35 m 1 nx 1 wmin 2.850 lmin 0.50 rho 319.8 val 624.831 dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 0 grc 0 gtc 1 gbc 0 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 0 wmax 2.850 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1701460012
<< nwell >>
rect 4660 3188 10894 3189
rect 4660 1868 24723 3188
rect 4660 -4741 10894 1569
rect 15633 1031 16473 1868
rect 19756 1031 20596 1868
rect 23879 1031 24719 1868
rect 4739 -6610 5032 -6466
rect 4660 -6791 10894 -6610
<< pwell >>
rect 4021 -10028 25495 -6990
<< pmos >>
rect 4856 590 4916 1190
rect 4974 590 5034 1190
rect 5092 590 5152 1190
rect 5210 590 5270 1190
rect 5328 590 5388 1190
rect 5446 590 5506 1190
rect 5564 590 5624 1190
rect 5682 590 5742 1190
rect 5800 590 5860 1190
rect 5918 590 5978 1190
rect 6036 590 6096 1190
rect 6154 590 6214 1190
rect 6272 590 6332 1190
rect 6390 590 6450 1190
rect 6508 590 6568 1190
rect 6626 590 6686 1190
rect 6744 590 6804 1190
rect 6862 590 6922 1190
rect 6980 590 7040 1190
rect 7098 590 7158 1190
rect 7216 590 7276 1190
rect 7334 590 7394 1190
rect 7452 590 7512 1190
rect 7570 590 7630 1190
rect 7688 590 7748 1190
rect 7806 590 7866 1190
rect 7924 590 7984 1190
rect 8042 590 8102 1190
rect 8160 590 8220 1190
rect 8278 590 8338 1190
rect 8396 590 8456 1190
rect 8514 590 8574 1190
rect 8632 590 8692 1190
rect 8750 590 8810 1190
rect 8868 590 8928 1190
rect 8986 590 9046 1190
rect 9104 590 9164 1190
rect 9222 590 9282 1190
rect 9340 590 9400 1190
rect 9458 590 9518 1190
rect 9576 590 9636 1190
rect 9694 590 9754 1190
rect 9812 590 9872 1190
rect 9930 590 9990 1190
rect 10048 590 10108 1190
rect 10166 590 10226 1190
rect 10284 590 10344 1190
rect 10402 590 10462 1190
rect 10520 590 10580 1190
rect 10638 590 10698 1190
rect 4856 -246 4916 354
rect 4974 -246 5034 354
rect 5092 -246 5152 354
rect 5210 -246 5270 354
rect 5328 -246 5388 354
rect 5446 -246 5506 354
rect 5564 -246 5624 354
rect 5682 -246 5742 354
rect 5800 -246 5860 354
rect 5918 -246 5978 354
rect 6036 -246 6096 354
rect 6154 -246 6214 354
rect 6272 -246 6332 354
rect 6390 -246 6450 354
rect 6508 -246 6568 354
rect 6626 -246 6686 354
rect 6744 -246 6804 354
rect 6862 -246 6922 354
rect 6980 -246 7040 354
rect 7098 -246 7158 354
rect 7216 -246 7276 354
rect 7334 -246 7394 354
rect 7452 -246 7512 354
rect 7570 -246 7630 354
rect 7688 -246 7748 354
rect 7806 -246 7866 354
rect 7924 -246 7984 354
rect 8042 -246 8102 354
rect 8160 -246 8220 354
rect 8278 -246 8338 354
rect 8396 -246 8456 354
rect 8514 -246 8574 354
rect 8632 -246 8692 354
rect 8750 -246 8810 354
rect 8868 -246 8928 354
rect 8986 -246 9046 354
rect 9104 -246 9164 354
rect 9222 -246 9282 354
rect 9340 -246 9400 354
rect 9458 -246 9518 354
rect 9576 -246 9636 354
rect 9694 -246 9754 354
rect 9812 -246 9872 354
rect 9930 -246 9990 354
rect 10048 -246 10108 354
rect 10166 -246 10226 354
rect 10284 -246 10344 354
rect 10402 -246 10462 354
rect 10520 -246 10580 354
rect 10638 -246 10698 354
rect 4856 -1460 4916 -860
rect 4974 -1460 5034 -860
rect 5092 -1460 5152 -860
rect 5210 -1460 5270 -860
rect 5328 -1460 5388 -860
rect 5446 -1460 5506 -860
rect 5564 -1460 5624 -860
rect 5682 -1460 5742 -860
rect 5800 -1460 5860 -860
rect 5918 -1460 5978 -860
rect 6036 -1460 6096 -860
rect 6154 -1460 6214 -860
rect 6272 -1460 6332 -860
rect 6390 -1460 6450 -860
rect 6508 -1460 6568 -860
rect 6626 -1460 6686 -860
rect 6744 -1460 6804 -860
rect 6862 -1460 6922 -860
rect 6980 -1460 7040 -860
rect 7098 -1460 7158 -860
rect 7216 -1460 7276 -860
rect 7334 -1460 7394 -860
rect 7452 -1460 7512 -860
rect 7570 -1460 7630 -860
rect 7688 -1460 7748 -860
rect 7806 -1460 7866 -860
rect 7924 -1460 7984 -860
rect 8042 -1460 8102 -860
rect 8160 -1460 8220 -860
rect 8278 -1460 8338 -860
rect 8396 -1460 8456 -860
rect 8514 -1460 8574 -860
rect 8632 -1460 8692 -860
rect 8750 -1460 8810 -860
rect 8868 -1460 8928 -860
rect 8986 -1460 9046 -860
rect 9104 -1460 9164 -860
rect 9222 -1460 9282 -860
rect 9340 -1460 9400 -860
rect 9458 -1460 9518 -860
rect 9576 -1460 9636 -860
rect 9694 -1460 9754 -860
rect 9812 -1460 9872 -860
rect 9930 -1460 9990 -860
rect 10048 -1460 10108 -860
rect 10166 -1460 10226 -860
rect 10284 -1460 10344 -860
rect 10402 -1460 10462 -860
rect 10520 -1460 10580 -860
rect 10638 -1460 10698 -860
rect 4856 -2296 4916 -1696
rect 4974 -2296 5034 -1696
rect 5092 -2296 5152 -1696
rect 5210 -2296 5270 -1696
rect 5328 -2296 5388 -1696
rect 5446 -2296 5506 -1696
rect 5564 -2296 5624 -1696
rect 5682 -2296 5742 -1696
rect 5800 -2296 5860 -1696
rect 5918 -2296 5978 -1696
rect 6036 -2296 6096 -1696
rect 6154 -2296 6214 -1696
rect 6272 -2296 6332 -1696
rect 6390 -2296 6450 -1696
rect 6508 -2296 6568 -1696
rect 6626 -2296 6686 -1696
rect 6744 -2296 6804 -1696
rect 6862 -2296 6922 -1696
rect 6980 -2296 7040 -1696
rect 7098 -2296 7158 -1696
rect 7216 -2296 7276 -1696
rect 7334 -2296 7394 -1696
rect 7452 -2296 7512 -1696
rect 7570 -2296 7630 -1696
rect 7688 -2296 7748 -1696
rect 7806 -2296 7866 -1696
rect 7924 -2296 7984 -1696
rect 8042 -2296 8102 -1696
rect 8160 -2296 8220 -1696
rect 8278 -2296 8338 -1696
rect 8396 -2296 8456 -1696
rect 8514 -2296 8574 -1696
rect 8632 -2296 8692 -1696
rect 8750 -2296 8810 -1696
rect 8868 -2296 8928 -1696
rect 8986 -2296 9046 -1696
rect 9104 -2296 9164 -1696
rect 9222 -2296 9282 -1696
rect 9340 -2296 9400 -1696
rect 9458 -2296 9518 -1696
rect 9576 -2296 9636 -1696
rect 9694 -2296 9754 -1696
rect 9812 -2296 9872 -1696
rect 9930 -2296 9990 -1696
rect 10048 -2296 10108 -1696
rect 10166 -2296 10226 -1696
rect 10284 -2296 10344 -1696
rect 10402 -2296 10462 -1696
rect 10520 -2296 10580 -1696
rect 10638 -2296 10698 -1696
rect 4856 -3510 4916 -2910
rect 4974 -3510 5034 -2910
rect 5092 -3510 5152 -2910
rect 5210 -3510 5270 -2910
rect 5328 -3510 5388 -2910
rect 5446 -3510 5506 -2910
rect 5564 -3510 5624 -2910
rect 5682 -3510 5742 -2910
rect 5800 -3510 5860 -2910
rect 5918 -3510 5978 -2910
rect 6036 -3510 6096 -2910
rect 6154 -3510 6214 -2910
rect 6272 -3510 6332 -2910
rect 6390 -3510 6450 -2910
rect 6508 -3510 6568 -2910
rect 6626 -3510 6686 -2910
rect 6744 -3510 6804 -2910
rect 6862 -3510 6922 -2910
rect 6980 -3510 7040 -2910
rect 7098 -3510 7158 -2910
rect 7216 -3510 7276 -2910
rect 7334 -3510 7394 -2910
rect 7452 -3510 7512 -2910
rect 7570 -3510 7630 -2910
rect 7688 -3510 7748 -2910
rect 7806 -3510 7866 -2910
rect 7924 -3510 7984 -2910
rect 8042 -3510 8102 -2910
rect 8160 -3510 8220 -2910
rect 8278 -3510 8338 -2910
rect 8396 -3510 8456 -2910
rect 8514 -3510 8574 -2910
rect 8632 -3510 8692 -2910
rect 8750 -3510 8810 -2910
rect 8868 -3510 8928 -2910
rect 8986 -3510 9046 -2910
rect 9104 -3510 9164 -2910
rect 9222 -3510 9282 -2910
rect 9340 -3510 9400 -2910
rect 9458 -3510 9518 -2910
rect 9576 -3510 9636 -2910
rect 9694 -3510 9754 -2910
rect 9812 -3510 9872 -2910
rect 9930 -3510 9990 -2910
rect 10048 -3510 10108 -2910
rect 10166 -3510 10226 -2910
rect 10284 -3510 10344 -2910
rect 10402 -3510 10462 -2910
rect 10520 -3510 10580 -2910
rect 10638 -3510 10698 -2910
rect 4856 -4346 4916 -3746
rect 4974 -4346 5034 -3746
rect 5092 -4346 5152 -3746
rect 5210 -4346 5270 -3746
rect 5328 -4346 5388 -3746
rect 5446 -4346 5506 -3746
rect 5564 -4346 5624 -3746
rect 5682 -4346 5742 -3746
rect 5800 -4346 5860 -3746
rect 5918 -4346 5978 -3746
rect 6036 -4346 6096 -3746
rect 6154 -4346 6214 -3746
rect 6272 -4346 6332 -3746
rect 6390 -4346 6450 -3746
rect 6508 -4346 6568 -3746
rect 6626 -4346 6686 -3746
rect 6744 -4346 6804 -3746
rect 6862 -4346 6922 -3746
rect 6980 -4346 7040 -3746
rect 7098 -4346 7158 -3746
rect 7216 -4346 7276 -3746
rect 7334 -4346 7394 -3746
rect 7452 -4346 7512 -3746
rect 7570 -4346 7630 -3746
rect 7688 -4346 7748 -3746
rect 7806 -4346 7866 -3746
rect 7924 -4346 7984 -3746
rect 8042 -4346 8102 -3746
rect 8160 -4346 8220 -3746
rect 8278 -4346 8338 -3746
rect 8396 -4346 8456 -3746
rect 8514 -4346 8574 -3746
rect 8632 -4346 8692 -3746
rect 8750 -4346 8810 -3746
rect 8868 -4346 8928 -3746
rect 8986 -4346 9046 -3746
rect 9104 -4346 9164 -3746
rect 9222 -4346 9282 -3746
rect 9340 -4346 9400 -3746
rect 9458 -4346 9518 -3746
rect 9576 -4346 9636 -3746
rect 9694 -4346 9754 -3746
rect 9812 -4346 9872 -3746
rect 9930 -4346 9990 -3746
rect 10048 -4346 10108 -3746
rect 10166 -4346 10226 -3746
rect 10284 -4346 10344 -3746
rect 10402 -4346 10462 -3746
rect 10520 -4346 10580 -3746
rect 10638 -4346 10698 -3746
<< ndiff >>
rect 10839 -7377 10897 -7365
rect 10839 -7503 10851 -7377
rect 10885 -7503 10897 -7377
rect 10839 -7515 10897 -7503
rect 10927 -7377 10985 -7365
rect 10927 -7503 10939 -7377
rect 10973 -7503 10985 -7377
rect 10927 -7515 10985 -7503
rect 11155 -7377 11213 -7365
rect 11155 -7503 11167 -7377
rect 11201 -7503 11213 -7377
rect 11155 -7515 11213 -7503
rect 11243 -7377 11301 -7365
rect 11243 -7503 11255 -7377
rect 11289 -7503 11301 -7377
rect 11243 -7515 11301 -7503
rect 11471 -7377 11529 -7365
rect 11471 -7503 11483 -7377
rect 11517 -7503 11529 -7377
rect 11471 -7515 11529 -7503
rect 11559 -7377 11617 -7365
rect 11559 -7503 11571 -7377
rect 11605 -7503 11617 -7377
rect 11559 -7515 11617 -7503
rect 11787 -7377 11845 -7365
rect 11787 -7503 11799 -7377
rect 11833 -7503 11845 -7377
rect 11787 -7515 11845 -7503
rect 11875 -7377 11933 -7365
rect 11875 -7503 11887 -7377
rect 11921 -7503 11933 -7377
rect 11875 -7515 11933 -7503
rect 12103 -7377 12161 -7365
rect 12103 -7503 12115 -7377
rect 12149 -7503 12161 -7377
rect 12103 -7515 12161 -7503
rect 12191 -7377 12249 -7365
rect 12191 -7503 12203 -7377
rect 12237 -7503 12249 -7377
rect 12191 -7515 12249 -7503
<< pdiff >>
rect 4798 1178 4856 1190
rect 4798 602 4810 1178
rect 4844 602 4856 1178
rect 4798 590 4856 602
rect 4916 1178 4974 1190
rect 4916 602 4928 1178
rect 4962 602 4974 1178
rect 4916 590 4974 602
rect 5034 1178 5092 1190
rect 5034 602 5046 1178
rect 5080 602 5092 1178
rect 5034 590 5092 602
rect 5152 1178 5210 1190
rect 5152 602 5164 1178
rect 5198 602 5210 1178
rect 5152 590 5210 602
rect 5270 1178 5328 1190
rect 5270 602 5282 1178
rect 5316 602 5328 1178
rect 5270 590 5328 602
rect 5388 1178 5446 1190
rect 5388 602 5400 1178
rect 5434 602 5446 1178
rect 5388 590 5446 602
rect 5506 1178 5564 1190
rect 5506 602 5518 1178
rect 5552 602 5564 1178
rect 5506 590 5564 602
rect 5624 1178 5682 1190
rect 5624 602 5636 1178
rect 5670 602 5682 1178
rect 5624 590 5682 602
rect 5742 1178 5800 1190
rect 5742 602 5754 1178
rect 5788 602 5800 1178
rect 5742 590 5800 602
rect 5860 1178 5918 1190
rect 5860 602 5872 1178
rect 5906 602 5918 1178
rect 5860 590 5918 602
rect 5978 1178 6036 1190
rect 5978 602 5990 1178
rect 6024 602 6036 1178
rect 5978 590 6036 602
rect 6096 1178 6154 1190
rect 6096 602 6108 1178
rect 6142 602 6154 1178
rect 6096 590 6154 602
rect 6214 1178 6272 1190
rect 6214 602 6226 1178
rect 6260 602 6272 1178
rect 6214 590 6272 602
rect 6332 1178 6390 1190
rect 6332 602 6344 1178
rect 6378 602 6390 1178
rect 6332 590 6390 602
rect 6450 1178 6508 1190
rect 6450 602 6462 1178
rect 6496 602 6508 1178
rect 6450 590 6508 602
rect 6568 1178 6626 1190
rect 6568 602 6580 1178
rect 6614 602 6626 1178
rect 6568 590 6626 602
rect 6686 1178 6744 1190
rect 6686 602 6698 1178
rect 6732 602 6744 1178
rect 6686 590 6744 602
rect 6804 1178 6862 1190
rect 6804 602 6816 1178
rect 6850 602 6862 1178
rect 6804 590 6862 602
rect 6922 1178 6980 1190
rect 6922 602 6934 1178
rect 6968 602 6980 1178
rect 6922 590 6980 602
rect 7040 1178 7098 1190
rect 7040 602 7052 1178
rect 7086 602 7098 1178
rect 7040 590 7098 602
rect 7158 1178 7216 1190
rect 7158 602 7170 1178
rect 7204 602 7216 1178
rect 7158 590 7216 602
rect 7276 1178 7334 1190
rect 7276 602 7288 1178
rect 7322 602 7334 1178
rect 7276 590 7334 602
rect 7394 1178 7452 1190
rect 7394 602 7406 1178
rect 7440 602 7452 1178
rect 7394 590 7452 602
rect 7512 1178 7570 1190
rect 7512 602 7524 1178
rect 7558 602 7570 1178
rect 7512 590 7570 602
rect 7630 1178 7688 1190
rect 7630 602 7642 1178
rect 7676 602 7688 1178
rect 7630 590 7688 602
rect 7748 1178 7806 1190
rect 7748 602 7760 1178
rect 7794 602 7806 1178
rect 7748 590 7806 602
rect 7866 1178 7924 1190
rect 7866 602 7878 1178
rect 7912 602 7924 1178
rect 7866 590 7924 602
rect 7984 1178 8042 1190
rect 7984 602 7996 1178
rect 8030 602 8042 1178
rect 7984 590 8042 602
rect 8102 1178 8160 1190
rect 8102 602 8114 1178
rect 8148 602 8160 1178
rect 8102 590 8160 602
rect 8220 1178 8278 1190
rect 8220 602 8232 1178
rect 8266 602 8278 1178
rect 8220 590 8278 602
rect 8338 1178 8396 1190
rect 8338 602 8350 1178
rect 8384 602 8396 1178
rect 8338 590 8396 602
rect 8456 1178 8514 1190
rect 8456 602 8468 1178
rect 8502 602 8514 1178
rect 8456 590 8514 602
rect 8574 1178 8632 1190
rect 8574 602 8586 1178
rect 8620 602 8632 1178
rect 8574 590 8632 602
rect 8692 1178 8750 1190
rect 8692 602 8704 1178
rect 8738 602 8750 1178
rect 8692 590 8750 602
rect 8810 1178 8868 1190
rect 8810 602 8822 1178
rect 8856 602 8868 1178
rect 8810 590 8868 602
rect 8928 1178 8986 1190
rect 8928 602 8940 1178
rect 8974 602 8986 1178
rect 8928 590 8986 602
rect 9046 1178 9104 1190
rect 9046 602 9058 1178
rect 9092 602 9104 1178
rect 9046 590 9104 602
rect 9164 1178 9222 1190
rect 9164 602 9176 1178
rect 9210 602 9222 1178
rect 9164 590 9222 602
rect 9282 1178 9340 1190
rect 9282 602 9294 1178
rect 9328 602 9340 1178
rect 9282 590 9340 602
rect 9400 1178 9458 1190
rect 9400 602 9412 1178
rect 9446 602 9458 1178
rect 9400 590 9458 602
rect 9518 1178 9576 1190
rect 9518 602 9530 1178
rect 9564 602 9576 1178
rect 9518 590 9576 602
rect 9636 1178 9694 1190
rect 9636 602 9648 1178
rect 9682 602 9694 1178
rect 9636 590 9694 602
rect 9754 1178 9812 1190
rect 9754 602 9766 1178
rect 9800 602 9812 1178
rect 9754 590 9812 602
rect 9872 1178 9930 1190
rect 9872 602 9884 1178
rect 9918 602 9930 1178
rect 9872 590 9930 602
rect 9990 1178 10048 1190
rect 9990 602 10002 1178
rect 10036 602 10048 1178
rect 9990 590 10048 602
rect 10108 1178 10166 1190
rect 10108 602 10120 1178
rect 10154 602 10166 1178
rect 10108 590 10166 602
rect 10226 1178 10284 1190
rect 10226 602 10238 1178
rect 10272 602 10284 1178
rect 10226 590 10284 602
rect 10344 1178 10402 1190
rect 10344 602 10356 1178
rect 10390 602 10402 1178
rect 10344 590 10402 602
rect 10462 1178 10520 1190
rect 10462 602 10474 1178
rect 10508 602 10520 1178
rect 10462 590 10520 602
rect 10580 1178 10638 1190
rect 10580 602 10592 1178
rect 10626 602 10638 1178
rect 10580 590 10638 602
rect 10698 1178 10756 1190
rect 10698 602 10710 1178
rect 10744 602 10756 1178
rect 10698 590 10756 602
rect 4798 342 4856 354
rect 4798 -234 4810 342
rect 4844 -234 4856 342
rect 4798 -246 4856 -234
rect 4916 342 4974 354
rect 4916 -234 4928 342
rect 4962 -234 4974 342
rect 4916 -246 4974 -234
rect 5034 342 5092 354
rect 5034 -234 5046 342
rect 5080 -234 5092 342
rect 5034 -246 5092 -234
rect 5152 342 5210 354
rect 5152 -234 5164 342
rect 5198 -234 5210 342
rect 5152 -246 5210 -234
rect 5270 342 5328 354
rect 5270 -234 5282 342
rect 5316 -234 5328 342
rect 5270 -246 5328 -234
rect 5388 342 5446 354
rect 5388 -234 5400 342
rect 5434 -234 5446 342
rect 5388 -246 5446 -234
rect 5506 342 5564 354
rect 5506 -234 5518 342
rect 5552 -234 5564 342
rect 5506 -246 5564 -234
rect 5624 342 5682 354
rect 5624 -234 5636 342
rect 5670 -234 5682 342
rect 5624 -246 5682 -234
rect 5742 342 5800 354
rect 5742 -234 5754 342
rect 5788 -234 5800 342
rect 5742 -246 5800 -234
rect 5860 342 5918 354
rect 5860 -234 5872 342
rect 5906 -234 5918 342
rect 5860 -246 5918 -234
rect 5978 342 6036 354
rect 5978 -234 5990 342
rect 6024 -234 6036 342
rect 5978 -246 6036 -234
rect 6096 342 6154 354
rect 6096 -234 6108 342
rect 6142 -234 6154 342
rect 6096 -246 6154 -234
rect 6214 342 6272 354
rect 6214 -234 6226 342
rect 6260 -234 6272 342
rect 6214 -246 6272 -234
rect 6332 342 6390 354
rect 6332 -234 6344 342
rect 6378 -234 6390 342
rect 6332 -246 6390 -234
rect 6450 342 6508 354
rect 6450 -234 6462 342
rect 6496 -234 6508 342
rect 6450 -246 6508 -234
rect 6568 342 6626 354
rect 6568 -234 6580 342
rect 6614 -234 6626 342
rect 6568 -246 6626 -234
rect 6686 342 6744 354
rect 6686 -234 6698 342
rect 6732 -234 6744 342
rect 6686 -246 6744 -234
rect 6804 342 6862 354
rect 6804 -234 6816 342
rect 6850 -234 6862 342
rect 6804 -246 6862 -234
rect 6922 342 6980 354
rect 6922 -234 6934 342
rect 6968 -234 6980 342
rect 6922 -246 6980 -234
rect 7040 342 7098 354
rect 7040 -234 7052 342
rect 7086 -234 7098 342
rect 7040 -246 7098 -234
rect 7158 342 7216 354
rect 7158 -234 7170 342
rect 7204 -234 7216 342
rect 7158 -246 7216 -234
rect 7276 342 7334 354
rect 7276 -234 7288 342
rect 7322 -234 7334 342
rect 7276 -246 7334 -234
rect 7394 342 7452 354
rect 7394 -234 7406 342
rect 7440 -234 7452 342
rect 7394 -246 7452 -234
rect 7512 342 7570 354
rect 7512 -234 7524 342
rect 7558 -234 7570 342
rect 7512 -246 7570 -234
rect 7630 342 7688 354
rect 7630 -234 7642 342
rect 7676 -234 7688 342
rect 7630 -246 7688 -234
rect 7748 342 7806 354
rect 7748 -234 7760 342
rect 7794 -234 7806 342
rect 7748 -246 7806 -234
rect 7866 342 7924 354
rect 7866 -234 7878 342
rect 7912 -234 7924 342
rect 7866 -246 7924 -234
rect 7984 342 8042 354
rect 7984 -234 7996 342
rect 8030 -234 8042 342
rect 7984 -246 8042 -234
rect 8102 342 8160 354
rect 8102 -234 8114 342
rect 8148 -234 8160 342
rect 8102 -246 8160 -234
rect 8220 342 8278 354
rect 8220 -234 8232 342
rect 8266 -234 8278 342
rect 8220 -246 8278 -234
rect 8338 342 8396 354
rect 8338 -234 8350 342
rect 8384 -234 8396 342
rect 8338 -246 8396 -234
rect 8456 342 8514 354
rect 8456 -234 8468 342
rect 8502 -234 8514 342
rect 8456 -246 8514 -234
rect 8574 342 8632 354
rect 8574 -234 8586 342
rect 8620 -234 8632 342
rect 8574 -246 8632 -234
rect 8692 342 8750 354
rect 8692 -234 8704 342
rect 8738 -234 8750 342
rect 8692 -246 8750 -234
rect 8810 342 8868 354
rect 8810 -234 8822 342
rect 8856 -234 8868 342
rect 8810 -246 8868 -234
rect 8928 342 8986 354
rect 8928 -234 8940 342
rect 8974 -234 8986 342
rect 8928 -246 8986 -234
rect 9046 342 9104 354
rect 9046 -234 9058 342
rect 9092 -234 9104 342
rect 9046 -246 9104 -234
rect 9164 342 9222 354
rect 9164 -234 9176 342
rect 9210 -234 9222 342
rect 9164 -246 9222 -234
rect 9282 342 9340 354
rect 9282 -234 9294 342
rect 9328 -234 9340 342
rect 9282 -246 9340 -234
rect 9400 342 9458 354
rect 9400 -234 9412 342
rect 9446 -234 9458 342
rect 9400 -246 9458 -234
rect 9518 342 9576 354
rect 9518 -234 9530 342
rect 9564 -234 9576 342
rect 9518 -246 9576 -234
rect 9636 342 9694 354
rect 9636 -234 9648 342
rect 9682 -234 9694 342
rect 9636 -246 9694 -234
rect 9754 342 9812 354
rect 9754 -234 9766 342
rect 9800 -234 9812 342
rect 9754 -246 9812 -234
rect 9872 342 9930 354
rect 9872 -234 9884 342
rect 9918 -234 9930 342
rect 9872 -246 9930 -234
rect 9990 342 10048 354
rect 9990 -234 10002 342
rect 10036 -234 10048 342
rect 9990 -246 10048 -234
rect 10108 342 10166 354
rect 10108 -234 10120 342
rect 10154 -234 10166 342
rect 10108 -246 10166 -234
rect 10226 342 10284 354
rect 10226 -234 10238 342
rect 10272 -234 10284 342
rect 10226 -246 10284 -234
rect 10344 342 10402 354
rect 10344 -234 10356 342
rect 10390 -234 10402 342
rect 10344 -246 10402 -234
rect 10462 342 10520 354
rect 10462 -234 10474 342
rect 10508 -234 10520 342
rect 10462 -246 10520 -234
rect 10580 342 10638 354
rect 10580 -234 10592 342
rect 10626 -234 10638 342
rect 10580 -246 10638 -234
rect 10698 342 10756 354
rect 10698 -234 10710 342
rect 10744 -234 10756 342
rect 10698 -246 10756 -234
rect 4798 -872 4856 -860
rect 4798 -1448 4810 -872
rect 4844 -1448 4856 -872
rect 4798 -1460 4856 -1448
rect 4916 -872 4974 -860
rect 4916 -1448 4928 -872
rect 4962 -1448 4974 -872
rect 4916 -1460 4974 -1448
rect 5034 -872 5092 -860
rect 5034 -1448 5046 -872
rect 5080 -1448 5092 -872
rect 5034 -1460 5092 -1448
rect 5152 -872 5210 -860
rect 5152 -1448 5164 -872
rect 5198 -1448 5210 -872
rect 5152 -1460 5210 -1448
rect 5270 -872 5328 -860
rect 5270 -1448 5282 -872
rect 5316 -1448 5328 -872
rect 5270 -1460 5328 -1448
rect 5388 -872 5446 -860
rect 5388 -1448 5400 -872
rect 5434 -1448 5446 -872
rect 5388 -1460 5446 -1448
rect 5506 -872 5564 -860
rect 5506 -1448 5518 -872
rect 5552 -1448 5564 -872
rect 5506 -1460 5564 -1448
rect 5624 -872 5682 -860
rect 5624 -1448 5636 -872
rect 5670 -1448 5682 -872
rect 5624 -1460 5682 -1448
rect 5742 -872 5800 -860
rect 5742 -1448 5754 -872
rect 5788 -1448 5800 -872
rect 5742 -1460 5800 -1448
rect 5860 -872 5918 -860
rect 5860 -1448 5872 -872
rect 5906 -1448 5918 -872
rect 5860 -1460 5918 -1448
rect 5978 -872 6036 -860
rect 5978 -1448 5990 -872
rect 6024 -1448 6036 -872
rect 5978 -1460 6036 -1448
rect 6096 -872 6154 -860
rect 6096 -1448 6108 -872
rect 6142 -1448 6154 -872
rect 6096 -1460 6154 -1448
rect 6214 -872 6272 -860
rect 6214 -1448 6226 -872
rect 6260 -1448 6272 -872
rect 6214 -1460 6272 -1448
rect 6332 -872 6390 -860
rect 6332 -1448 6344 -872
rect 6378 -1448 6390 -872
rect 6332 -1460 6390 -1448
rect 6450 -872 6508 -860
rect 6450 -1448 6462 -872
rect 6496 -1448 6508 -872
rect 6450 -1460 6508 -1448
rect 6568 -872 6626 -860
rect 6568 -1448 6580 -872
rect 6614 -1448 6626 -872
rect 6568 -1460 6626 -1448
rect 6686 -872 6744 -860
rect 6686 -1448 6698 -872
rect 6732 -1448 6744 -872
rect 6686 -1460 6744 -1448
rect 6804 -872 6862 -860
rect 6804 -1448 6816 -872
rect 6850 -1448 6862 -872
rect 6804 -1460 6862 -1448
rect 6922 -872 6980 -860
rect 6922 -1448 6934 -872
rect 6968 -1448 6980 -872
rect 6922 -1460 6980 -1448
rect 7040 -872 7098 -860
rect 7040 -1448 7052 -872
rect 7086 -1448 7098 -872
rect 7040 -1460 7098 -1448
rect 7158 -872 7216 -860
rect 7158 -1448 7170 -872
rect 7204 -1448 7216 -872
rect 7158 -1460 7216 -1448
rect 7276 -872 7334 -860
rect 7276 -1448 7288 -872
rect 7322 -1448 7334 -872
rect 7276 -1460 7334 -1448
rect 7394 -872 7452 -860
rect 7394 -1448 7406 -872
rect 7440 -1448 7452 -872
rect 7394 -1460 7452 -1448
rect 7512 -872 7570 -860
rect 7512 -1448 7524 -872
rect 7558 -1448 7570 -872
rect 7512 -1460 7570 -1448
rect 7630 -872 7688 -860
rect 7630 -1448 7642 -872
rect 7676 -1448 7688 -872
rect 7630 -1460 7688 -1448
rect 7748 -872 7806 -860
rect 7748 -1448 7760 -872
rect 7794 -1448 7806 -872
rect 7748 -1460 7806 -1448
rect 7866 -872 7924 -860
rect 7866 -1448 7878 -872
rect 7912 -1448 7924 -872
rect 7866 -1460 7924 -1448
rect 7984 -872 8042 -860
rect 7984 -1448 7996 -872
rect 8030 -1448 8042 -872
rect 7984 -1460 8042 -1448
rect 8102 -872 8160 -860
rect 8102 -1448 8114 -872
rect 8148 -1448 8160 -872
rect 8102 -1460 8160 -1448
rect 8220 -872 8278 -860
rect 8220 -1448 8232 -872
rect 8266 -1448 8278 -872
rect 8220 -1460 8278 -1448
rect 8338 -872 8396 -860
rect 8338 -1448 8350 -872
rect 8384 -1448 8396 -872
rect 8338 -1460 8396 -1448
rect 8456 -872 8514 -860
rect 8456 -1448 8468 -872
rect 8502 -1448 8514 -872
rect 8456 -1460 8514 -1448
rect 8574 -872 8632 -860
rect 8574 -1448 8586 -872
rect 8620 -1448 8632 -872
rect 8574 -1460 8632 -1448
rect 8692 -872 8750 -860
rect 8692 -1448 8704 -872
rect 8738 -1448 8750 -872
rect 8692 -1460 8750 -1448
rect 8810 -872 8868 -860
rect 8810 -1448 8822 -872
rect 8856 -1448 8868 -872
rect 8810 -1460 8868 -1448
rect 8928 -872 8986 -860
rect 8928 -1448 8940 -872
rect 8974 -1448 8986 -872
rect 8928 -1460 8986 -1448
rect 9046 -872 9104 -860
rect 9046 -1448 9058 -872
rect 9092 -1448 9104 -872
rect 9046 -1460 9104 -1448
rect 9164 -872 9222 -860
rect 9164 -1448 9176 -872
rect 9210 -1448 9222 -872
rect 9164 -1460 9222 -1448
rect 9282 -872 9340 -860
rect 9282 -1448 9294 -872
rect 9328 -1448 9340 -872
rect 9282 -1460 9340 -1448
rect 9400 -872 9458 -860
rect 9400 -1448 9412 -872
rect 9446 -1448 9458 -872
rect 9400 -1460 9458 -1448
rect 9518 -872 9576 -860
rect 9518 -1448 9530 -872
rect 9564 -1448 9576 -872
rect 9518 -1460 9576 -1448
rect 9636 -872 9694 -860
rect 9636 -1448 9648 -872
rect 9682 -1448 9694 -872
rect 9636 -1460 9694 -1448
rect 9754 -872 9812 -860
rect 9754 -1448 9766 -872
rect 9800 -1448 9812 -872
rect 9754 -1460 9812 -1448
rect 9872 -872 9930 -860
rect 9872 -1448 9884 -872
rect 9918 -1448 9930 -872
rect 9872 -1460 9930 -1448
rect 9990 -872 10048 -860
rect 9990 -1448 10002 -872
rect 10036 -1448 10048 -872
rect 9990 -1460 10048 -1448
rect 10108 -872 10166 -860
rect 10108 -1448 10120 -872
rect 10154 -1448 10166 -872
rect 10108 -1460 10166 -1448
rect 10226 -872 10284 -860
rect 10226 -1448 10238 -872
rect 10272 -1448 10284 -872
rect 10226 -1460 10284 -1448
rect 10344 -872 10402 -860
rect 10344 -1448 10356 -872
rect 10390 -1448 10402 -872
rect 10344 -1460 10402 -1448
rect 10462 -872 10520 -860
rect 10462 -1448 10474 -872
rect 10508 -1448 10520 -872
rect 10462 -1460 10520 -1448
rect 10580 -872 10638 -860
rect 10580 -1448 10592 -872
rect 10626 -1448 10638 -872
rect 10580 -1460 10638 -1448
rect 10698 -872 10756 -860
rect 10698 -1448 10710 -872
rect 10744 -1448 10756 -872
rect 10698 -1460 10756 -1448
rect 4798 -1708 4856 -1696
rect 4798 -2284 4810 -1708
rect 4844 -2284 4856 -1708
rect 4798 -2296 4856 -2284
rect 4916 -1708 4974 -1696
rect 4916 -2284 4928 -1708
rect 4962 -2284 4974 -1708
rect 4916 -2296 4974 -2284
rect 5034 -1708 5092 -1696
rect 5034 -2284 5046 -1708
rect 5080 -2284 5092 -1708
rect 5034 -2296 5092 -2284
rect 5152 -1708 5210 -1696
rect 5152 -2284 5164 -1708
rect 5198 -2284 5210 -1708
rect 5152 -2296 5210 -2284
rect 5270 -1708 5328 -1696
rect 5270 -2284 5282 -1708
rect 5316 -2284 5328 -1708
rect 5270 -2296 5328 -2284
rect 5388 -1708 5446 -1696
rect 5388 -2284 5400 -1708
rect 5434 -2284 5446 -1708
rect 5388 -2296 5446 -2284
rect 5506 -1708 5564 -1696
rect 5506 -2284 5518 -1708
rect 5552 -2284 5564 -1708
rect 5506 -2296 5564 -2284
rect 5624 -1708 5682 -1696
rect 5624 -2284 5636 -1708
rect 5670 -2284 5682 -1708
rect 5624 -2296 5682 -2284
rect 5742 -1708 5800 -1696
rect 5742 -2284 5754 -1708
rect 5788 -2284 5800 -1708
rect 5742 -2296 5800 -2284
rect 5860 -1708 5918 -1696
rect 5860 -2284 5872 -1708
rect 5906 -2284 5918 -1708
rect 5860 -2296 5918 -2284
rect 5978 -1708 6036 -1696
rect 5978 -2284 5990 -1708
rect 6024 -2284 6036 -1708
rect 5978 -2296 6036 -2284
rect 6096 -1708 6154 -1696
rect 6096 -2284 6108 -1708
rect 6142 -2284 6154 -1708
rect 6096 -2296 6154 -2284
rect 6214 -1708 6272 -1696
rect 6214 -2284 6226 -1708
rect 6260 -2284 6272 -1708
rect 6214 -2296 6272 -2284
rect 6332 -1708 6390 -1696
rect 6332 -2284 6344 -1708
rect 6378 -2284 6390 -1708
rect 6332 -2296 6390 -2284
rect 6450 -1708 6508 -1696
rect 6450 -2284 6462 -1708
rect 6496 -2284 6508 -1708
rect 6450 -2296 6508 -2284
rect 6568 -1708 6626 -1696
rect 6568 -2284 6580 -1708
rect 6614 -2284 6626 -1708
rect 6568 -2296 6626 -2284
rect 6686 -1708 6744 -1696
rect 6686 -2284 6698 -1708
rect 6732 -2284 6744 -1708
rect 6686 -2296 6744 -2284
rect 6804 -1708 6862 -1696
rect 6804 -2284 6816 -1708
rect 6850 -2284 6862 -1708
rect 6804 -2296 6862 -2284
rect 6922 -1708 6980 -1696
rect 6922 -2284 6934 -1708
rect 6968 -2284 6980 -1708
rect 6922 -2296 6980 -2284
rect 7040 -1708 7098 -1696
rect 7040 -2284 7052 -1708
rect 7086 -2284 7098 -1708
rect 7040 -2296 7098 -2284
rect 7158 -1708 7216 -1696
rect 7158 -2284 7170 -1708
rect 7204 -2284 7216 -1708
rect 7158 -2296 7216 -2284
rect 7276 -1708 7334 -1696
rect 7276 -2284 7288 -1708
rect 7322 -2284 7334 -1708
rect 7276 -2296 7334 -2284
rect 7394 -1708 7452 -1696
rect 7394 -2284 7406 -1708
rect 7440 -2284 7452 -1708
rect 7394 -2296 7452 -2284
rect 7512 -1708 7570 -1696
rect 7512 -2284 7524 -1708
rect 7558 -2284 7570 -1708
rect 7512 -2296 7570 -2284
rect 7630 -1708 7688 -1696
rect 7630 -2284 7642 -1708
rect 7676 -2284 7688 -1708
rect 7630 -2296 7688 -2284
rect 7748 -1708 7806 -1696
rect 7748 -2284 7760 -1708
rect 7794 -2284 7806 -1708
rect 7748 -2296 7806 -2284
rect 7866 -1708 7924 -1696
rect 7866 -2284 7878 -1708
rect 7912 -2284 7924 -1708
rect 7866 -2296 7924 -2284
rect 7984 -1708 8042 -1696
rect 7984 -2284 7996 -1708
rect 8030 -2284 8042 -1708
rect 7984 -2296 8042 -2284
rect 8102 -1708 8160 -1696
rect 8102 -2284 8114 -1708
rect 8148 -2284 8160 -1708
rect 8102 -2296 8160 -2284
rect 8220 -1708 8278 -1696
rect 8220 -2284 8232 -1708
rect 8266 -2284 8278 -1708
rect 8220 -2296 8278 -2284
rect 8338 -1708 8396 -1696
rect 8338 -2284 8350 -1708
rect 8384 -2284 8396 -1708
rect 8338 -2296 8396 -2284
rect 8456 -1708 8514 -1696
rect 8456 -2284 8468 -1708
rect 8502 -2284 8514 -1708
rect 8456 -2296 8514 -2284
rect 8574 -1708 8632 -1696
rect 8574 -2284 8586 -1708
rect 8620 -2284 8632 -1708
rect 8574 -2296 8632 -2284
rect 8692 -1708 8750 -1696
rect 8692 -2284 8704 -1708
rect 8738 -2284 8750 -1708
rect 8692 -2296 8750 -2284
rect 8810 -1708 8868 -1696
rect 8810 -2284 8822 -1708
rect 8856 -2284 8868 -1708
rect 8810 -2296 8868 -2284
rect 8928 -1708 8986 -1696
rect 8928 -2284 8940 -1708
rect 8974 -2284 8986 -1708
rect 8928 -2296 8986 -2284
rect 9046 -1708 9104 -1696
rect 9046 -2284 9058 -1708
rect 9092 -2284 9104 -1708
rect 9046 -2296 9104 -2284
rect 9164 -1708 9222 -1696
rect 9164 -2284 9176 -1708
rect 9210 -2284 9222 -1708
rect 9164 -2296 9222 -2284
rect 9282 -1708 9340 -1696
rect 9282 -2284 9294 -1708
rect 9328 -2284 9340 -1708
rect 9282 -2296 9340 -2284
rect 9400 -1708 9458 -1696
rect 9400 -2284 9412 -1708
rect 9446 -2284 9458 -1708
rect 9400 -2296 9458 -2284
rect 9518 -1708 9576 -1696
rect 9518 -2284 9530 -1708
rect 9564 -2284 9576 -1708
rect 9518 -2296 9576 -2284
rect 9636 -1708 9694 -1696
rect 9636 -2284 9648 -1708
rect 9682 -2284 9694 -1708
rect 9636 -2296 9694 -2284
rect 9754 -1708 9812 -1696
rect 9754 -2284 9766 -1708
rect 9800 -2284 9812 -1708
rect 9754 -2296 9812 -2284
rect 9872 -1708 9930 -1696
rect 9872 -2284 9884 -1708
rect 9918 -2284 9930 -1708
rect 9872 -2296 9930 -2284
rect 9990 -1708 10048 -1696
rect 9990 -2284 10002 -1708
rect 10036 -2284 10048 -1708
rect 9990 -2296 10048 -2284
rect 10108 -1708 10166 -1696
rect 10108 -2284 10120 -1708
rect 10154 -2284 10166 -1708
rect 10108 -2296 10166 -2284
rect 10226 -1708 10284 -1696
rect 10226 -2284 10238 -1708
rect 10272 -2284 10284 -1708
rect 10226 -2296 10284 -2284
rect 10344 -1708 10402 -1696
rect 10344 -2284 10356 -1708
rect 10390 -2284 10402 -1708
rect 10344 -2296 10402 -2284
rect 10462 -1708 10520 -1696
rect 10462 -2284 10474 -1708
rect 10508 -2284 10520 -1708
rect 10462 -2296 10520 -2284
rect 10580 -1708 10638 -1696
rect 10580 -2284 10592 -1708
rect 10626 -2284 10638 -1708
rect 10580 -2296 10638 -2284
rect 10698 -1708 10756 -1696
rect 10698 -2284 10710 -1708
rect 10744 -2284 10756 -1708
rect 10698 -2296 10756 -2284
rect 4798 -2922 4856 -2910
rect 4798 -3498 4810 -2922
rect 4844 -3498 4856 -2922
rect 4798 -3510 4856 -3498
rect 4916 -2922 4974 -2910
rect 4916 -3498 4928 -2922
rect 4962 -3498 4974 -2922
rect 4916 -3510 4974 -3498
rect 5034 -2922 5092 -2910
rect 5034 -3498 5046 -2922
rect 5080 -3498 5092 -2922
rect 5034 -3510 5092 -3498
rect 5152 -2922 5210 -2910
rect 5152 -3498 5164 -2922
rect 5198 -3498 5210 -2922
rect 5152 -3510 5210 -3498
rect 5270 -2922 5328 -2910
rect 5270 -3498 5282 -2922
rect 5316 -3498 5328 -2922
rect 5270 -3510 5328 -3498
rect 5388 -2922 5446 -2910
rect 5388 -3498 5400 -2922
rect 5434 -3498 5446 -2922
rect 5388 -3510 5446 -3498
rect 5506 -2922 5564 -2910
rect 5506 -3498 5518 -2922
rect 5552 -3498 5564 -2922
rect 5506 -3510 5564 -3498
rect 5624 -2922 5682 -2910
rect 5624 -3498 5636 -2922
rect 5670 -3498 5682 -2922
rect 5624 -3510 5682 -3498
rect 5742 -2922 5800 -2910
rect 5742 -3498 5754 -2922
rect 5788 -3498 5800 -2922
rect 5742 -3510 5800 -3498
rect 5860 -2922 5918 -2910
rect 5860 -3498 5872 -2922
rect 5906 -3498 5918 -2922
rect 5860 -3510 5918 -3498
rect 5978 -2922 6036 -2910
rect 5978 -3498 5990 -2922
rect 6024 -3498 6036 -2922
rect 5978 -3510 6036 -3498
rect 6096 -2922 6154 -2910
rect 6096 -3498 6108 -2922
rect 6142 -3498 6154 -2922
rect 6096 -3510 6154 -3498
rect 6214 -2922 6272 -2910
rect 6214 -3498 6226 -2922
rect 6260 -3498 6272 -2922
rect 6214 -3510 6272 -3498
rect 6332 -2922 6390 -2910
rect 6332 -3498 6344 -2922
rect 6378 -3498 6390 -2922
rect 6332 -3510 6390 -3498
rect 6450 -2922 6508 -2910
rect 6450 -3498 6462 -2922
rect 6496 -3498 6508 -2922
rect 6450 -3510 6508 -3498
rect 6568 -2922 6626 -2910
rect 6568 -3498 6580 -2922
rect 6614 -3498 6626 -2922
rect 6568 -3510 6626 -3498
rect 6686 -2922 6744 -2910
rect 6686 -3498 6698 -2922
rect 6732 -3498 6744 -2922
rect 6686 -3510 6744 -3498
rect 6804 -2922 6862 -2910
rect 6804 -3498 6816 -2922
rect 6850 -3498 6862 -2922
rect 6804 -3510 6862 -3498
rect 6922 -2922 6980 -2910
rect 6922 -3498 6934 -2922
rect 6968 -3498 6980 -2922
rect 6922 -3510 6980 -3498
rect 7040 -2922 7098 -2910
rect 7040 -3498 7052 -2922
rect 7086 -3498 7098 -2922
rect 7040 -3510 7098 -3498
rect 7158 -2922 7216 -2910
rect 7158 -3498 7170 -2922
rect 7204 -3498 7216 -2922
rect 7158 -3510 7216 -3498
rect 7276 -2922 7334 -2910
rect 7276 -3498 7288 -2922
rect 7322 -3498 7334 -2922
rect 7276 -3510 7334 -3498
rect 7394 -2922 7452 -2910
rect 7394 -3498 7406 -2922
rect 7440 -3498 7452 -2922
rect 7394 -3510 7452 -3498
rect 7512 -2922 7570 -2910
rect 7512 -3498 7524 -2922
rect 7558 -3498 7570 -2922
rect 7512 -3510 7570 -3498
rect 7630 -2922 7688 -2910
rect 7630 -3498 7642 -2922
rect 7676 -3498 7688 -2922
rect 7630 -3510 7688 -3498
rect 7748 -2922 7806 -2910
rect 7748 -3498 7760 -2922
rect 7794 -3498 7806 -2922
rect 7748 -3510 7806 -3498
rect 7866 -2922 7924 -2910
rect 7866 -3498 7878 -2922
rect 7912 -3498 7924 -2922
rect 7866 -3510 7924 -3498
rect 7984 -2922 8042 -2910
rect 7984 -3498 7996 -2922
rect 8030 -3498 8042 -2922
rect 7984 -3510 8042 -3498
rect 8102 -2922 8160 -2910
rect 8102 -3498 8114 -2922
rect 8148 -3498 8160 -2922
rect 8102 -3510 8160 -3498
rect 8220 -2922 8278 -2910
rect 8220 -3498 8232 -2922
rect 8266 -3498 8278 -2922
rect 8220 -3510 8278 -3498
rect 8338 -2922 8396 -2910
rect 8338 -3498 8350 -2922
rect 8384 -3498 8396 -2922
rect 8338 -3510 8396 -3498
rect 8456 -2922 8514 -2910
rect 8456 -3498 8468 -2922
rect 8502 -3498 8514 -2922
rect 8456 -3510 8514 -3498
rect 8574 -2922 8632 -2910
rect 8574 -3498 8586 -2922
rect 8620 -3498 8632 -2922
rect 8574 -3510 8632 -3498
rect 8692 -2922 8750 -2910
rect 8692 -3498 8704 -2922
rect 8738 -3498 8750 -2922
rect 8692 -3510 8750 -3498
rect 8810 -2922 8868 -2910
rect 8810 -3498 8822 -2922
rect 8856 -3498 8868 -2922
rect 8810 -3510 8868 -3498
rect 8928 -2922 8986 -2910
rect 8928 -3498 8940 -2922
rect 8974 -3498 8986 -2922
rect 8928 -3510 8986 -3498
rect 9046 -2922 9104 -2910
rect 9046 -3498 9058 -2922
rect 9092 -3498 9104 -2922
rect 9046 -3510 9104 -3498
rect 9164 -2922 9222 -2910
rect 9164 -3498 9176 -2922
rect 9210 -3498 9222 -2922
rect 9164 -3510 9222 -3498
rect 9282 -2922 9340 -2910
rect 9282 -3498 9294 -2922
rect 9328 -3498 9340 -2922
rect 9282 -3510 9340 -3498
rect 9400 -2922 9458 -2910
rect 9400 -3498 9412 -2922
rect 9446 -3498 9458 -2922
rect 9400 -3510 9458 -3498
rect 9518 -2922 9576 -2910
rect 9518 -3498 9530 -2922
rect 9564 -3498 9576 -2922
rect 9518 -3510 9576 -3498
rect 9636 -2922 9694 -2910
rect 9636 -3498 9648 -2922
rect 9682 -3498 9694 -2922
rect 9636 -3510 9694 -3498
rect 9754 -2922 9812 -2910
rect 9754 -3498 9766 -2922
rect 9800 -3498 9812 -2922
rect 9754 -3510 9812 -3498
rect 9872 -2922 9930 -2910
rect 9872 -3498 9884 -2922
rect 9918 -3498 9930 -2922
rect 9872 -3510 9930 -3498
rect 9990 -2922 10048 -2910
rect 9990 -3498 10002 -2922
rect 10036 -3498 10048 -2922
rect 9990 -3510 10048 -3498
rect 10108 -2922 10166 -2910
rect 10108 -3498 10120 -2922
rect 10154 -3498 10166 -2922
rect 10108 -3510 10166 -3498
rect 10226 -2922 10284 -2910
rect 10226 -3498 10238 -2922
rect 10272 -3498 10284 -2922
rect 10226 -3510 10284 -3498
rect 10344 -2922 10402 -2910
rect 10344 -3498 10356 -2922
rect 10390 -3498 10402 -2922
rect 10344 -3510 10402 -3498
rect 10462 -2922 10520 -2910
rect 10462 -3498 10474 -2922
rect 10508 -3498 10520 -2922
rect 10462 -3510 10520 -3498
rect 10580 -2922 10638 -2910
rect 10580 -3498 10592 -2922
rect 10626 -3498 10638 -2922
rect 10580 -3510 10638 -3498
rect 10698 -2922 10756 -2910
rect 10698 -3498 10710 -2922
rect 10744 -3498 10756 -2922
rect 10698 -3510 10756 -3498
rect 4798 -3758 4856 -3746
rect 4798 -4334 4810 -3758
rect 4844 -4334 4856 -3758
rect 4798 -4346 4856 -4334
rect 4916 -3758 4974 -3746
rect 4916 -4334 4928 -3758
rect 4962 -4334 4974 -3758
rect 4916 -4346 4974 -4334
rect 5034 -3758 5092 -3746
rect 5034 -4334 5046 -3758
rect 5080 -4334 5092 -3758
rect 5034 -4346 5092 -4334
rect 5152 -3758 5210 -3746
rect 5152 -4334 5164 -3758
rect 5198 -4334 5210 -3758
rect 5152 -4346 5210 -4334
rect 5270 -3758 5328 -3746
rect 5270 -4334 5282 -3758
rect 5316 -4334 5328 -3758
rect 5270 -4346 5328 -4334
rect 5388 -3758 5446 -3746
rect 5388 -4334 5400 -3758
rect 5434 -4334 5446 -3758
rect 5388 -4346 5446 -4334
rect 5506 -3758 5564 -3746
rect 5506 -4334 5518 -3758
rect 5552 -4334 5564 -3758
rect 5506 -4346 5564 -4334
rect 5624 -3758 5682 -3746
rect 5624 -4334 5636 -3758
rect 5670 -4334 5682 -3758
rect 5624 -4346 5682 -4334
rect 5742 -3758 5800 -3746
rect 5742 -4334 5754 -3758
rect 5788 -4334 5800 -3758
rect 5742 -4346 5800 -4334
rect 5860 -3758 5918 -3746
rect 5860 -4334 5872 -3758
rect 5906 -4334 5918 -3758
rect 5860 -4346 5918 -4334
rect 5978 -3758 6036 -3746
rect 5978 -4334 5990 -3758
rect 6024 -4334 6036 -3758
rect 5978 -4346 6036 -4334
rect 6096 -3758 6154 -3746
rect 6096 -4334 6108 -3758
rect 6142 -4334 6154 -3758
rect 6096 -4346 6154 -4334
rect 6214 -3758 6272 -3746
rect 6214 -4334 6226 -3758
rect 6260 -4334 6272 -3758
rect 6214 -4346 6272 -4334
rect 6332 -3758 6390 -3746
rect 6332 -4334 6344 -3758
rect 6378 -4334 6390 -3758
rect 6332 -4346 6390 -4334
rect 6450 -3758 6508 -3746
rect 6450 -4334 6462 -3758
rect 6496 -4334 6508 -3758
rect 6450 -4346 6508 -4334
rect 6568 -3758 6626 -3746
rect 6568 -4334 6580 -3758
rect 6614 -4334 6626 -3758
rect 6568 -4346 6626 -4334
rect 6686 -3758 6744 -3746
rect 6686 -4334 6698 -3758
rect 6732 -4334 6744 -3758
rect 6686 -4346 6744 -4334
rect 6804 -3758 6862 -3746
rect 6804 -4334 6816 -3758
rect 6850 -4334 6862 -3758
rect 6804 -4346 6862 -4334
rect 6922 -3758 6980 -3746
rect 6922 -4334 6934 -3758
rect 6968 -4334 6980 -3758
rect 6922 -4346 6980 -4334
rect 7040 -3758 7098 -3746
rect 7040 -4334 7052 -3758
rect 7086 -4334 7098 -3758
rect 7040 -4346 7098 -4334
rect 7158 -3758 7216 -3746
rect 7158 -4334 7170 -3758
rect 7204 -4334 7216 -3758
rect 7158 -4346 7216 -4334
rect 7276 -3758 7334 -3746
rect 7276 -4334 7288 -3758
rect 7322 -4334 7334 -3758
rect 7276 -4346 7334 -4334
rect 7394 -3758 7452 -3746
rect 7394 -4334 7406 -3758
rect 7440 -4334 7452 -3758
rect 7394 -4346 7452 -4334
rect 7512 -3758 7570 -3746
rect 7512 -4334 7524 -3758
rect 7558 -4334 7570 -3758
rect 7512 -4346 7570 -4334
rect 7630 -3758 7688 -3746
rect 7630 -4334 7642 -3758
rect 7676 -4334 7688 -3758
rect 7630 -4346 7688 -4334
rect 7748 -3758 7806 -3746
rect 7748 -4334 7760 -3758
rect 7794 -4334 7806 -3758
rect 7748 -4346 7806 -4334
rect 7866 -3758 7924 -3746
rect 7866 -4334 7878 -3758
rect 7912 -4334 7924 -3758
rect 7866 -4346 7924 -4334
rect 7984 -3758 8042 -3746
rect 7984 -4334 7996 -3758
rect 8030 -4334 8042 -3758
rect 7984 -4346 8042 -4334
rect 8102 -3758 8160 -3746
rect 8102 -4334 8114 -3758
rect 8148 -4334 8160 -3758
rect 8102 -4346 8160 -4334
rect 8220 -3758 8278 -3746
rect 8220 -4334 8232 -3758
rect 8266 -4334 8278 -3758
rect 8220 -4346 8278 -4334
rect 8338 -3758 8396 -3746
rect 8338 -4334 8350 -3758
rect 8384 -4334 8396 -3758
rect 8338 -4346 8396 -4334
rect 8456 -3758 8514 -3746
rect 8456 -4334 8468 -3758
rect 8502 -4334 8514 -3758
rect 8456 -4346 8514 -4334
rect 8574 -3758 8632 -3746
rect 8574 -4334 8586 -3758
rect 8620 -4334 8632 -3758
rect 8574 -4346 8632 -4334
rect 8692 -3758 8750 -3746
rect 8692 -4334 8704 -3758
rect 8738 -4334 8750 -3758
rect 8692 -4346 8750 -4334
rect 8810 -3758 8868 -3746
rect 8810 -4334 8822 -3758
rect 8856 -4334 8868 -3758
rect 8810 -4346 8868 -4334
rect 8928 -3758 8986 -3746
rect 8928 -4334 8940 -3758
rect 8974 -4334 8986 -3758
rect 8928 -4346 8986 -4334
rect 9046 -3758 9104 -3746
rect 9046 -4334 9058 -3758
rect 9092 -4334 9104 -3758
rect 9046 -4346 9104 -4334
rect 9164 -3758 9222 -3746
rect 9164 -4334 9176 -3758
rect 9210 -4334 9222 -3758
rect 9164 -4346 9222 -4334
rect 9282 -3758 9340 -3746
rect 9282 -4334 9294 -3758
rect 9328 -4334 9340 -3758
rect 9282 -4346 9340 -4334
rect 9400 -3758 9458 -3746
rect 9400 -4334 9412 -3758
rect 9446 -4334 9458 -3758
rect 9400 -4346 9458 -4334
rect 9518 -3758 9576 -3746
rect 9518 -4334 9530 -3758
rect 9564 -4334 9576 -3758
rect 9518 -4346 9576 -4334
rect 9636 -3758 9694 -3746
rect 9636 -4334 9648 -3758
rect 9682 -4334 9694 -3758
rect 9636 -4346 9694 -4334
rect 9754 -3758 9812 -3746
rect 9754 -4334 9766 -3758
rect 9800 -4334 9812 -3758
rect 9754 -4346 9812 -4334
rect 9872 -3758 9930 -3746
rect 9872 -4334 9884 -3758
rect 9918 -4334 9930 -3758
rect 9872 -4346 9930 -4334
rect 9990 -3758 10048 -3746
rect 9990 -4334 10002 -3758
rect 10036 -4334 10048 -3758
rect 9990 -4346 10048 -4334
rect 10108 -3758 10166 -3746
rect 10108 -4334 10120 -3758
rect 10154 -4334 10166 -3758
rect 10108 -4346 10166 -4334
rect 10226 -3758 10284 -3746
rect 10226 -4334 10238 -3758
rect 10272 -4334 10284 -3758
rect 10226 -4346 10284 -4334
rect 10344 -3758 10402 -3746
rect 10344 -4334 10356 -3758
rect 10390 -4334 10402 -3758
rect 10344 -4346 10402 -4334
rect 10462 -3758 10520 -3746
rect 10462 -4334 10474 -3758
rect 10508 -4334 10520 -3758
rect 10462 -4346 10520 -4334
rect 10580 -3758 10638 -3746
rect 10580 -4334 10592 -3758
rect 10626 -4334 10638 -3758
rect 10580 -4346 10638 -4334
rect 10698 -3758 10756 -3746
rect 10698 -4334 10710 -3758
rect 10744 -4334 10756 -3758
rect 10698 -4346 10756 -4334
<< ndiffc >>
rect 6348 -7791 6382 -7215
rect 6466 -7791 6500 -7215
rect 6584 -7791 6618 -7215
rect 6702 -7791 6736 -7215
rect 7874 -7791 7908 -7215
rect 7992 -7791 8026 -7215
rect 8110 -7791 8144 -7215
rect 8228 -7791 8262 -7215
rect 8346 -7791 8380 -7215
rect 8464 -7791 8498 -7215
rect 8582 -7791 8616 -7215
rect 8700 -7791 8734 -7215
rect 8818 -7791 8852 -7215
rect 8936 -7791 8970 -7215
rect 9054 -7791 9088 -7215
rect 9172 -7791 9206 -7215
rect 9290 -7791 9324 -7215
rect 9408 -7791 9442 -7215
rect 9526 -7791 9560 -7215
rect 9644 -7791 9678 -7215
rect 10851 -7503 10885 -7377
rect 10939 -7503 10973 -7377
rect 11167 -7503 11201 -7377
rect 11255 -7503 11289 -7377
rect 11483 -7503 11517 -7377
rect 11571 -7503 11605 -7377
rect 11799 -7503 11833 -7377
rect 11887 -7503 11921 -7377
rect 12115 -7503 12149 -7377
rect 12203 -7503 12237 -7377
rect 6348 -8609 6382 -8033
rect 6466 -8609 6500 -8033
rect 6584 -8609 6618 -8033
rect 6702 -8609 6736 -8033
rect 7874 -8609 7908 -8033
rect 7992 -8609 8026 -8033
rect 8110 -8609 8144 -8033
rect 8228 -8609 8262 -8033
rect 8346 -8609 8380 -8033
rect 8464 -8609 8498 -8033
rect 8582 -8609 8616 -8033
rect 8700 -8609 8734 -8033
rect 8818 -8609 8852 -8033
rect 8936 -8609 8970 -8033
rect 9054 -8609 9088 -8033
rect 9172 -8609 9206 -8033
rect 9290 -8609 9324 -8033
rect 9408 -8609 9442 -8033
rect 9526 -8609 9560 -8033
rect 9644 -8609 9678 -8033
rect 13718 -8091 13752 -7215
rect 13866 -8091 13900 -7215
rect 14014 -8091 14048 -7215
rect 14162 -8091 14196 -7215
rect 14310 -8091 14344 -7215
rect 14458 -8091 14492 -7215
rect 14606 -8091 14640 -7215
rect 14754 -8091 14788 -7215
rect 14902 -8091 14936 -7215
rect 15050 -8091 15084 -7215
rect 15198 -8091 15232 -7215
rect 15346 -8091 15380 -7215
rect 15494 -8091 15528 -7215
rect 15642 -8091 15676 -7215
rect 15790 -8091 15824 -7215
rect 15938 -8091 15972 -7215
rect 16086 -8091 16120 -7215
rect 16234 -8091 16268 -7215
rect 16382 -8091 16416 -7215
rect 16530 -8091 16564 -7215
rect 16678 -8091 16712 -7215
rect 16826 -8091 16860 -7215
rect 16974 -8091 17008 -7215
rect 17122 -8091 17156 -7215
rect 17270 -8091 17304 -7215
rect 17418 -8091 17452 -7215
rect 17566 -8091 17600 -7215
rect 17714 -8091 17748 -7215
rect 17862 -8091 17896 -7215
rect 18010 -8091 18044 -7215
rect 18158 -8091 18192 -7215
rect 18306 -8091 18340 -7215
rect 18454 -8091 18488 -7215
rect 18602 -8091 18636 -7215
rect 18750 -8091 18784 -7215
rect 18898 -8091 18932 -7215
rect 19046 -8091 19080 -7215
rect 19194 -8091 19228 -7215
rect 19342 -8091 19376 -7215
rect 19490 -8091 19524 -7215
rect 19638 -8091 19672 -7215
rect 19786 -8091 19820 -7215
rect 19934 -8091 19968 -7215
rect 20082 -8091 20116 -7215
rect 20230 -8091 20264 -7215
rect 20378 -8091 20412 -7215
rect 20526 -8091 20560 -7215
rect 20674 -8091 20708 -7215
rect 20822 -8091 20856 -7215
rect 20970 -8091 21004 -7215
rect 21118 -8091 21152 -7215
rect 21266 -8091 21300 -7215
rect 21414 -8091 21448 -7215
rect 21562 -8091 21596 -7215
rect 21710 -8091 21744 -7215
rect 21858 -8091 21892 -7215
rect 22006 -8091 22040 -7215
rect 22154 -8091 22188 -7215
rect 22302 -8091 22336 -7215
rect 22450 -8091 22484 -7215
rect 22598 -8091 22632 -7215
rect 22746 -8091 22780 -7215
rect 22894 -8091 22928 -7215
rect 23042 -8091 23076 -7215
rect 21414 -9209 21448 -8333
rect 21562 -9209 21596 -8333
rect 21710 -9209 21744 -8333
rect 21858 -9209 21892 -8333
rect 22006 -9209 22040 -8333
rect 22154 -9209 22188 -8333
rect 22302 -9209 22336 -8333
rect 22450 -9209 22484 -8333
<< pdiffc >>
rect 12972 2098 13006 2674
rect 13090 2098 13124 2674
rect 13208 2098 13242 2674
rect 13326 2098 13360 2674
rect 13444 2098 13478 2674
rect 13562 2098 13596 2674
rect 13680 2098 13714 2674
rect 13798 2098 13832 2674
rect 13916 2098 13950 2674
rect 14034 2098 14068 2674
rect 14152 2098 14186 2674
rect 14270 2098 14304 2674
rect 14388 2098 14422 2674
rect 14506 2098 14540 2674
rect 14624 2098 14658 2674
rect 14742 2098 14776 2674
rect 14860 2098 14894 2674
rect 14978 2098 15012 2674
rect 15096 2098 15130 2674
rect 15214 2098 15248 2674
rect 15332 2098 15366 2674
rect 15450 2098 15484 2674
rect 17095 2098 17129 2674
rect 17213 2098 17247 2674
rect 17331 2098 17365 2674
rect 17449 2098 17483 2674
rect 17567 2098 17601 2674
rect 17685 2098 17719 2674
rect 17803 2098 17837 2674
rect 17921 2098 17955 2674
rect 18039 2098 18073 2674
rect 18157 2098 18191 2674
rect 18275 2098 18309 2674
rect 18393 2098 18427 2674
rect 18511 2098 18545 2674
rect 18629 2098 18663 2674
rect 18747 2098 18781 2674
rect 18865 2098 18899 2674
rect 18983 2098 19017 2674
rect 19101 2098 19135 2674
rect 19219 2098 19253 2674
rect 19337 2098 19371 2674
rect 19455 2098 19489 2674
rect 19573 2098 19607 2674
rect 21218 2098 21252 2674
rect 21336 2098 21370 2674
rect 21454 2098 21488 2674
rect 21572 2098 21606 2674
rect 21690 2098 21724 2674
rect 21808 2098 21842 2674
rect 21926 2098 21960 2674
rect 22044 2098 22078 2674
rect 22162 2098 22196 2674
rect 22280 2098 22314 2674
rect 22398 2098 22432 2674
rect 22516 2098 22550 2674
rect 22634 2098 22668 2674
rect 22752 2098 22786 2674
rect 22870 2098 22904 2674
rect 22988 2098 23022 2674
rect 23106 2098 23140 2674
rect 23224 2098 23258 2674
rect 23342 2098 23376 2674
rect 23460 2098 23494 2674
rect 23578 2098 23612 2674
rect 23696 2098 23730 2674
rect 4810 602 4844 1178
rect 4928 602 4962 1178
rect 5046 602 5080 1178
rect 5164 602 5198 1178
rect 5282 602 5316 1178
rect 5400 602 5434 1178
rect 5518 602 5552 1178
rect 5636 602 5670 1178
rect 5754 602 5788 1178
rect 5872 602 5906 1178
rect 5990 602 6024 1178
rect 6108 602 6142 1178
rect 6226 602 6260 1178
rect 6344 602 6378 1178
rect 6462 602 6496 1178
rect 6580 602 6614 1178
rect 6698 602 6732 1178
rect 6816 602 6850 1178
rect 6934 602 6968 1178
rect 7052 602 7086 1178
rect 7170 602 7204 1178
rect 7288 602 7322 1178
rect 7406 602 7440 1178
rect 7524 602 7558 1178
rect 7642 602 7676 1178
rect 7760 602 7794 1178
rect 7878 602 7912 1178
rect 7996 602 8030 1178
rect 8114 602 8148 1178
rect 8232 602 8266 1178
rect 8350 602 8384 1178
rect 8468 602 8502 1178
rect 8586 602 8620 1178
rect 8704 602 8738 1178
rect 8822 602 8856 1178
rect 8940 602 8974 1178
rect 9058 602 9092 1178
rect 9176 602 9210 1178
rect 9294 602 9328 1178
rect 9412 602 9446 1178
rect 9530 602 9564 1178
rect 9648 602 9682 1178
rect 9766 602 9800 1178
rect 9884 602 9918 1178
rect 10002 602 10036 1178
rect 10120 602 10154 1178
rect 10238 602 10272 1178
rect 10356 602 10390 1178
rect 10474 602 10508 1178
rect 10592 602 10626 1178
rect 10710 602 10744 1178
rect 4810 -234 4844 342
rect 4928 -234 4962 342
rect 5046 -234 5080 342
rect 5164 -234 5198 342
rect 5282 -234 5316 342
rect 5400 -234 5434 342
rect 5518 -234 5552 342
rect 5636 -234 5670 342
rect 5754 -234 5788 342
rect 5872 -234 5906 342
rect 5990 -234 6024 342
rect 6108 -234 6142 342
rect 6226 -234 6260 342
rect 6344 -234 6378 342
rect 6462 -234 6496 342
rect 6580 -234 6614 342
rect 6698 -234 6732 342
rect 6816 -234 6850 342
rect 6934 -234 6968 342
rect 7052 -234 7086 342
rect 7170 -234 7204 342
rect 7288 -234 7322 342
rect 7406 -234 7440 342
rect 7524 -234 7558 342
rect 7642 -234 7676 342
rect 7760 -234 7794 342
rect 7878 -234 7912 342
rect 7996 -234 8030 342
rect 8114 -234 8148 342
rect 8232 -234 8266 342
rect 8350 -234 8384 342
rect 8468 -234 8502 342
rect 8586 -234 8620 342
rect 8704 -234 8738 342
rect 8822 -234 8856 342
rect 8940 -234 8974 342
rect 9058 -234 9092 342
rect 9176 -234 9210 342
rect 9294 -234 9328 342
rect 9412 -234 9446 342
rect 9530 -234 9564 342
rect 9648 -234 9682 342
rect 9766 -234 9800 342
rect 9884 -234 9918 342
rect 10002 -234 10036 342
rect 10120 -234 10154 342
rect 10238 -234 10272 342
rect 10356 -234 10390 342
rect 10474 -234 10508 342
rect 10592 -234 10626 342
rect 10710 -234 10744 342
rect 12972 1262 13006 1838
rect 13090 1262 13124 1838
rect 13208 1262 13242 1838
rect 13326 1262 13360 1838
rect 13444 1262 13478 1838
rect 13562 1262 13596 1838
rect 13680 1262 13714 1838
rect 13798 1262 13832 1838
rect 13916 1262 13950 1838
rect 14034 1262 14068 1838
rect 14152 1262 14186 1838
rect 14270 1262 14304 1838
rect 14388 1262 14422 1838
rect 14506 1262 14540 1838
rect 14624 1262 14658 1838
rect 14742 1262 14776 1838
rect 14860 1262 14894 1838
rect 14978 1262 15012 1838
rect 15096 1262 15130 1838
rect 15214 1262 15248 1838
rect 15332 1262 15366 1838
rect 15450 1262 15484 1838
rect 17095 1262 17129 1838
rect 17213 1262 17247 1838
rect 17331 1262 17365 1838
rect 17449 1262 17483 1838
rect 17567 1262 17601 1838
rect 17685 1262 17719 1838
rect 17803 1262 17837 1838
rect 17921 1262 17955 1838
rect 18039 1262 18073 1838
rect 18157 1262 18191 1838
rect 18275 1262 18309 1838
rect 18393 1262 18427 1838
rect 18511 1262 18545 1838
rect 18629 1262 18663 1838
rect 18747 1262 18781 1838
rect 18865 1262 18899 1838
rect 18983 1262 19017 1838
rect 19101 1262 19135 1838
rect 19219 1262 19253 1838
rect 19337 1262 19371 1838
rect 19455 1262 19489 1838
rect 19573 1262 19607 1838
rect 21218 1262 21252 1838
rect 21336 1262 21370 1838
rect 21454 1262 21488 1838
rect 21572 1262 21606 1838
rect 21690 1262 21724 1838
rect 21808 1262 21842 1838
rect 21926 1262 21960 1838
rect 22044 1262 22078 1838
rect 22162 1262 22196 1838
rect 22280 1262 22314 1838
rect 22398 1262 22432 1838
rect 22516 1262 22550 1838
rect 22634 1262 22668 1838
rect 22752 1262 22786 1838
rect 22870 1262 22904 1838
rect 22988 1262 23022 1838
rect 23106 1262 23140 1838
rect 23224 1262 23258 1838
rect 23342 1262 23376 1838
rect 23460 1262 23494 1838
rect 23578 1262 23612 1838
rect 23696 1262 23730 1838
rect 4810 -1448 4844 -872
rect 4928 -1448 4962 -872
rect 5046 -1448 5080 -872
rect 5164 -1448 5198 -872
rect 5282 -1448 5316 -872
rect 5400 -1448 5434 -872
rect 5518 -1448 5552 -872
rect 5636 -1448 5670 -872
rect 5754 -1448 5788 -872
rect 5872 -1448 5906 -872
rect 5990 -1448 6024 -872
rect 6108 -1448 6142 -872
rect 6226 -1448 6260 -872
rect 6344 -1448 6378 -872
rect 6462 -1448 6496 -872
rect 6580 -1448 6614 -872
rect 6698 -1448 6732 -872
rect 6816 -1448 6850 -872
rect 6934 -1448 6968 -872
rect 7052 -1448 7086 -872
rect 7170 -1448 7204 -872
rect 7288 -1448 7322 -872
rect 7406 -1448 7440 -872
rect 7524 -1448 7558 -872
rect 7642 -1448 7676 -872
rect 7760 -1448 7794 -872
rect 7878 -1448 7912 -872
rect 7996 -1448 8030 -872
rect 8114 -1448 8148 -872
rect 8232 -1448 8266 -872
rect 8350 -1448 8384 -872
rect 8468 -1448 8502 -872
rect 8586 -1448 8620 -872
rect 8704 -1448 8738 -872
rect 8822 -1448 8856 -872
rect 8940 -1448 8974 -872
rect 9058 -1448 9092 -872
rect 9176 -1448 9210 -872
rect 9294 -1448 9328 -872
rect 9412 -1448 9446 -872
rect 9530 -1448 9564 -872
rect 9648 -1448 9682 -872
rect 9766 -1448 9800 -872
rect 9884 -1448 9918 -872
rect 10002 -1448 10036 -872
rect 10120 -1448 10154 -872
rect 10238 -1448 10272 -872
rect 10356 -1448 10390 -872
rect 10474 -1448 10508 -872
rect 10592 -1448 10626 -872
rect 10710 -1448 10744 -872
rect 4810 -2284 4844 -1708
rect 4928 -2284 4962 -1708
rect 5046 -2284 5080 -1708
rect 5164 -2284 5198 -1708
rect 5282 -2284 5316 -1708
rect 5400 -2284 5434 -1708
rect 5518 -2284 5552 -1708
rect 5636 -2284 5670 -1708
rect 5754 -2284 5788 -1708
rect 5872 -2284 5906 -1708
rect 5990 -2284 6024 -1708
rect 6108 -2284 6142 -1708
rect 6226 -2284 6260 -1708
rect 6344 -2284 6378 -1708
rect 6462 -2284 6496 -1708
rect 6580 -2284 6614 -1708
rect 6698 -2284 6732 -1708
rect 6816 -2284 6850 -1708
rect 6934 -2284 6968 -1708
rect 7052 -2284 7086 -1708
rect 7170 -2284 7204 -1708
rect 7288 -2284 7322 -1708
rect 7406 -2284 7440 -1708
rect 7524 -2284 7558 -1708
rect 7642 -2284 7676 -1708
rect 7760 -2284 7794 -1708
rect 7878 -2284 7912 -1708
rect 7996 -2284 8030 -1708
rect 8114 -2284 8148 -1708
rect 8232 -2284 8266 -1708
rect 8350 -2284 8384 -1708
rect 8468 -2284 8502 -1708
rect 8586 -2284 8620 -1708
rect 8704 -2284 8738 -1708
rect 8822 -2284 8856 -1708
rect 8940 -2284 8974 -1708
rect 9058 -2284 9092 -1708
rect 9176 -2284 9210 -1708
rect 9294 -2284 9328 -1708
rect 9412 -2284 9446 -1708
rect 9530 -2284 9564 -1708
rect 9648 -2284 9682 -1708
rect 9766 -2284 9800 -1708
rect 9884 -2284 9918 -1708
rect 10002 -2284 10036 -1708
rect 10120 -2284 10154 -1708
rect 10238 -2284 10272 -1708
rect 10356 -2284 10390 -1708
rect 10474 -2284 10508 -1708
rect 10592 -2284 10626 -1708
rect 10710 -2284 10744 -1708
rect 4810 -3498 4844 -2922
rect 4928 -3498 4962 -2922
rect 5046 -3498 5080 -2922
rect 5164 -3498 5198 -2922
rect 5282 -3498 5316 -2922
rect 5400 -3498 5434 -2922
rect 5518 -3498 5552 -2922
rect 5636 -3498 5670 -2922
rect 5754 -3498 5788 -2922
rect 5872 -3498 5906 -2922
rect 5990 -3498 6024 -2922
rect 6108 -3498 6142 -2922
rect 6226 -3498 6260 -2922
rect 6344 -3498 6378 -2922
rect 6462 -3498 6496 -2922
rect 6580 -3498 6614 -2922
rect 6698 -3498 6732 -2922
rect 6816 -3498 6850 -2922
rect 6934 -3498 6968 -2922
rect 7052 -3498 7086 -2922
rect 7170 -3498 7204 -2922
rect 7288 -3498 7322 -2922
rect 7406 -3498 7440 -2922
rect 7524 -3498 7558 -2922
rect 7642 -3498 7676 -2922
rect 7760 -3498 7794 -2922
rect 7878 -3498 7912 -2922
rect 7996 -3498 8030 -2922
rect 8114 -3498 8148 -2922
rect 8232 -3498 8266 -2922
rect 8350 -3498 8384 -2922
rect 8468 -3498 8502 -2922
rect 8586 -3498 8620 -2922
rect 8704 -3498 8738 -2922
rect 8822 -3498 8856 -2922
rect 8940 -3498 8974 -2922
rect 9058 -3498 9092 -2922
rect 9176 -3498 9210 -2922
rect 9294 -3498 9328 -2922
rect 9412 -3498 9446 -2922
rect 9530 -3498 9564 -2922
rect 9648 -3498 9682 -2922
rect 9766 -3498 9800 -2922
rect 9884 -3498 9918 -2922
rect 10002 -3498 10036 -2922
rect 10120 -3498 10154 -2922
rect 10238 -3498 10272 -2922
rect 10356 -3498 10390 -2922
rect 10474 -3498 10508 -2922
rect 10592 -3498 10626 -2922
rect 10710 -3498 10744 -2922
rect 4810 -4334 4844 -3758
rect 4928 -4334 4962 -3758
rect 5046 -4334 5080 -3758
rect 5164 -4334 5198 -3758
rect 5282 -4334 5316 -3758
rect 5400 -4334 5434 -3758
rect 5518 -4334 5552 -3758
rect 5636 -4334 5670 -3758
rect 5754 -4334 5788 -3758
rect 5872 -4334 5906 -3758
rect 5990 -4334 6024 -3758
rect 6108 -4334 6142 -3758
rect 6226 -4334 6260 -3758
rect 6344 -4334 6378 -3758
rect 6462 -4334 6496 -3758
rect 6580 -4334 6614 -3758
rect 6698 -4334 6732 -3758
rect 6816 -4334 6850 -3758
rect 6934 -4334 6968 -3758
rect 7052 -4334 7086 -3758
rect 7170 -4334 7204 -3758
rect 7288 -4334 7322 -3758
rect 7406 -4334 7440 -3758
rect 7524 -4334 7558 -3758
rect 7642 -4334 7676 -3758
rect 7760 -4334 7794 -3758
rect 7878 -4334 7912 -3758
rect 7996 -4334 8030 -3758
rect 8114 -4334 8148 -3758
rect 8232 -4334 8266 -3758
rect 8350 -4334 8384 -3758
rect 8468 -4334 8502 -3758
rect 8586 -4334 8620 -3758
rect 8704 -4334 8738 -3758
rect 8822 -4334 8856 -3758
rect 8940 -4334 8974 -3758
rect 9058 -4334 9092 -3758
rect 9176 -4334 9210 -3758
rect 9294 -4334 9328 -3758
rect 9412 -4334 9446 -3758
rect 9530 -4334 9564 -3758
rect 9648 -4334 9682 -3758
rect 9766 -4334 9800 -3758
rect 9884 -4334 9918 -3758
rect 10002 -4334 10036 -3758
rect 10120 -4334 10154 -3758
rect 10238 -4334 10272 -3758
rect 10356 -4334 10390 -3758
rect 10474 -4334 10508 -3758
rect 10592 -4334 10626 -3758
rect 10710 -4334 10744 -3758
rect 5754 -5548 5788 -4972
rect 5872 -5548 5906 -4972
rect 5990 -5548 6024 -4972
rect 6108 -5548 6142 -4972
rect 9058 -5548 9092 -4972
rect 9176 -5548 9210 -4972
rect 9294 -5548 9328 -4972
rect 9412 -5548 9446 -4972
rect 9530 -5548 9564 -4972
rect 9648 -5548 9682 -4972
rect 9766 -5548 9800 -4972
rect 9884 -5548 9918 -4972
rect 10002 -5548 10036 -4972
rect 10120 -5548 10154 -4972
rect 10238 -5548 10272 -4972
rect 10356 -5548 10390 -4972
rect 5754 -6384 5788 -5808
rect 5872 -6384 5906 -5808
rect 5990 -6384 6024 -5808
rect 6108 -6384 6142 -5808
rect 9058 -6384 9092 -5808
rect 9176 -6384 9210 -5808
rect 9294 -6384 9328 -5808
rect 9412 -6384 9446 -5808
rect 9530 -6384 9564 -5808
rect 9648 -6384 9682 -5808
rect 9766 -6384 9800 -5808
rect 9884 -6384 9918 -5808
rect 10002 -6384 10036 -5808
rect 10120 -6384 10154 -5808
rect 10238 -6384 10272 -5808
rect 10356 -6384 10390 -5808
<< psubdiff >>
rect 10737 -7225 10777 -7191
rect 11053 -7225 11093 -7191
rect 11369 -7225 11409 -7191
rect 11685 -7225 11725 -7191
rect 12001 -7225 12041 -7191
rect 12317 -7225 12357 -7191
rect 10737 -7287 10771 -7225
rect 10421 -7640 10455 -7437
rect 11053 -7287 11087 -7225
rect 10737 -7649 10771 -7593
rect 11369 -7287 11403 -7225
rect 11053 -7649 11087 -7593
rect 11685 -7287 11719 -7225
rect 11369 -7649 11403 -7593
rect 12001 -7287 12035 -7225
rect 11685 -7649 11719 -7593
rect 12317 -7287 12351 -7225
rect 12001 -7649 12035 -7593
rect 12317 -7649 12351 -7593
rect 10440 -7689 12310 -7655
rect 5583 -8831 5697 -8797
rect 4056 -8865 5697 -8831
rect 4056 -8871 5750 -8865
rect 4056 -8905 4080 -8871
rect 4114 -8905 4152 -8871
rect 4186 -8905 4234 -8871
rect 4268 -8905 4306 -8871
rect 4340 -8905 4388 -8871
rect 4422 -8905 4460 -8871
rect 4494 -8905 4542 -8871
rect 4576 -8905 4614 -8871
rect 4648 -8905 4696 -8871
rect 4730 -8905 4768 -8871
rect 4802 -8905 4850 -8871
rect 4884 -8905 4922 -8871
rect 4956 -8905 5004 -8871
rect 5038 -8905 5076 -8871
rect 5110 -8905 5158 -8871
rect 5192 -8905 5230 -8871
rect 5264 -8905 5312 -8871
rect 5346 -8905 5384 -8871
rect 5418 -8905 5466 -8871
rect 5500 -8905 5538 -8871
rect 5572 -8905 5620 -8871
rect 5654 -8905 5692 -8871
rect 5726 -8877 5750 -8871
rect 5726 -8905 12064 -8877
rect 4056 -8945 12064 -8905
rect 4056 -8979 4080 -8945
rect 4114 -8979 4152 -8945
rect 4186 -8979 4234 -8945
rect 4268 -8979 4306 -8945
rect 4340 -8979 4388 -8945
rect 4422 -8979 4460 -8945
rect 4494 -8979 4542 -8945
rect 4576 -8979 4614 -8945
rect 4648 -8979 4696 -8945
rect 4730 -8979 4768 -8945
rect 4802 -8979 4850 -8945
rect 4884 -8979 4922 -8945
rect 4956 -8979 5004 -8945
rect 5038 -8979 5076 -8945
rect 5110 -8979 5158 -8945
rect 5192 -8979 5230 -8945
rect 5264 -8979 5312 -8945
rect 5346 -8979 5384 -8945
rect 5418 -8979 5466 -8945
rect 5500 -8979 5538 -8945
rect 5572 -8979 5620 -8945
rect 5654 -8979 5692 -8945
rect 5726 -8979 5774 -8945
rect 5808 -8979 5846 -8945
rect 5880 -8979 5928 -8945
rect 5962 -8979 6000 -8945
rect 6034 -8979 6082 -8945
rect 6116 -8979 6154 -8945
rect 6188 -8979 6236 -8945
rect 6270 -8979 6308 -8945
rect 6342 -8979 6390 -8945
rect 6424 -8979 6462 -8945
rect 6496 -8979 6544 -8945
rect 6578 -8979 6616 -8945
rect 6650 -8979 6698 -8945
rect 6732 -8979 6770 -8945
rect 6804 -8979 6852 -8945
rect 6886 -8979 6924 -8945
rect 6958 -8979 7006 -8945
rect 7040 -8979 7078 -8945
rect 7112 -8979 7160 -8945
rect 7194 -8979 7232 -8945
rect 7266 -8979 7314 -8945
rect 7348 -8979 7386 -8945
rect 7420 -8979 7468 -8945
rect 7502 -8979 7540 -8945
rect 7574 -8979 7622 -8945
rect 7656 -8979 7694 -8945
rect 7728 -8979 7776 -8945
rect 7810 -8979 7848 -8945
rect 7882 -8979 7930 -8945
rect 7964 -8979 8002 -8945
rect 8036 -8979 8084 -8945
rect 8118 -8979 8156 -8945
rect 8190 -8979 8238 -8945
rect 8272 -8979 8310 -8945
rect 8344 -8979 8392 -8945
rect 8426 -8979 8464 -8945
rect 8498 -8979 8546 -8945
rect 8580 -8979 8618 -8945
rect 8652 -8979 8700 -8945
rect 8734 -8979 8772 -8945
rect 8806 -8979 8854 -8945
rect 8888 -8979 8926 -8945
rect 8960 -8979 9008 -8945
rect 9042 -8979 9080 -8945
rect 9114 -8979 9162 -8945
rect 9196 -8979 9234 -8945
rect 9268 -8979 9316 -8945
rect 9350 -8979 9388 -8945
rect 9422 -8979 9470 -8945
rect 9504 -8979 9542 -8945
rect 9576 -8979 9624 -8945
rect 9658 -8979 9696 -8945
rect 9730 -8979 9778 -8945
rect 9812 -8979 9850 -8945
rect 9884 -8979 9932 -8945
rect 9966 -8979 10004 -8945
rect 10038 -8979 10086 -8945
rect 10120 -8979 10158 -8945
rect 10192 -8979 10240 -8945
rect 10274 -8979 10312 -8945
rect 10346 -8979 10394 -8945
rect 10428 -8979 10466 -8945
rect 10500 -8979 10548 -8945
rect 10582 -8979 10620 -8945
rect 10654 -8979 10702 -8945
rect 10736 -8979 10774 -8945
rect 10808 -8979 10856 -8945
rect 10890 -8979 10928 -8945
rect 10962 -8979 11010 -8945
rect 11044 -8979 11082 -8945
rect 11116 -8979 11164 -8945
rect 11198 -8979 11236 -8945
rect 11270 -8979 11318 -8945
rect 11352 -8979 11390 -8945
rect 11424 -8979 11472 -8945
rect 11506 -8979 11544 -8945
rect 11578 -8979 11626 -8945
rect 11660 -8979 11698 -8945
rect 11732 -8979 11780 -8945
rect 11814 -8979 11852 -8945
rect 11886 -8979 11934 -8945
rect 11968 -8979 12006 -8945
rect 12040 -8979 12064 -8945
rect 4056 -9019 12064 -8979
rect 4056 -9053 4080 -9019
rect 4114 -9053 4152 -9019
rect 4186 -9053 4234 -9019
rect 4268 -9053 4306 -9019
rect 4340 -9053 4388 -9019
rect 4422 -9053 4460 -9019
rect 4494 -9053 4542 -9019
rect 4576 -9053 4614 -9019
rect 4648 -9053 4696 -9019
rect 4730 -9053 4768 -9019
rect 4802 -9053 4850 -9019
rect 4884 -9053 4922 -9019
rect 4956 -9053 5004 -9019
rect 5038 -9053 5076 -9019
rect 5110 -9053 5158 -9019
rect 5192 -9053 5230 -9019
rect 5264 -9053 5312 -9019
rect 5346 -9053 5384 -9019
rect 5418 -9053 5466 -9019
rect 5500 -9053 5538 -9019
rect 5572 -9053 5620 -9019
rect 5654 -9053 5692 -9019
rect 5726 -9053 5774 -9019
rect 5808 -9053 5846 -9019
rect 5880 -9053 5928 -9019
rect 5962 -9053 6000 -9019
rect 6034 -9053 6082 -9019
rect 6116 -9053 6154 -9019
rect 6188 -9053 6236 -9019
rect 6270 -9053 6308 -9019
rect 6342 -9053 6390 -9019
rect 6424 -9053 6462 -9019
rect 6496 -9053 6544 -9019
rect 6578 -9053 6616 -9019
rect 6650 -9053 6698 -9019
rect 6732 -9053 6770 -9019
rect 6804 -9053 6852 -9019
rect 6886 -9053 6924 -9019
rect 6958 -9053 7006 -9019
rect 7040 -9053 7078 -9019
rect 7112 -9053 7160 -9019
rect 7194 -9053 7232 -9019
rect 7266 -9053 7314 -9019
rect 7348 -9053 7386 -9019
rect 7420 -9053 7468 -9019
rect 7502 -9053 7540 -9019
rect 7574 -9053 7622 -9019
rect 7656 -9053 7694 -9019
rect 7728 -9053 7776 -9019
rect 7810 -9053 7848 -9019
rect 7882 -9053 7930 -9019
rect 7964 -9053 8002 -9019
rect 8036 -9053 8084 -9019
rect 8118 -9053 8156 -9019
rect 8190 -9053 8238 -9019
rect 8272 -9053 8310 -9019
rect 8344 -9053 8392 -9019
rect 8426 -9053 8464 -9019
rect 8498 -9053 8546 -9019
rect 8580 -9053 8618 -9019
rect 8652 -9053 8700 -9019
rect 8734 -9053 8772 -9019
rect 8806 -9053 8854 -9019
rect 8888 -9053 8926 -9019
rect 8960 -9053 9008 -9019
rect 9042 -9053 9080 -9019
rect 9114 -9053 9162 -9019
rect 9196 -9053 9234 -9019
rect 9268 -9053 9316 -9019
rect 9350 -9053 9388 -9019
rect 9422 -9053 9470 -9019
rect 9504 -9053 9542 -9019
rect 9576 -9053 9624 -9019
rect 9658 -9053 9696 -9019
rect 9730 -9053 9778 -9019
rect 9812 -9053 9850 -9019
rect 9884 -9053 9932 -9019
rect 9966 -9053 10004 -9019
rect 10038 -9053 10086 -9019
rect 10120 -9053 10158 -9019
rect 10192 -9053 10240 -9019
rect 10274 -9053 10312 -9019
rect 10346 -9053 10394 -9019
rect 10428 -9053 10466 -9019
rect 10500 -9053 10548 -9019
rect 10582 -9053 10620 -9019
rect 10654 -9053 10702 -9019
rect 10736 -9053 10774 -9019
rect 10808 -9053 10856 -9019
rect 10890 -9053 10928 -9019
rect 10962 -9053 11010 -9019
rect 11044 -9053 11082 -9019
rect 11116 -9053 11164 -9019
rect 11198 -9053 11236 -9019
rect 11270 -9053 11318 -9019
rect 11352 -9053 11390 -9019
rect 11424 -9053 11472 -9019
rect 11506 -9053 11544 -9019
rect 11578 -9053 11626 -9019
rect 11660 -9053 11698 -9019
rect 11732 -9053 11780 -9019
rect 11814 -9053 11852 -9019
rect 11886 -9053 11934 -9019
rect 11968 -9053 12006 -9019
rect 12040 -9053 12064 -9019
rect 4056 -9093 12064 -9053
rect 4056 -9127 4080 -9093
rect 4114 -9127 4152 -9093
rect 4186 -9127 4234 -9093
rect 4268 -9127 4306 -9093
rect 4340 -9127 4388 -9093
rect 4422 -9127 4460 -9093
rect 4494 -9127 4542 -9093
rect 4576 -9127 4614 -9093
rect 4648 -9127 4696 -9093
rect 4730 -9127 4768 -9093
rect 4802 -9127 4850 -9093
rect 4884 -9127 4922 -9093
rect 4956 -9127 5004 -9093
rect 5038 -9127 5076 -9093
rect 5110 -9127 5158 -9093
rect 5192 -9127 5230 -9093
rect 5264 -9127 5312 -9093
rect 5346 -9127 5384 -9093
rect 5418 -9127 5466 -9093
rect 5500 -9127 5538 -9093
rect 5572 -9127 5620 -9093
rect 5654 -9127 5692 -9093
rect 5726 -9127 5774 -9093
rect 5808 -9127 5846 -9093
rect 5880 -9127 5928 -9093
rect 5962 -9127 6000 -9093
rect 6034 -9127 6082 -9093
rect 6116 -9127 6154 -9093
rect 6188 -9127 6236 -9093
rect 6270 -9127 6308 -9093
rect 6342 -9127 6390 -9093
rect 6424 -9127 6462 -9093
rect 6496 -9127 6544 -9093
rect 6578 -9127 6616 -9093
rect 6650 -9127 6698 -9093
rect 6732 -9127 6770 -9093
rect 6804 -9127 6852 -9093
rect 6886 -9127 6924 -9093
rect 6958 -9127 7006 -9093
rect 7040 -9127 7078 -9093
rect 7112 -9127 7160 -9093
rect 7194 -9127 7232 -9093
rect 7266 -9127 7314 -9093
rect 7348 -9127 7386 -9093
rect 7420 -9127 7468 -9093
rect 7502 -9127 7540 -9093
rect 7574 -9127 7622 -9093
rect 7656 -9127 7694 -9093
rect 7728 -9127 7776 -9093
rect 7810 -9127 7848 -9093
rect 7882 -9127 7930 -9093
rect 7964 -9127 8002 -9093
rect 8036 -9127 8084 -9093
rect 8118 -9127 8156 -9093
rect 8190 -9127 8238 -9093
rect 8272 -9127 8310 -9093
rect 8344 -9127 8392 -9093
rect 8426 -9127 8464 -9093
rect 8498 -9127 8546 -9093
rect 8580 -9127 8618 -9093
rect 8652 -9127 8700 -9093
rect 8734 -9127 8772 -9093
rect 8806 -9127 8854 -9093
rect 8888 -9127 8926 -9093
rect 8960 -9127 9008 -9093
rect 9042 -9127 9080 -9093
rect 9114 -9127 9162 -9093
rect 9196 -9127 9234 -9093
rect 9268 -9127 9316 -9093
rect 9350 -9127 9388 -9093
rect 9422 -9127 9470 -9093
rect 9504 -9127 9542 -9093
rect 9576 -9127 9624 -9093
rect 9658 -9127 9696 -9093
rect 9730 -9127 9778 -9093
rect 9812 -9127 9850 -9093
rect 9884 -9127 9932 -9093
rect 9966 -9127 10004 -9093
rect 10038 -9127 10086 -9093
rect 10120 -9127 10158 -9093
rect 10192 -9127 10240 -9093
rect 10274 -9127 10312 -9093
rect 10346 -9127 10394 -9093
rect 10428 -9127 10466 -9093
rect 10500 -9127 10548 -9093
rect 10582 -9127 10620 -9093
rect 10654 -9127 10702 -9093
rect 10736 -9127 10774 -9093
rect 10808 -9127 10856 -9093
rect 10890 -9127 10928 -9093
rect 10962 -9127 11010 -9093
rect 11044 -9127 11082 -9093
rect 11116 -9127 11164 -9093
rect 11198 -9127 11236 -9093
rect 11270 -9127 11318 -9093
rect 11352 -9127 11390 -9093
rect 11424 -9127 11472 -9093
rect 11506 -9127 11544 -9093
rect 11578 -9127 11626 -9093
rect 11660 -9127 11698 -9093
rect 11732 -9127 11780 -9093
rect 11814 -9127 11852 -9093
rect 11886 -9127 11934 -9093
rect 11968 -9127 12006 -9093
rect 12040 -9127 12064 -9093
rect 4056 -9167 12064 -9127
rect 4056 -9201 4080 -9167
rect 4114 -9201 4152 -9167
rect 4186 -9201 4234 -9167
rect 4268 -9201 4306 -9167
rect 4340 -9201 4388 -9167
rect 4422 -9201 4460 -9167
rect 4494 -9201 4542 -9167
rect 4576 -9201 4614 -9167
rect 4648 -9201 4696 -9167
rect 4730 -9201 4768 -9167
rect 4802 -9201 4850 -9167
rect 4884 -9201 4922 -9167
rect 4956 -9201 5004 -9167
rect 5038 -9201 5076 -9167
rect 5110 -9201 5158 -9167
rect 5192 -9201 5230 -9167
rect 5264 -9201 5312 -9167
rect 5346 -9201 5384 -9167
rect 5418 -9201 5466 -9167
rect 5500 -9201 5538 -9167
rect 5572 -9201 5620 -9167
rect 5654 -9201 5692 -9167
rect 5726 -9201 5774 -9167
rect 5808 -9201 5846 -9167
rect 5880 -9201 5928 -9167
rect 5962 -9201 6000 -9167
rect 6034 -9201 6082 -9167
rect 6116 -9201 6154 -9167
rect 6188 -9201 6236 -9167
rect 6270 -9201 6308 -9167
rect 6342 -9201 6390 -9167
rect 6424 -9201 6462 -9167
rect 6496 -9201 6544 -9167
rect 6578 -9201 6616 -9167
rect 6650 -9201 6698 -9167
rect 6732 -9201 6770 -9167
rect 6804 -9201 6852 -9167
rect 6886 -9201 6924 -9167
rect 6958 -9201 7006 -9167
rect 7040 -9201 7078 -9167
rect 7112 -9201 7160 -9167
rect 7194 -9201 7232 -9167
rect 7266 -9201 7314 -9167
rect 7348 -9201 7386 -9167
rect 7420 -9201 7468 -9167
rect 7502 -9201 7540 -9167
rect 7574 -9201 7622 -9167
rect 7656 -9201 7694 -9167
rect 7728 -9201 7776 -9167
rect 7810 -9201 7848 -9167
rect 7882 -9201 7930 -9167
rect 7964 -9201 8002 -9167
rect 8036 -9201 8084 -9167
rect 8118 -9201 8156 -9167
rect 8190 -9201 8238 -9167
rect 8272 -9201 8310 -9167
rect 8344 -9201 8392 -9167
rect 8426 -9201 8464 -9167
rect 8498 -9201 8546 -9167
rect 8580 -9201 8618 -9167
rect 8652 -9201 8700 -9167
rect 8734 -9201 8772 -9167
rect 8806 -9201 8854 -9167
rect 8888 -9201 8926 -9167
rect 8960 -9201 9008 -9167
rect 9042 -9201 9080 -9167
rect 9114 -9201 9162 -9167
rect 9196 -9201 9234 -9167
rect 9268 -9201 9316 -9167
rect 9350 -9201 9388 -9167
rect 9422 -9201 9470 -9167
rect 9504 -9201 9542 -9167
rect 9576 -9201 9624 -9167
rect 9658 -9201 9696 -9167
rect 9730 -9201 9778 -9167
rect 9812 -9201 9850 -9167
rect 9884 -9201 9932 -9167
rect 9966 -9201 10004 -9167
rect 10038 -9201 10086 -9167
rect 10120 -9201 10158 -9167
rect 10192 -9201 10240 -9167
rect 10274 -9201 10312 -9167
rect 10346 -9201 10394 -9167
rect 10428 -9201 10466 -9167
rect 10500 -9201 10548 -9167
rect 10582 -9201 10620 -9167
rect 10654 -9201 10702 -9167
rect 10736 -9201 10774 -9167
rect 10808 -9201 10856 -9167
rect 10890 -9201 10928 -9167
rect 10962 -9201 11010 -9167
rect 11044 -9201 11082 -9167
rect 11116 -9201 11164 -9167
rect 11198 -9201 11236 -9167
rect 11270 -9201 11318 -9167
rect 11352 -9201 11390 -9167
rect 11424 -9201 11472 -9167
rect 11506 -9201 11544 -9167
rect 11578 -9201 11626 -9167
rect 11660 -9201 11698 -9167
rect 11732 -9201 11780 -9167
rect 11814 -9201 11852 -9167
rect 11886 -9201 11934 -9167
rect 11968 -9201 12006 -9167
rect 12040 -9201 12064 -9167
rect 4056 -9241 12064 -9201
rect 4056 -9275 4080 -9241
rect 4114 -9275 4152 -9241
rect 4186 -9275 4234 -9241
rect 4268 -9275 4306 -9241
rect 4340 -9275 4388 -9241
rect 4422 -9275 4460 -9241
rect 4494 -9275 4542 -9241
rect 4576 -9275 4614 -9241
rect 4648 -9275 4696 -9241
rect 4730 -9275 4768 -9241
rect 4802 -9275 4850 -9241
rect 4884 -9275 4922 -9241
rect 4956 -9275 5004 -9241
rect 5038 -9275 5076 -9241
rect 5110 -9275 5158 -9241
rect 5192 -9275 5230 -9241
rect 5264 -9275 5312 -9241
rect 5346 -9275 5384 -9241
rect 5418 -9275 5466 -9241
rect 5500 -9275 5538 -9241
rect 5572 -9275 5620 -9241
rect 5654 -9275 5692 -9241
rect 5726 -9275 5774 -9241
rect 5808 -9275 5846 -9241
rect 5880 -9275 5928 -9241
rect 5962 -9275 6000 -9241
rect 6034 -9275 6082 -9241
rect 6116 -9275 6154 -9241
rect 6188 -9275 6236 -9241
rect 6270 -9275 6308 -9241
rect 6342 -9275 6390 -9241
rect 6424 -9275 6462 -9241
rect 6496 -9275 6544 -9241
rect 6578 -9275 6616 -9241
rect 6650 -9275 6698 -9241
rect 6732 -9275 6770 -9241
rect 6804 -9275 6852 -9241
rect 6886 -9275 6924 -9241
rect 6958 -9275 7006 -9241
rect 7040 -9275 7078 -9241
rect 7112 -9275 7160 -9241
rect 7194 -9275 7232 -9241
rect 7266 -9275 7314 -9241
rect 7348 -9275 7386 -9241
rect 7420 -9275 7468 -9241
rect 7502 -9275 7540 -9241
rect 7574 -9275 7622 -9241
rect 7656 -9275 7694 -9241
rect 7728 -9275 7776 -9241
rect 7810 -9275 7848 -9241
rect 7882 -9275 7930 -9241
rect 7964 -9275 8002 -9241
rect 8036 -9275 8084 -9241
rect 8118 -9275 8156 -9241
rect 8190 -9275 8238 -9241
rect 8272 -9275 8310 -9241
rect 8344 -9275 8392 -9241
rect 8426 -9275 8464 -9241
rect 8498 -9275 8546 -9241
rect 8580 -9275 8618 -9241
rect 8652 -9275 8700 -9241
rect 8734 -9275 8772 -9241
rect 8806 -9275 8854 -9241
rect 8888 -9275 8926 -9241
rect 8960 -9275 9008 -9241
rect 9042 -9275 9080 -9241
rect 9114 -9275 9162 -9241
rect 9196 -9275 9234 -9241
rect 9268 -9275 9316 -9241
rect 9350 -9275 9388 -9241
rect 9422 -9275 9470 -9241
rect 9504 -9275 9542 -9241
rect 9576 -9275 9624 -9241
rect 9658 -9275 9696 -9241
rect 9730 -9275 9778 -9241
rect 9812 -9275 9850 -9241
rect 9884 -9275 9932 -9241
rect 9966 -9275 10004 -9241
rect 10038 -9275 10086 -9241
rect 10120 -9275 10158 -9241
rect 10192 -9275 10240 -9241
rect 10274 -9275 10312 -9241
rect 10346 -9275 10394 -9241
rect 10428 -9275 10466 -9241
rect 10500 -9275 10548 -9241
rect 10582 -9275 10620 -9241
rect 10654 -9275 10702 -9241
rect 10736 -9275 10774 -9241
rect 10808 -9275 10856 -9241
rect 10890 -9275 10928 -9241
rect 10962 -9275 11010 -9241
rect 11044 -9275 11082 -9241
rect 11116 -9275 11164 -9241
rect 11198 -9275 11236 -9241
rect 11270 -9275 11318 -9241
rect 11352 -9275 11390 -9241
rect 11424 -9275 11472 -9241
rect 11506 -9275 11544 -9241
rect 11578 -9275 11626 -9241
rect 11660 -9275 11698 -9241
rect 11732 -9275 11780 -9241
rect 11814 -9275 11852 -9241
rect 11886 -9275 11934 -9241
rect 11968 -9275 12006 -9241
rect 12040 -9275 12064 -9241
rect 4056 -9315 12064 -9275
rect 4056 -9349 4080 -9315
rect 4114 -9349 4152 -9315
rect 4186 -9349 4234 -9315
rect 4268 -9349 4306 -9315
rect 4340 -9349 4388 -9315
rect 4422 -9349 4460 -9315
rect 4494 -9349 4542 -9315
rect 4576 -9349 4614 -9315
rect 4648 -9349 4696 -9315
rect 4730 -9349 4768 -9315
rect 4802 -9349 4850 -9315
rect 4884 -9349 4922 -9315
rect 4956 -9349 5004 -9315
rect 5038 -9349 5076 -9315
rect 5110 -9349 5158 -9315
rect 5192 -9349 5230 -9315
rect 5264 -9349 5312 -9315
rect 5346 -9349 5384 -9315
rect 5418 -9349 5466 -9315
rect 5500 -9349 5538 -9315
rect 5572 -9349 5620 -9315
rect 5654 -9349 5692 -9315
rect 5726 -9349 5774 -9315
rect 5808 -9349 5846 -9315
rect 5880 -9349 5928 -9315
rect 5962 -9349 6000 -9315
rect 6034 -9349 6082 -9315
rect 6116 -9349 6154 -9315
rect 6188 -9349 6236 -9315
rect 6270 -9349 6308 -9315
rect 6342 -9349 6390 -9315
rect 6424 -9349 6462 -9315
rect 6496 -9349 6544 -9315
rect 6578 -9349 6616 -9315
rect 6650 -9349 6698 -9315
rect 6732 -9349 6770 -9315
rect 6804 -9349 6852 -9315
rect 6886 -9349 6924 -9315
rect 6958 -9349 7006 -9315
rect 7040 -9349 7078 -9315
rect 7112 -9349 7160 -9315
rect 7194 -9349 7232 -9315
rect 7266 -9349 7314 -9315
rect 7348 -9349 7386 -9315
rect 7420 -9349 7468 -9315
rect 7502 -9349 7540 -9315
rect 7574 -9349 7622 -9315
rect 7656 -9349 7694 -9315
rect 7728 -9349 7776 -9315
rect 7810 -9349 7848 -9315
rect 7882 -9349 7930 -9315
rect 7964 -9349 8002 -9315
rect 8036 -9349 8084 -9315
rect 8118 -9349 8156 -9315
rect 8190 -9349 8238 -9315
rect 8272 -9349 8310 -9315
rect 8344 -9349 8392 -9315
rect 8426 -9349 8464 -9315
rect 8498 -9349 8546 -9315
rect 8580 -9349 8618 -9315
rect 8652 -9349 8700 -9315
rect 8734 -9349 8772 -9315
rect 8806 -9349 8854 -9315
rect 8888 -9349 8926 -9315
rect 8960 -9349 9008 -9315
rect 9042 -9349 9080 -9315
rect 9114 -9349 9162 -9315
rect 9196 -9349 9234 -9315
rect 9268 -9349 9316 -9315
rect 9350 -9349 9388 -9315
rect 9422 -9349 9470 -9315
rect 9504 -9349 9542 -9315
rect 9576 -9349 9624 -9315
rect 9658 -9349 9696 -9315
rect 9730 -9349 9778 -9315
rect 9812 -9349 9850 -9315
rect 9884 -9349 9932 -9315
rect 9966 -9349 10004 -9315
rect 10038 -9349 10086 -9315
rect 10120 -9349 10158 -9315
rect 10192 -9349 10240 -9315
rect 10274 -9349 10312 -9315
rect 10346 -9349 10394 -9315
rect 10428 -9349 10466 -9315
rect 10500 -9349 10548 -9315
rect 10582 -9349 10620 -9315
rect 10654 -9349 10702 -9315
rect 10736 -9349 10774 -9315
rect 10808 -9349 10856 -9315
rect 10890 -9349 10928 -9315
rect 10962 -9349 11010 -9315
rect 11044 -9349 11082 -9315
rect 11116 -9349 11164 -9315
rect 11198 -9349 11236 -9315
rect 11270 -9349 11318 -9315
rect 11352 -9349 11390 -9315
rect 11424 -9349 11472 -9315
rect 11506 -9349 11544 -9315
rect 11578 -9349 11626 -9315
rect 11660 -9349 11698 -9315
rect 11732 -9349 11780 -9315
rect 11814 -9349 11852 -9315
rect 11886 -9349 11934 -9315
rect 11968 -9349 12006 -9315
rect 12040 -9349 12064 -9315
rect 4056 -9389 12064 -9349
rect 4056 -9423 4080 -9389
rect 4114 -9423 4152 -9389
rect 4186 -9423 4234 -9389
rect 4268 -9423 4306 -9389
rect 4340 -9423 4388 -9389
rect 4422 -9423 4460 -9389
rect 4494 -9423 4542 -9389
rect 4576 -9423 4614 -9389
rect 4648 -9423 4696 -9389
rect 4730 -9423 4768 -9389
rect 4802 -9423 4850 -9389
rect 4884 -9423 4922 -9389
rect 4956 -9423 5004 -9389
rect 5038 -9423 5076 -9389
rect 5110 -9423 5158 -9389
rect 5192 -9423 5230 -9389
rect 5264 -9423 5312 -9389
rect 5346 -9423 5384 -9389
rect 5418 -9423 5466 -9389
rect 5500 -9423 5538 -9389
rect 5572 -9423 5620 -9389
rect 5654 -9423 5692 -9389
rect 5726 -9423 5774 -9389
rect 5808 -9423 5846 -9389
rect 5880 -9423 5928 -9389
rect 5962 -9423 6000 -9389
rect 6034 -9423 6082 -9389
rect 6116 -9423 6154 -9389
rect 6188 -9423 6236 -9389
rect 6270 -9423 6308 -9389
rect 6342 -9423 6390 -9389
rect 6424 -9423 6462 -9389
rect 6496 -9423 6544 -9389
rect 6578 -9423 6616 -9389
rect 6650 -9423 6698 -9389
rect 6732 -9423 6770 -9389
rect 6804 -9423 6852 -9389
rect 6886 -9423 6924 -9389
rect 6958 -9423 7006 -9389
rect 7040 -9423 7078 -9389
rect 7112 -9423 7160 -9389
rect 7194 -9423 7232 -9389
rect 7266 -9423 7314 -9389
rect 7348 -9423 7386 -9389
rect 7420 -9423 7468 -9389
rect 7502 -9423 7540 -9389
rect 7574 -9423 7622 -9389
rect 7656 -9423 7694 -9389
rect 7728 -9423 7776 -9389
rect 7810 -9423 7848 -9389
rect 7882 -9423 7930 -9389
rect 7964 -9423 8002 -9389
rect 8036 -9423 8084 -9389
rect 8118 -9423 8156 -9389
rect 8190 -9423 8238 -9389
rect 8272 -9423 8310 -9389
rect 8344 -9423 8392 -9389
rect 8426 -9423 8464 -9389
rect 8498 -9423 8546 -9389
rect 8580 -9423 8618 -9389
rect 8652 -9423 8700 -9389
rect 8734 -9423 8772 -9389
rect 8806 -9423 8854 -9389
rect 8888 -9423 8926 -9389
rect 8960 -9423 9008 -9389
rect 9042 -9423 9080 -9389
rect 9114 -9423 9162 -9389
rect 9196 -9423 9234 -9389
rect 9268 -9423 9316 -9389
rect 9350 -9423 9388 -9389
rect 9422 -9423 9470 -9389
rect 9504 -9423 9542 -9389
rect 9576 -9423 9624 -9389
rect 9658 -9423 9696 -9389
rect 9730 -9423 9778 -9389
rect 9812 -9423 9850 -9389
rect 9884 -9423 9932 -9389
rect 9966 -9423 10004 -9389
rect 10038 -9423 10086 -9389
rect 10120 -9423 10158 -9389
rect 10192 -9423 10240 -9389
rect 10274 -9423 10312 -9389
rect 10346 -9423 10394 -9389
rect 10428 -9423 10466 -9389
rect 10500 -9423 10548 -9389
rect 10582 -9423 10620 -9389
rect 10654 -9423 10702 -9389
rect 10736 -9423 10774 -9389
rect 10808 -9423 10856 -9389
rect 10890 -9423 10928 -9389
rect 10962 -9423 11010 -9389
rect 11044 -9423 11082 -9389
rect 11116 -9423 11164 -9389
rect 11198 -9423 11236 -9389
rect 11270 -9423 11318 -9389
rect 11352 -9423 11390 -9389
rect 11424 -9423 11472 -9389
rect 11506 -9423 11544 -9389
rect 11578 -9423 11626 -9389
rect 11660 -9423 11698 -9389
rect 11732 -9423 11780 -9389
rect 11814 -9423 11852 -9389
rect 11886 -9423 11934 -9389
rect 11968 -9423 12006 -9389
rect 12040 -9423 12064 -9389
rect 4056 -9577 12064 -9423
rect 4020 -9682 4060 -9678
rect 4019 -9712 4060 -9682
rect 4094 -9712 4134 -9678
rect 4168 -9712 4208 -9678
rect 4242 -9712 4282 -9678
rect 4316 -9712 4356 -9678
rect 4390 -9712 4430 -9678
rect 4464 -9712 4504 -9678
rect 4538 -9712 4578 -9678
rect 4612 -9712 4652 -9678
rect 4686 -9712 4726 -9678
rect 4760 -9712 4800 -9678
rect 4834 -9712 4874 -9678
rect 4908 -9712 4948 -9678
rect 4982 -9712 5022 -9678
rect 5056 -9712 5096 -9678
rect 5130 -9712 5170 -9678
rect 5204 -9712 5244 -9678
rect 5278 -9712 5318 -9678
rect 5352 -9712 5392 -9678
rect 5426 -9712 5466 -9678
rect 5500 -9712 5540 -9678
rect 5574 -9712 5614 -9678
rect 5648 -9712 5688 -9678
rect 5722 -9712 5762 -9678
rect 5796 -9712 5836 -9678
rect 5870 -9712 5910 -9678
rect 5944 -9712 5984 -9678
rect 6018 -9712 6058 -9678
rect 6092 -9712 6132 -9678
rect 6166 -9712 6206 -9678
rect 6240 -9712 6280 -9678
rect 6314 -9712 6354 -9678
rect 6388 -9712 6428 -9678
rect 6462 -9712 6502 -9678
rect 6536 -9712 6576 -9678
rect 6610 -9712 6650 -9678
rect 6684 -9712 6724 -9678
rect 6758 -9712 6798 -9678
rect 6832 -9712 6872 -9678
rect 6906 -9712 6946 -9678
rect 6980 -9712 7020 -9678
rect 7054 -9712 7094 -9678
rect 7128 -9712 7168 -9678
rect 7202 -9712 7242 -9678
rect 7276 -9712 7316 -9678
rect 7350 -9712 7390 -9678
rect 7424 -9712 7464 -9678
rect 7498 -9712 7538 -9678
rect 7572 -9712 7612 -9678
rect 7646 -9712 7686 -9678
rect 7720 -9712 7760 -9678
rect 7794 -9712 7834 -9678
rect 7868 -9712 7908 -9678
rect 7942 -9712 7982 -9678
rect 8016 -9712 8056 -9678
rect 8090 -9712 8130 -9678
rect 8164 -9712 8204 -9678
rect 8238 -9712 8278 -9678
rect 8312 -9712 8352 -9678
rect 8386 -9712 8426 -9678
rect 8460 -9712 8500 -9678
rect 8534 -9712 8574 -9678
rect 8608 -9712 8648 -9678
rect 8682 -9712 8722 -9678
rect 8756 -9712 8796 -9678
rect 8830 -9712 8870 -9678
rect 8904 -9712 8944 -9678
rect 8978 -9712 9018 -9678
rect 9052 -9712 9092 -9678
rect 9126 -9712 9166 -9678
rect 9200 -9712 9240 -9678
rect 9274 -9712 9314 -9678
rect 9348 -9712 9388 -9678
rect 9422 -9712 9462 -9678
rect 9496 -9712 9536 -9678
rect 9570 -9712 9610 -9678
rect 9644 -9712 9684 -9678
rect 9718 -9712 9758 -9678
rect 9792 -9712 9832 -9678
rect 9866 -9712 9906 -9678
rect 9940 -9712 9980 -9678
rect 10014 -9712 10054 -9678
rect 10088 -9712 10128 -9678
rect 10162 -9712 10202 -9678
rect 10236 -9712 10276 -9678
rect 10310 -9712 10350 -9678
rect 10384 -9712 10424 -9678
rect 10458 -9712 10498 -9678
rect 10532 -9712 10572 -9678
rect 10606 -9712 10646 -9678
rect 10680 -9712 10720 -9678
rect 10754 -9712 10794 -9678
rect 10828 -9712 10868 -9678
rect 10902 -9712 10942 -9678
rect 10976 -9712 11016 -9678
rect 11050 -9712 11090 -9678
rect 11124 -9712 11164 -9678
rect 11198 -9712 11238 -9678
rect 11272 -9712 11312 -9678
rect 11346 -9712 11386 -9678
rect 11420 -9712 11460 -9678
rect 11494 -9712 11534 -9678
rect 11568 -9712 11608 -9678
rect 11642 -9712 11682 -9678
rect 11716 -9712 11756 -9678
rect 11790 -9712 11830 -9678
rect 11864 -9712 11904 -9678
rect 11938 -9712 11978 -9678
rect 12012 -9712 12052 -9678
rect 12086 -9712 12126 -9678
rect 12160 -9712 12200 -9678
rect 12234 -9712 12274 -9678
rect 12308 -9712 12348 -9678
rect 12382 -9712 12422 -9678
rect 12456 -9712 12496 -9678
rect 12530 -9712 12570 -9678
rect 12604 -9712 12644 -9678
rect 12678 -9712 12718 -9678
rect 12752 -9712 12792 -9678
rect 12826 -9712 12866 -9678
rect 12900 -9712 12940 -9678
rect 12974 -9712 13014 -9678
rect 13048 -9712 13088 -9678
rect 13122 -9712 13162 -9678
rect 13196 -9712 13236 -9678
rect 13270 -9712 13310 -9678
rect 13344 -9712 13384 -9678
rect 13418 -9712 13458 -9678
rect 13492 -9712 13532 -9678
rect 13566 -9712 13606 -9678
rect 13640 -9712 13680 -9678
rect 13714 -9712 13754 -9678
rect 13788 -9712 13828 -9678
rect 13862 -9712 13902 -9678
rect 13936 -9712 13976 -9678
rect 14010 -9712 14050 -9678
rect 14084 -9712 14124 -9678
rect 14158 -9712 14198 -9678
rect 14232 -9712 14272 -9678
rect 14306 -9712 14346 -9678
rect 14380 -9712 14420 -9678
rect 14454 -9712 14494 -9678
rect 14528 -9712 14568 -9678
rect 14602 -9712 14642 -9678
rect 14676 -9712 14716 -9678
rect 14750 -9712 14790 -9678
rect 14824 -9712 14864 -9678
rect 14898 -9712 14938 -9678
rect 14972 -9712 15012 -9678
rect 15046 -9712 15086 -9678
rect 15120 -9712 15160 -9678
rect 15194 -9712 15234 -9678
rect 15268 -9712 15308 -9678
rect 15342 -9712 15382 -9678
rect 15416 -9712 15456 -9678
rect 15490 -9712 15530 -9678
rect 15564 -9712 15604 -9678
rect 15638 -9712 15678 -9678
rect 15712 -9712 15752 -9678
rect 15786 -9712 15826 -9678
rect 15860 -9712 15900 -9678
rect 15934 -9712 15974 -9678
rect 16008 -9712 16048 -9678
rect 16082 -9712 16122 -9678
rect 16156 -9712 16196 -9678
rect 16230 -9712 16270 -9678
rect 16304 -9712 16344 -9678
rect 16378 -9712 16418 -9678
rect 16452 -9712 16492 -9678
rect 16526 -9712 16566 -9678
rect 16600 -9712 16640 -9678
rect 16674 -9712 16714 -9678
rect 16748 -9712 16788 -9678
rect 16822 -9712 16862 -9678
rect 16896 -9712 16936 -9678
rect 16970 -9712 17010 -9678
rect 17044 -9712 17084 -9678
rect 17118 -9712 17158 -9678
rect 17192 -9712 17232 -9678
rect 17266 -9712 17306 -9678
rect 17340 -9712 17380 -9678
rect 17414 -9712 17454 -9678
rect 17488 -9712 17528 -9678
rect 17562 -9712 17602 -9678
rect 17636 -9712 17676 -9678
rect 17710 -9712 17750 -9678
rect 17784 -9712 17824 -9678
rect 17858 -9712 17898 -9678
rect 17932 -9712 17972 -9678
rect 18006 -9712 18046 -9678
rect 18080 -9712 18120 -9678
rect 18154 -9712 18194 -9678
rect 18228 -9712 18268 -9678
rect 18302 -9712 18342 -9678
rect 18376 -9712 18416 -9678
rect 18450 -9712 18490 -9678
rect 18524 -9712 18564 -9678
rect 18598 -9712 18638 -9678
rect 18672 -9712 18712 -9678
rect 18746 -9712 18786 -9678
rect 18820 -9712 18860 -9678
rect 18894 -9712 18934 -9678
rect 18968 -9712 19008 -9678
rect 19042 -9712 19082 -9678
rect 19116 -9712 19156 -9678
rect 19190 -9712 19230 -9678
rect 19264 -9712 19304 -9678
rect 19338 -9712 19378 -9678
rect 19412 -9712 19452 -9678
rect 19486 -9712 19526 -9678
rect 19560 -9712 19600 -9678
rect 19634 -9712 19674 -9678
rect 19708 -9712 19748 -9678
rect 19782 -9712 19822 -9678
rect 19856 -9712 19896 -9678
rect 19930 -9712 19970 -9678
rect 20004 -9712 20044 -9678
rect 20078 -9712 20118 -9678
rect 20152 -9712 20192 -9678
rect 20226 -9712 20266 -9678
rect 20300 -9712 20340 -9678
rect 20374 -9712 20414 -9678
rect 20448 -9712 20488 -9678
rect 20522 -9712 20562 -9678
rect 20596 -9712 20636 -9678
rect 20670 -9712 20710 -9678
rect 20744 -9712 20784 -9678
rect 20818 -9712 20858 -9678
rect 20892 -9712 20932 -9678
rect 20966 -9712 21006 -9678
rect 21040 -9712 21080 -9678
rect 21114 -9712 21154 -9678
rect 21188 -9712 21228 -9678
rect 21262 -9712 21302 -9678
rect 21336 -9712 21376 -9678
rect 21410 -9712 21450 -9678
rect 21484 -9712 21524 -9678
rect 21558 -9712 21598 -9678
rect 21632 -9712 21672 -9678
rect 21706 -9712 21746 -9678
rect 21780 -9712 21820 -9678
rect 21854 -9712 21894 -9678
rect 21928 -9712 21968 -9678
rect 22002 -9712 22042 -9678
rect 22076 -9712 22116 -9678
rect 22150 -9712 22190 -9678
rect 22224 -9712 22264 -9678
rect 22298 -9712 22338 -9678
rect 22372 -9712 22412 -9678
rect 22446 -9712 22486 -9678
rect 22520 -9712 22560 -9678
rect 22594 -9712 22634 -9678
rect 22668 -9712 22708 -9678
rect 22742 -9712 22782 -9678
rect 22816 -9712 22856 -9678
rect 22890 -9712 22930 -9678
rect 22964 -9712 23004 -9678
rect 23038 -9712 23078 -9678
rect 23112 -9712 23152 -9678
rect 23186 -9712 23226 -9678
rect 23260 -9712 23300 -9678
rect 23334 -9712 23374 -9678
rect 23408 -9712 23448 -9678
rect 23482 -9712 23522 -9678
rect 23556 -9712 23596 -9678
rect 23630 -9712 23670 -9678
rect 23704 -9712 23744 -9678
rect 23778 -9712 23818 -9678
rect 23852 -9712 23892 -9678
rect 23926 -9712 23966 -9678
rect 24000 -9712 24040 -9678
rect 24074 -9712 24114 -9678
rect 24148 -9712 24188 -9678
rect 24222 -9712 24262 -9678
rect 24296 -9712 24336 -9678
rect 24370 -9712 24410 -9678
rect 24444 -9712 24484 -9678
rect 24518 -9712 24558 -9678
rect 24592 -9712 24632 -9678
rect 24666 -9712 24706 -9678
rect 24740 -9712 24780 -9678
rect 24814 -9712 24854 -9678
rect 24888 -9712 24928 -9678
rect 24962 -9712 25002 -9678
rect 25036 -9712 25076 -9678
rect 25110 -9712 25150 -9678
rect 25184 -9712 25224 -9678
rect 4019 -9752 25224 -9712
rect 4019 -9786 4060 -9752
rect 4094 -9786 4134 -9752
rect 4168 -9786 4208 -9752
rect 4242 -9786 4282 -9752
rect 4316 -9786 4356 -9752
rect 4390 -9786 4430 -9752
rect 4464 -9786 4504 -9752
rect 4538 -9786 4578 -9752
rect 4612 -9786 4652 -9752
rect 4686 -9786 4726 -9752
rect 4760 -9786 4800 -9752
rect 4834 -9786 4874 -9752
rect 4908 -9786 4948 -9752
rect 4982 -9786 5022 -9752
rect 5056 -9786 5096 -9752
rect 5130 -9786 5170 -9752
rect 5204 -9786 5244 -9752
rect 5278 -9786 5318 -9752
rect 5352 -9786 5392 -9752
rect 5426 -9786 5466 -9752
rect 5500 -9786 5540 -9752
rect 5574 -9786 5614 -9752
rect 5648 -9786 5688 -9752
rect 5722 -9786 5762 -9752
rect 5796 -9786 5836 -9752
rect 5870 -9786 5910 -9752
rect 5944 -9786 5984 -9752
rect 6018 -9786 6058 -9752
rect 6092 -9786 6132 -9752
rect 6166 -9786 6206 -9752
rect 6240 -9786 6280 -9752
rect 6314 -9786 6354 -9752
rect 6388 -9786 6428 -9752
rect 6462 -9786 6502 -9752
rect 6536 -9786 6576 -9752
rect 6610 -9786 6650 -9752
rect 6684 -9786 6724 -9752
rect 6758 -9786 6798 -9752
rect 6832 -9786 6872 -9752
rect 6906 -9786 6946 -9752
rect 6980 -9786 7020 -9752
rect 7054 -9786 7094 -9752
rect 7128 -9786 7168 -9752
rect 7202 -9786 7242 -9752
rect 7276 -9786 7316 -9752
rect 7350 -9786 7390 -9752
rect 7424 -9786 7464 -9752
rect 7498 -9786 7538 -9752
rect 7572 -9786 7612 -9752
rect 7646 -9786 7686 -9752
rect 7720 -9786 7760 -9752
rect 7794 -9786 7834 -9752
rect 7868 -9786 7908 -9752
rect 7942 -9786 7982 -9752
rect 8016 -9786 8056 -9752
rect 8090 -9786 8130 -9752
rect 8164 -9786 8204 -9752
rect 8238 -9786 8278 -9752
rect 8312 -9786 8352 -9752
rect 8386 -9786 8426 -9752
rect 8460 -9786 8500 -9752
rect 8534 -9786 8574 -9752
rect 8608 -9786 8648 -9752
rect 8682 -9786 8722 -9752
rect 8756 -9786 8796 -9752
rect 8830 -9786 8870 -9752
rect 8904 -9786 8944 -9752
rect 8978 -9786 9018 -9752
rect 9052 -9786 9092 -9752
rect 9126 -9786 9166 -9752
rect 9200 -9786 9240 -9752
rect 9274 -9786 9314 -9752
rect 9348 -9786 9388 -9752
rect 9422 -9786 9462 -9752
rect 9496 -9786 9536 -9752
rect 9570 -9786 9610 -9752
rect 9644 -9786 9684 -9752
rect 9718 -9786 9758 -9752
rect 9792 -9786 9832 -9752
rect 9866 -9786 9906 -9752
rect 9940 -9786 9980 -9752
rect 10014 -9786 10054 -9752
rect 10088 -9786 10128 -9752
rect 10162 -9786 10202 -9752
rect 10236 -9786 10276 -9752
rect 10310 -9786 10350 -9752
rect 10384 -9786 10424 -9752
rect 10458 -9786 10498 -9752
rect 10532 -9786 10572 -9752
rect 10606 -9786 10646 -9752
rect 10680 -9786 10720 -9752
rect 10754 -9786 10794 -9752
rect 10828 -9786 10868 -9752
rect 10902 -9786 10942 -9752
rect 10976 -9786 11016 -9752
rect 11050 -9786 11090 -9752
rect 11124 -9786 11164 -9752
rect 11198 -9786 11238 -9752
rect 11272 -9786 11312 -9752
rect 11346 -9786 11386 -9752
rect 11420 -9786 11460 -9752
rect 11494 -9786 11534 -9752
rect 11568 -9786 11608 -9752
rect 11642 -9786 11682 -9752
rect 11716 -9786 11756 -9752
rect 11790 -9786 11830 -9752
rect 11864 -9786 11904 -9752
rect 11938 -9786 11978 -9752
rect 12012 -9786 12052 -9752
rect 12086 -9786 12126 -9752
rect 12160 -9786 12200 -9752
rect 12234 -9786 12274 -9752
rect 12308 -9786 12348 -9752
rect 12382 -9786 12422 -9752
rect 12456 -9786 12496 -9752
rect 12530 -9786 12570 -9752
rect 12604 -9786 12644 -9752
rect 12678 -9786 12718 -9752
rect 12752 -9786 12792 -9752
rect 12826 -9786 12866 -9752
rect 12900 -9786 12940 -9752
rect 12974 -9786 13014 -9752
rect 13048 -9786 13088 -9752
rect 13122 -9786 13162 -9752
rect 13196 -9786 13236 -9752
rect 13270 -9786 13310 -9752
rect 13344 -9786 13384 -9752
rect 13418 -9786 13458 -9752
rect 13492 -9786 13532 -9752
rect 13566 -9786 13606 -9752
rect 13640 -9786 13680 -9752
rect 13714 -9786 13754 -9752
rect 13788 -9786 13828 -9752
rect 13862 -9786 13902 -9752
rect 13936 -9786 13976 -9752
rect 14010 -9786 14050 -9752
rect 14084 -9786 14124 -9752
rect 14158 -9786 14198 -9752
rect 14232 -9786 14272 -9752
rect 14306 -9786 14346 -9752
rect 14380 -9786 14420 -9752
rect 14454 -9786 14494 -9752
rect 14528 -9786 14568 -9752
rect 14602 -9786 14642 -9752
rect 14676 -9786 14716 -9752
rect 14750 -9786 14790 -9752
rect 14824 -9786 14864 -9752
rect 14898 -9786 14938 -9752
rect 14972 -9786 15012 -9752
rect 15046 -9786 15086 -9752
rect 15120 -9786 15160 -9752
rect 15194 -9786 15234 -9752
rect 15268 -9786 15308 -9752
rect 15342 -9786 15382 -9752
rect 15416 -9786 15456 -9752
rect 15490 -9786 15530 -9752
rect 15564 -9786 15604 -9752
rect 15638 -9786 15678 -9752
rect 15712 -9786 15752 -9752
rect 15786 -9786 15826 -9752
rect 15860 -9786 15900 -9752
rect 15934 -9786 15974 -9752
rect 16008 -9786 16048 -9752
rect 16082 -9786 16122 -9752
rect 16156 -9786 16196 -9752
rect 16230 -9786 16270 -9752
rect 16304 -9786 16344 -9752
rect 16378 -9786 16418 -9752
rect 16452 -9786 16492 -9752
rect 16526 -9786 16566 -9752
rect 16600 -9786 16640 -9752
rect 16674 -9786 16714 -9752
rect 16748 -9786 16788 -9752
rect 16822 -9786 16862 -9752
rect 16896 -9786 16936 -9752
rect 16970 -9786 17010 -9752
rect 17044 -9786 17084 -9752
rect 17118 -9786 17158 -9752
rect 17192 -9786 17232 -9752
rect 17266 -9786 17306 -9752
rect 17340 -9786 17380 -9752
rect 17414 -9786 17454 -9752
rect 17488 -9786 17528 -9752
rect 17562 -9786 17602 -9752
rect 17636 -9786 17676 -9752
rect 17710 -9786 17750 -9752
rect 17784 -9786 17824 -9752
rect 17858 -9786 17898 -9752
rect 17932 -9786 17972 -9752
rect 18006 -9786 18046 -9752
rect 18080 -9786 18120 -9752
rect 18154 -9786 18194 -9752
rect 18228 -9786 18268 -9752
rect 18302 -9786 18342 -9752
rect 18376 -9786 18416 -9752
rect 18450 -9786 18490 -9752
rect 18524 -9786 18564 -9752
rect 18598 -9786 18638 -9752
rect 18672 -9786 18712 -9752
rect 18746 -9786 18786 -9752
rect 18820 -9786 18860 -9752
rect 18894 -9786 18934 -9752
rect 18968 -9786 19008 -9752
rect 19042 -9786 19082 -9752
rect 19116 -9786 19156 -9752
rect 19190 -9786 19230 -9752
rect 19264 -9786 19304 -9752
rect 19338 -9786 19378 -9752
rect 19412 -9786 19452 -9752
rect 19486 -9786 19526 -9752
rect 19560 -9786 19600 -9752
rect 19634 -9786 19674 -9752
rect 19708 -9786 19748 -9752
rect 19782 -9786 19822 -9752
rect 19856 -9786 19896 -9752
rect 19930 -9786 19970 -9752
rect 20004 -9786 20044 -9752
rect 20078 -9786 20118 -9752
rect 20152 -9786 20192 -9752
rect 20226 -9786 20266 -9752
rect 20300 -9786 20340 -9752
rect 20374 -9786 20414 -9752
rect 20448 -9786 20488 -9752
rect 20522 -9786 20562 -9752
rect 20596 -9786 20636 -9752
rect 20670 -9786 20710 -9752
rect 20744 -9786 20784 -9752
rect 20818 -9786 20858 -9752
rect 20892 -9786 20932 -9752
rect 20966 -9786 21006 -9752
rect 21040 -9786 21080 -9752
rect 21114 -9786 21154 -9752
rect 21188 -9786 21228 -9752
rect 21262 -9786 21302 -9752
rect 21336 -9786 21376 -9752
rect 21410 -9786 21450 -9752
rect 21484 -9786 21524 -9752
rect 21558 -9786 21598 -9752
rect 21632 -9786 21672 -9752
rect 21706 -9786 21746 -9752
rect 21780 -9786 21820 -9752
rect 21854 -9786 21894 -9752
rect 21928 -9786 21968 -9752
rect 22002 -9786 22042 -9752
rect 22076 -9786 22116 -9752
rect 22150 -9786 22190 -9752
rect 22224 -9786 22264 -9752
rect 22298 -9786 22338 -9752
rect 22372 -9786 22412 -9752
rect 22446 -9786 22486 -9752
rect 22520 -9786 22560 -9752
rect 22594 -9786 22634 -9752
rect 22668 -9786 22708 -9752
rect 22742 -9786 22782 -9752
rect 22816 -9786 22856 -9752
rect 22890 -9786 22930 -9752
rect 22964 -9786 23004 -9752
rect 23038 -9786 23078 -9752
rect 23112 -9786 23152 -9752
rect 23186 -9786 23226 -9752
rect 23260 -9786 23300 -9752
rect 23334 -9786 23374 -9752
rect 23408 -9786 23448 -9752
rect 23482 -9786 23522 -9752
rect 23556 -9786 23596 -9752
rect 23630 -9786 23670 -9752
rect 23704 -9786 23744 -9752
rect 23778 -9786 23818 -9752
rect 23852 -9786 23892 -9752
rect 23926 -9786 23966 -9752
rect 24000 -9786 24040 -9752
rect 24074 -9786 24114 -9752
rect 24148 -9786 24188 -9752
rect 24222 -9786 24262 -9752
rect 24296 -9786 24336 -9752
rect 24370 -9786 24410 -9752
rect 24444 -9786 24484 -9752
rect 24518 -9786 24558 -9752
rect 24592 -9786 24632 -9752
rect 24666 -9786 24706 -9752
rect 24740 -9786 24780 -9752
rect 24814 -9786 24854 -9752
rect 24888 -9786 24928 -9752
rect 24962 -9786 25002 -9752
rect 25036 -9786 25076 -9752
rect 25110 -9786 25150 -9752
rect 25184 -9786 25224 -9752
rect 4019 -9826 25224 -9786
rect 4019 -9860 4060 -9826
rect 4094 -9860 4134 -9826
rect 4168 -9860 4208 -9826
rect 4242 -9860 4282 -9826
rect 4316 -9860 4356 -9826
rect 4390 -9860 4430 -9826
rect 4464 -9860 4504 -9826
rect 4538 -9860 4578 -9826
rect 4612 -9860 4652 -9826
rect 4686 -9860 4726 -9826
rect 4760 -9860 4800 -9826
rect 4834 -9860 4874 -9826
rect 4908 -9860 4948 -9826
rect 4982 -9860 5022 -9826
rect 5056 -9860 5096 -9826
rect 5130 -9860 5170 -9826
rect 5204 -9860 5244 -9826
rect 5278 -9860 5318 -9826
rect 5352 -9860 5392 -9826
rect 5426 -9860 5466 -9826
rect 5500 -9860 5540 -9826
rect 5574 -9860 5614 -9826
rect 5648 -9860 5688 -9826
rect 5722 -9860 5762 -9826
rect 5796 -9860 5836 -9826
rect 5870 -9860 5910 -9826
rect 5944 -9860 5984 -9826
rect 6018 -9860 6058 -9826
rect 6092 -9860 6132 -9826
rect 6166 -9860 6206 -9826
rect 6240 -9860 6280 -9826
rect 6314 -9860 6354 -9826
rect 6388 -9860 6428 -9826
rect 6462 -9860 6502 -9826
rect 6536 -9860 6576 -9826
rect 6610 -9860 6650 -9826
rect 6684 -9860 6724 -9826
rect 6758 -9860 6798 -9826
rect 6832 -9860 6872 -9826
rect 6906 -9860 6946 -9826
rect 6980 -9860 7020 -9826
rect 7054 -9860 7094 -9826
rect 7128 -9860 7168 -9826
rect 7202 -9860 7242 -9826
rect 7276 -9860 7316 -9826
rect 7350 -9860 7390 -9826
rect 7424 -9860 7464 -9826
rect 7498 -9860 7538 -9826
rect 7572 -9860 7612 -9826
rect 7646 -9860 7686 -9826
rect 7720 -9860 7760 -9826
rect 7794 -9860 7834 -9826
rect 7868 -9860 7908 -9826
rect 7942 -9860 7982 -9826
rect 8016 -9860 8056 -9826
rect 8090 -9860 8130 -9826
rect 8164 -9860 8204 -9826
rect 8238 -9860 8278 -9826
rect 8312 -9860 8352 -9826
rect 8386 -9860 8426 -9826
rect 8460 -9860 8500 -9826
rect 8534 -9860 8574 -9826
rect 8608 -9860 8648 -9826
rect 8682 -9860 8722 -9826
rect 8756 -9860 8796 -9826
rect 8830 -9860 8870 -9826
rect 8904 -9860 8944 -9826
rect 8978 -9860 9018 -9826
rect 9052 -9860 9092 -9826
rect 9126 -9860 9166 -9826
rect 9200 -9860 9240 -9826
rect 9274 -9860 9314 -9826
rect 9348 -9860 9388 -9826
rect 9422 -9860 9462 -9826
rect 9496 -9860 9536 -9826
rect 9570 -9860 9610 -9826
rect 9644 -9860 9684 -9826
rect 9718 -9860 9758 -9826
rect 9792 -9860 9832 -9826
rect 9866 -9860 9906 -9826
rect 9940 -9860 9980 -9826
rect 10014 -9860 10054 -9826
rect 10088 -9860 10128 -9826
rect 10162 -9860 10202 -9826
rect 10236 -9860 10276 -9826
rect 10310 -9860 10350 -9826
rect 10384 -9860 10424 -9826
rect 10458 -9860 10498 -9826
rect 10532 -9860 10572 -9826
rect 10606 -9860 10646 -9826
rect 10680 -9860 10720 -9826
rect 10754 -9860 10794 -9826
rect 10828 -9860 10868 -9826
rect 10902 -9860 10942 -9826
rect 10976 -9860 11016 -9826
rect 11050 -9860 11090 -9826
rect 11124 -9860 11164 -9826
rect 11198 -9860 11238 -9826
rect 11272 -9860 11312 -9826
rect 11346 -9860 11386 -9826
rect 11420 -9860 11460 -9826
rect 11494 -9860 11534 -9826
rect 11568 -9860 11608 -9826
rect 11642 -9860 11682 -9826
rect 11716 -9860 11756 -9826
rect 11790 -9860 11830 -9826
rect 11864 -9860 11904 -9826
rect 11938 -9860 11978 -9826
rect 12012 -9860 12052 -9826
rect 12086 -9860 12126 -9826
rect 12160 -9860 12200 -9826
rect 12234 -9860 12274 -9826
rect 12308 -9860 12348 -9826
rect 12382 -9860 12422 -9826
rect 12456 -9860 12496 -9826
rect 12530 -9860 12570 -9826
rect 12604 -9860 12644 -9826
rect 12678 -9860 12718 -9826
rect 12752 -9860 12792 -9826
rect 12826 -9860 12866 -9826
rect 12900 -9860 12940 -9826
rect 12974 -9860 13014 -9826
rect 13048 -9860 13088 -9826
rect 13122 -9860 13162 -9826
rect 13196 -9860 13236 -9826
rect 13270 -9860 13310 -9826
rect 13344 -9860 13384 -9826
rect 13418 -9860 13458 -9826
rect 13492 -9860 13532 -9826
rect 13566 -9860 13606 -9826
rect 13640 -9860 13680 -9826
rect 13714 -9860 13754 -9826
rect 13788 -9860 13828 -9826
rect 13862 -9860 13902 -9826
rect 13936 -9860 13976 -9826
rect 14010 -9860 14050 -9826
rect 14084 -9860 14124 -9826
rect 14158 -9860 14198 -9826
rect 14232 -9860 14272 -9826
rect 14306 -9860 14346 -9826
rect 14380 -9860 14420 -9826
rect 14454 -9860 14494 -9826
rect 14528 -9860 14568 -9826
rect 14602 -9860 14642 -9826
rect 14676 -9860 14716 -9826
rect 14750 -9860 14790 -9826
rect 14824 -9860 14864 -9826
rect 14898 -9860 14938 -9826
rect 14972 -9860 15012 -9826
rect 15046 -9860 15086 -9826
rect 15120 -9860 15160 -9826
rect 15194 -9860 15234 -9826
rect 15268 -9860 15308 -9826
rect 15342 -9860 15382 -9826
rect 15416 -9860 15456 -9826
rect 15490 -9860 15530 -9826
rect 15564 -9860 15604 -9826
rect 15638 -9860 15678 -9826
rect 15712 -9860 15752 -9826
rect 15786 -9860 15826 -9826
rect 15860 -9860 15900 -9826
rect 15934 -9860 15974 -9826
rect 16008 -9860 16048 -9826
rect 16082 -9860 16122 -9826
rect 16156 -9860 16196 -9826
rect 16230 -9860 16270 -9826
rect 16304 -9860 16344 -9826
rect 16378 -9860 16418 -9826
rect 16452 -9860 16492 -9826
rect 16526 -9860 16566 -9826
rect 16600 -9860 16640 -9826
rect 16674 -9860 16714 -9826
rect 16748 -9860 16788 -9826
rect 16822 -9860 16862 -9826
rect 16896 -9860 16936 -9826
rect 16970 -9860 17010 -9826
rect 17044 -9860 17084 -9826
rect 17118 -9860 17158 -9826
rect 17192 -9860 17232 -9826
rect 17266 -9860 17306 -9826
rect 17340 -9860 17380 -9826
rect 17414 -9860 17454 -9826
rect 17488 -9860 17528 -9826
rect 17562 -9860 17602 -9826
rect 17636 -9860 17676 -9826
rect 17710 -9860 17750 -9826
rect 17784 -9860 17824 -9826
rect 17858 -9860 17898 -9826
rect 17932 -9860 17972 -9826
rect 18006 -9860 18046 -9826
rect 18080 -9860 18120 -9826
rect 18154 -9860 18194 -9826
rect 18228 -9860 18268 -9826
rect 18302 -9860 18342 -9826
rect 18376 -9860 18416 -9826
rect 18450 -9860 18490 -9826
rect 18524 -9860 18564 -9826
rect 18598 -9860 18638 -9826
rect 18672 -9860 18712 -9826
rect 18746 -9860 18786 -9826
rect 18820 -9860 18860 -9826
rect 18894 -9860 18934 -9826
rect 18968 -9860 19008 -9826
rect 19042 -9860 19082 -9826
rect 19116 -9860 19156 -9826
rect 19190 -9860 19230 -9826
rect 19264 -9860 19304 -9826
rect 19338 -9860 19378 -9826
rect 19412 -9860 19452 -9826
rect 19486 -9860 19526 -9826
rect 19560 -9860 19600 -9826
rect 19634 -9860 19674 -9826
rect 19708 -9860 19748 -9826
rect 19782 -9860 19822 -9826
rect 19856 -9860 19896 -9826
rect 19930 -9860 19970 -9826
rect 20004 -9860 20044 -9826
rect 20078 -9860 20118 -9826
rect 20152 -9860 20192 -9826
rect 20226 -9860 20266 -9826
rect 20300 -9860 20340 -9826
rect 20374 -9860 20414 -9826
rect 20448 -9860 20488 -9826
rect 20522 -9860 20562 -9826
rect 20596 -9860 20636 -9826
rect 20670 -9860 20710 -9826
rect 20744 -9860 20784 -9826
rect 20818 -9860 20858 -9826
rect 20892 -9860 20932 -9826
rect 20966 -9860 21006 -9826
rect 21040 -9860 21080 -9826
rect 21114 -9860 21154 -9826
rect 21188 -9860 21228 -9826
rect 21262 -9860 21302 -9826
rect 21336 -9860 21376 -9826
rect 21410 -9860 21450 -9826
rect 21484 -9860 21524 -9826
rect 21558 -9860 21598 -9826
rect 21632 -9860 21672 -9826
rect 21706 -9860 21746 -9826
rect 21780 -9860 21820 -9826
rect 21854 -9860 21894 -9826
rect 21928 -9860 21968 -9826
rect 22002 -9860 22042 -9826
rect 22076 -9860 22116 -9826
rect 22150 -9860 22190 -9826
rect 22224 -9860 22264 -9826
rect 22298 -9860 22338 -9826
rect 22372 -9860 22412 -9826
rect 22446 -9860 22486 -9826
rect 22520 -9860 22560 -9826
rect 22594 -9860 22634 -9826
rect 22668 -9860 22708 -9826
rect 22742 -9860 22782 -9826
rect 22816 -9860 22856 -9826
rect 22890 -9860 22930 -9826
rect 22964 -9860 23004 -9826
rect 23038 -9860 23078 -9826
rect 23112 -9860 23152 -9826
rect 23186 -9860 23226 -9826
rect 23260 -9860 23300 -9826
rect 23334 -9860 23374 -9826
rect 23408 -9860 23448 -9826
rect 23482 -9860 23522 -9826
rect 23556 -9860 23596 -9826
rect 23630 -9860 23670 -9826
rect 23704 -9860 23744 -9826
rect 23778 -9860 23818 -9826
rect 23852 -9860 23892 -9826
rect 23926 -9860 23966 -9826
rect 24000 -9860 24040 -9826
rect 24074 -9860 24114 -9826
rect 24148 -9860 24188 -9826
rect 24222 -9860 24262 -9826
rect 24296 -9860 24336 -9826
rect 24370 -9860 24410 -9826
rect 24444 -9860 24484 -9826
rect 24518 -9860 24558 -9826
rect 24592 -9860 24632 -9826
rect 24666 -9860 24706 -9826
rect 24740 -9860 24780 -9826
rect 24814 -9860 24854 -9826
rect 24888 -9860 24928 -9826
rect 24962 -9860 25002 -9826
rect 25036 -9860 25076 -9826
rect 25110 -9860 25150 -9826
rect 25184 -9860 25224 -9826
rect 4019 -9900 25224 -9860
rect 4019 -9933 4060 -9900
rect 4020 -9934 4060 -9933
rect 4094 -9934 4134 -9900
rect 4168 -9934 4208 -9900
rect 4242 -9934 4282 -9900
rect 4316 -9934 4356 -9900
rect 4390 -9934 4430 -9900
rect 4464 -9934 4504 -9900
rect 4538 -9934 4578 -9900
rect 4612 -9934 4652 -9900
rect 4686 -9934 4726 -9900
rect 4760 -9934 4800 -9900
rect 4834 -9934 4874 -9900
rect 4908 -9934 4948 -9900
rect 4982 -9934 5022 -9900
rect 5056 -9934 5096 -9900
rect 5130 -9934 5170 -9900
rect 5204 -9934 5244 -9900
rect 5278 -9934 5318 -9900
rect 5352 -9934 5392 -9900
rect 5426 -9934 5466 -9900
rect 5500 -9934 5540 -9900
rect 5574 -9934 5614 -9900
rect 5648 -9934 5688 -9900
rect 5722 -9934 5762 -9900
rect 5796 -9934 5836 -9900
rect 5870 -9934 5910 -9900
rect 5944 -9934 5984 -9900
rect 6018 -9934 6058 -9900
rect 6092 -9934 6132 -9900
rect 6166 -9934 6206 -9900
rect 6240 -9934 6280 -9900
rect 6314 -9934 6354 -9900
rect 6388 -9934 6428 -9900
rect 6462 -9934 6502 -9900
rect 6536 -9934 6576 -9900
rect 6610 -9934 6650 -9900
rect 6684 -9934 6724 -9900
rect 6758 -9934 6798 -9900
rect 6832 -9934 6872 -9900
rect 6906 -9934 6946 -9900
rect 6980 -9934 7020 -9900
rect 7054 -9934 7094 -9900
rect 7128 -9934 7168 -9900
rect 7202 -9934 7242 -9900
rect 7276 -9934 7316 -9900
rect 7350 -9934 7390 -9900
rect 7424 -9934 7464 -9900
rect 7498 -9934 7538 -9900
rect 7572 -9934 7612 -9900
rect 7646 -9934 7686 -9900
rect 7720 -9934 7760 -9900
rect 7794 -9934 7834 -9900
rect 7868 -9934 7908 -9900
rect 7942 -9934 7982 -9900
rect 8016 -9934 8056 -9900
rect 8090 -9934 8130 -9900
rect 8164 -9934 8204 -9900
rect 8238 -9934 8278 -9900
rect 8312 -9934 8352 -9900
rect 8386 -9934 8426 -9900
rect 8460 -9934 8500 -9900
rect 8534 -9934 8574 -9900
rect 8608 -9934 8648 -9900
rect 8682 -9934 8722 -9900
rect 8756 -9934 8796 -9900
rect 8830 -9934 8870 -9900
rect 8904 -9934 8944 -9900
rect 8978 -9934 9018 -9900
rect 9052 -9934 9092 -9900
rect 9126 -9934 9166 -9900
rect 9200 -9934 9240 -9900
rect 9274 -9934 9314 -9900
rect 9348 -9934 9388 -9900
rect 9422 -9934 9462 -9900
rect 9496 -9934 9536 -9900
rect 9570 -9934 9610 -9900
rect 9644 -9934 9684 -9900
rect 9718 -9934 9758 -9900
rect 9792 -9934 9832 -9900
rect 9866 -9934 9906 -9900
rect 9940 -9934 9980 -9900
rect 10014 -9934 10054 -9900
rect 10088 -9934 10128 -9900
rect 10162 -9934 10202 -9900
rect 10236 -9934 10276 -9900
rect 10310 -9934 10350 -9900
rect 10384 -9934 10424 -9900
rect 10458 -9934 10498 -9900
rect 10532 -9934 10572 -9900
rect 10606 -9934 10646 -9900
rect 10680 -9934 10720 -9900
rect 10754 -9934 10794 -9900
rect 10828 -9934 10868 -9900
rect 10902 -9934 10942 -9900
rect 10976 -9934 11016 -9900
rect 11050 -9934 11090 -9900
rect 11124 -9934 11164 -9900
rect 11198 -9934 11238 -9900
rect 11272 -9934 11312 -9900
rect 11346 -9934 11386 -9900
rect 11420 -9934 11460 -9900
rect 11494 -9934 11534 -9900
rect 11568 -9934 11608 -9900
rect 11642 -9934 11682 -9900
rect 11716 -9934 11756 -9900
rect 11790 -9934 11830 -9900
rect 11864 -9934 11904 -9900
rect 11938 -9934 11978 -9900
rect 12012 -9934 12052 -9900
rect 12086 -9934 12126 -9900
rect 12160 -9934 12200 -9900
rect 12234 -9934 12274 -9900
rect 12308 -9934 12348 -9900
rect 12382 -9934 12422 -9900
rect 12456 -9934 12496 -9900
rect 12530 -9934 12570 -9900
rect 12604 -9934 12644 -9900
rect 12678 -9934 12718 -9900
rect 12752 -9934 12792 -9900
rect 12826 -9934 12866 -9900
rect 12900 -9934 12940 -9900
rect 12974 -9934 13014 -9900
rect 13048 -9934 13088 -9900
rect 13122 -9934 13162 -9900
rect 13196 -9934 13236 -9900
rect 13270 -9934 13310 -9900
rect 13344 -9934 13384 -9900
rect 13418 -9934 13458 -9900
rect 13492 -9934 13532 -9900
rect 13566 -9934 13606 -9900
rect 13640 -9934 13680 -9900
rect 13714 -9934 13754 -9900
rect 13788 -9934 13828 -9900
rect 13862 -9934 13902 -9900
rect 13936 -9934 13976 -9900
rect 14010 -9934 14050 -9900
rect 14084 -9934 14124 -9900
rect 14158 -9934 14198 -9900
rect 14232 -9934 14272 -9900
rect 14306 -9934 14346 -9900
rect 14380 -9934 14420 -9900
rect 14454 -9934 14494 -9900
rect 14528 -9934 14568 -9900
rect 14602 -9934 14642 -9900
rect 14676 -9934 14716 -9900
rect 14750 -9934 14790 -9900
rect 14824 -9934 14864 -9900
rect 14898 -9934 14938 -9900
rect 14972 -9934 15012 -9900
rect 15046 -9934 15086 -9900
rect 15120 -9934 15160 -9900
rect 15194 -9934 15234 -9900
rect 15268 -9934 15308 -9900
rect 15342 -9934 15382 -9900
rect 15416 -9934 15456 -9900
rect 15490 -9934 15530 -9900
rect 15564 -9934 15604 -9900
rect 15638 -9934 15678 -9900
rect 15712 -9934 15752 -9900
rect 15786 -9934 15826 -9900
rect 15860 -9934 15900 -9900
rect 15934 -9934 15974 -9900
rect 16008 -9934 16048 -9900
rect 16082 -9934 16122 -9900
rect 16156 -9934 16196 -9900
rect 16230 -9934 16270 -9900
rect 16304 -9934 16344 -9900
rect 16378 -9934 16418 -9900
rect 16452 -9934 16492 -9900
rect 16526 -9934 16566 -9900
rect 16600 -9934 16640 -9900
rect 16674 -9934 16714 -9900
rect 16748 -9934 16788 -9900
rect 16822 -9934 16862 -9900
rect 16896 -9934 16936 -9900
rect 16970 -9934 17010 -9900
rect 17044 -9934 17084 -9900
rect 17118 -9934 17158 -9900
rect 17192 -9934 17232 -9900
rect 17266 -9934 17306 -9900
rect 17340 -9934 17380 -9900
rect 17414 -9934 17454 -9900
rect 17488 -9934 17528 -9900
rect 17562 -9934 17602 -9900
rect 17636 -9934 17676 -9900
rect 17710 -9934 17750 -9900
rect 17784 -9934 17824 -9900
rect 17858 -9934 17898 -9900
rect 17932 -9934 17972 -9900
rect 18006 -9934 18046 -9900
rect 18080 -9934 18120 -9900
rect 18154 -9934 18194 -9900
rect 18228 -9934 18268 -9900
rect 18302 -9934 18342 -9900
rect 18376 -9934 18416 -9900
rect 18450 -9934 18490 -9900
rect 18524 -9934 18564 -9900
rect 18598 -9934 18638 -9900
rect 18672 -9934 18712 -9900
rect 18746 -9934 18786 -9900
rect 18820 -9934 18860 -9900
rect 18894 -9934 18934 -9900
rect 18968 -9934 19008 -9900
rect 19042 -9934 19082 -9900
rect 19116 -9934 19156 -9900
rect 19190 -9934 19230 -9900
rect 19264 -9934 19304 -9900
rect 19338 -9934 19378 -9900
rect 19412 -9934 19452 -9900
rect 19486 -9934 19526 -9900
rect 19560 -9934 19600 -9900
rect 19634 -9934 19674 -9900
rect 19708 -9934 19748 -9900
rect 19782 -9934 19822 -9900
rect 19856 -9934 19896 -9900
rect 19930 -9934 19970 -9900
rect 20004 -9934 20044 -9900
rect 20078 -9934 20118 -9900
rect 20152 -9934 20192 -9900
rect 20226 -9934 20266 -9900
rect 20300 -9934 20340 -9900
rect 20374 -9934 20414 -9900
rect 20448 -9934 20488 -9900
rect 20522 -9934 20562 -9900
rect 20596 -9934 20636 -9900
rect 20670 -9934 20710 -9900
rect 20744 -9934 20784 -9900
rect 20818 -9934 20858 -9900
rect 20892 -9934 20932 -9900
rect 20966 -9934 21006 -9900
rect 21040 -9934 21080 -9900
rect 21114 -9934 21154 -9900
rect 21188 -9934 21228 -9900
rect 21262 -9934 21302 -9900
rect 21336 -9934 21376 -9900
rect 21410 -9934 21450 -9900
rect 21484 -9934 21524 -9900
rect 21558 -9934 21598 -9900
rect 21632 -9934 21672 -9900
rect 21706 -9934 21746 -9900
rect 21780 -9934 21820 -9900
rect 21854 -9934 21894 -9900
rect 21928 -9934 21968 -9900
rect 22002 -9934 22042 -9900
rect 22076 -9934 22116 -9900
rect 22150 -9934 22190 -9900
rect 22224 -9934 22264 -9900
rect 22298 -9934 22338 -9900
rect 22372 -9934 22412 -9900
rect 22446 -9934 22486 -9900
rect 22520 -9934 22560 -9900
rect 22594 -9934 22634 -9900
rect 22668 -9934 22708 -9900
rect 22742 -9934 22782 -9900
rect 22816 -9934 22856 -9900
rect 22890 -9934 22930 -9900
rect 22964 -9934 23004 -9900
rect 23038 -9934 23078 -9900
rect 23112 -9934 23152 -9900
rect 23186 -9934 23226 -9900
rect 23260 -9934 23300 -9900
rect 23334 -9934 23374 -9900
rect 23408 -9934 23448 -9900
rect 23482 -9934 23522 -9900
rect 23556 -9934 23596 -9900
rect 23630 -9934 23670 -9900
rect 23704 -9934 23744 -9900
rect 23778 -9934 23818 -9900
rect 23852 -9934 23892 -9900
rect 23926 -9934 23966 -9900
rect 24000 -9934 24040 -9900
rect 24074 -9934 24114 -9900
rect 24148 -9934 24188 -9900
rect 24222 -9934 24262 -9900
rect 24296 -9934 24336 -9900
rect 24370 -9934 24410 -9900
rect 24444 -9934 24484 -9900
rect 24518 -9934 24558 -9900
rect 24592 -9934 24632 -9900
rect 24666 -9934 24706 -9900
rect 24740 -9934 24780 -9900
rect 24814 -9934 24854 -9900
rect 24888 -9934 24928 -9900
rect 24962 -9934 25002 -9900
rect 25036 -9934 25076 -9900
rect 25110 -9934 25150 -9900
rect 25184 -9934 25224 -9900
<< nsubdiff >>
rect 4730 3118 4792 3152
rect 10762 3118 10824 3152
rect 12420 3117 12482 3151
rect 18452 3117 18621 3151
rect 24591 3117 24653 3151
rect 4768 3030 4792 3064
rect 10762 3030 10786 3064
rect 12458 3029 12482 3063
rect 18452 3029 18476 3063
rect 18597 3029 18621 3063
rect 24591 3029 24615 3063
rect 4768 2942 4792 2976
rect 10762 2942 10786 2976
rect 12458 2941 12482 2975
rect 18452 2941 18621 2975
rect 24591 2941 24615 2975
rect 4768 1427 4792 1461
rect 10762 1427 10786 1461
rect 4696 1339 4792 1373
rect 10762 1339 10858 1373
rect 4696 1277 4730 1339
rect 10824 1277 10858 1339
rect 4696 -395 4730 -333
rect 10824 -395 10858 -333
rect 4696 -429 4792 -395
rect 10762 -429 10858 -395
rect 4768 -517 4792 -483
rect 10762 -517 10786 -483
rect 4768 -605 4792 -571
rect 10762 -605 10786 -571
rect 4696 -711 4792 -677
rect 10762 -711 10858 -677
rect 4696 -773 4730 -711
rect 10824 -773 10858 -711
rect 4696 -2445 4730 -2383
rect 10824 -2445 10858 -2383
rect 4696 -2479 4792 -2445
rect 10762 -2479 10858 -2445
rect 4768 -2567 4792 -2533
rect 10762 -2567 10786 -2533
rect 4768 -2655 4792 -2621
rect 10762 -2655 10786 -2621
rect 4696 -2761 4792 -2727
rect 10762 -2761 10858 -2727
rect 4696 -2823 4730 -2761
rect 10824 -2823 10858 -2761
rect 4696 -4495 4730 -4433
rect 10824 -4495 10858 -4433
rect 4696 -4529 4792 -4495
rect 10762 -4529 10858 -4495
rect 4768 -4617 4792 -4583
rect 10762 -4617 10786 -4583
rect 4768 -4705 4792 -4671
rect 10762 -4705 10786 -4671
rect 4768 -6667 4792 -6633
rect 10762 -6667 10786 -6633
rect 4768 -6755 4792 -6721
rect 10762 -6755 10786 -6721
<< psubdiffcont >>
rect 10737 -7593 10771 -7287
rect 11053 -7593 11087 -7287
rect 11369 -7593 11403 -7287
rect 11685 -7593 11719 -7287
rect 12001 -7593 12035 -7287
rect 12317 -7593 12351 -7287
rect 4080 -8905 4114 -8871
rect 4152 -8905 4186 -8871
rect 4234 -8905 4268 -8871
rect 4306 -8905 4340 -8871
rect 4388 -8905 4422 -8871
rect 4460 -8905 4494 -8871
rect 4542 -8905 4576 -8871
rect 4614 -8905 4648 -8871
rect 4696 -8905 4730 -8871
rect 4768 -8905 4802 -8871
rect 4850 -8905 4884 -8871
rect 4922 -8905 4956 -8871
rect 5004 -8905 5038 -8871
rect 5076 -8905 5110 -8871
rect 5158 -8905 5192 -8871
rect 5230 -8905 5264 -8871
rect 5312 -8905 5346 -8871
rect 5384 -8905 5418 -8871
rect 5466 -8905 5500 -8871
rect 5538 -8905 5572 -8871
rect 5620 -8905 5654 -8871
rect 5692 -8905 5726 -8871
rect 4080 -8979 4114 -8945
rect 4152 -8979 4186 -8945
rect 4234 -8979 4268 -8945
rect 4306 -8979 4340 -8945
rect 4388 -8979 4422 -8945
rect 4460 -8979 4494 -8945
rect 4542 -8979 4576 -8945
rect 4614 -8979 4648 -8945
rect 4696 -8979 4730 -8945
rect 4768 -8979 4802 -8945
rect 4850 -8979 4884 -8945
rect 4922 -8979 4956 -8945
rect 5004 -8979 5038 -8945
rect 5076 -8979 5110 -8945
rect 5158 -8979 5192 -8945
rect 5230 -8979 5264 -8945
rect 5312 -8979 5346 -8945
rect 5384 -8979 5418 -8945
rect 5466 -8979 5500 -8945
rect 5538 -8979 5572 -8945
rect 5620 -8979 5654 -8945
rect 5692 -8979 5726 -8945
rect 5774 -8979 5808 -8945
rect 5846 -8979 5880 -8945
rect 5928 -8979 5962 -8945
rect 6000 -8979 6034 -8945
rect 6082 -8979 6116 -8945
rect 6154 -8979 6188 -8945
rect 6236 -8979 6270 -8945
rect 6308 -8979 6342 -8945
rect 6390 -8979 6424 -8945
rect 6462 -8979 6496 -8945
rect 6544 -8979 6578 -8945
rect 6616 -8979 6650 -8945
rect 6698 -8979 6732 -8945
rect 6770 -8979 6804 -8945
rect 6852 -8979 6886 -8945
rect 6924 -8979 6958 -8945
rect 7006 -8979 7040 -8945
rect 7078 -8979 7112 -8945
rect 7160 -8979 7194 -8945
rect 7232 -8979 7266 -8945
rect 7314 -8979 7348 -8945
rect 7386 -8979 7420 -8945
rect 7468 -8979 7502 -8945
rect 7540 -8979 7574 -8945
rect 7622 -8979 7656 -8945
rect 7694 -8979 7728 -8945
rect 7776 -8979 7810 -8945
rect 7848 -8979 7882 -8945
rect 7930 -8979 7964 -8945
rect 8002 -8979 8036 -8945
rect 8084 -8979 8118 -8945
rect 8156 -8979 8190 -8945
rect 8238 -8979 8272 -8945
rect 8310 -8979 8344 -8945
rect 8392 -8979 8426 -8945
rect 8464 -8979 8498 -8945
rect 8546 -8979 8580 -8945
rect 8618 -8979 8652 -8945
rect 8700 -8979 8734 -8945
rect 8772 -8979 8806 -8945
rect 8854 -8979 8888 -8945
rect 8926 -8979 8960 -8945
rect 9008 -8979 9042 -8945
rect 9080 -8979 9114 -8945
rect 9162 -8979 9196 -8945
rect 9234 -8979 9268 -8945
rect 9316 -8979 9350 -8945
rect 9388 -8979 9422 -8945
rect 9470 -8979 9504 -8945
rect 9542 -8979 9576 -8945
rect 9624 -8979 9658 -8945
rect 9696 -8979 9730 -8945
rect 9778 -8979 9812 -8945
rect 9850 -8979 9884 -8945
rect 9932 -8979 9966 -8945
rect 10004 -8979 10038 -8945
rect 10086 -8979 10120 -8945
rect 10158 -8979 10192 -8945
rect 10240 -8979 10274 -8945
rect 10312 -8979 10346 -8945
rect 10394 -8979 10428 -8945
rect 10466 -8979 10500 -8945
rect 10548 -8979 10582 -8945
rect 10620 -8979 10654 -8945
rect 10702 -8979 10736 -8945
rect 10774 -8979 10808 -8945
rect 10856 -8979 10890 -8945
rect 10928 -8979 10962 -8945
rect 11010 -8979 11044 -8945
rect 11082 -8979 11116 -8945
rect 11164 -8979 11198 -8945
rect 11236 -8979 11270 -8945
rect 11318 -8979 11352 -8945
rect 11390 -8979 11424 -8945
rect 11472 -8979 11506 -8945
rect 11544 -8979 11578 -8945
rect 11626 -8979 11660 -8945
rect 11698 -8979 11732 -8945
rect 11780 -8979 11814 -8945
rect 11852 -8979 11886 -8945
rect 11934 -8979 11968 -8945
rect 12006 -8979 12040 -8945
rect 4080 -9053 4114 -9019
rect 4152 -9053 4186 -9019
rect 4234 -9053 4268 -9019
rect 4306 -9053 4340 -9019
rect 4388 -9053 4422 -9019
rect 4460 -9053 4494 -9019
rect 4542 -9053 4576 -9019
rect 4614 -9053 4648 -9019
rect 4696 -9053 4730 -9019
rect 4768 -9053 4802 -9019
rect 4850 -9053 4884 -9019
rect 4922 -9053 4956 -9019
rect 5004 -9053 5038 -9019
rect 5076 -9053 5110 -9019
rect 5158 -9053 5192 -9019
rect 5230 -9053 5264 -9019
rect 5312 -9053 5346 -9019
rect 5384 -9053 5418 -9019
rect 5466 -9053 5500 -9019
rect 5538 -9053 5572 -9019
rect 5620 -9053 5654 -9019
rect 5692 -9053 5726 -9019
rect 5774 -9053 5808 -9019
rect 5846 -9053 5880 -9019
rect 5928 -9053 5962 -9019
rect 6000 -9053 6034 -9019
rect 6082 -9053 6116 -9019
rect 6154 -9053 6188 -9019
rect 6236 -9053 6270 -9019
rect 6308 -9053 6342 -9019
rect 6390 -9053 6424 -9019
rect 6462 -9053 6496 -9019
rect 6544 -9053 6578 -9019
rect 6616 -9053 6650 -9019
rect 6698 -9053 6732 -9019
rect 6770 -9053 6804 -9019
rect 6852 -9053 6886 -9019
rect 6924 -9053 6958 -9019
rect 7006 -9053 7040 -9019
rect 7078 -9053 7112 -9019
rect 7160 -9053 7194 -9019
rect 7232 -9053 7266 -9019
rect 7314 -9053 7348 -9019
rect 7386 -9053 7420 -9019
rect 7468 -9053 7502 -9019
rect 7540 -9053 7574 -9019
rect 7622 -9053 7656 -9019
rect 7694 -9053 7728 -9019
rect 7776 -9053 7810 -9019
rect 7848 -9053 7882 -9019
rect 7930 -9053 7964 -9019
rect 8002 -9053 8036 -9019
rect 8084 -9053 8118 -9019
rect 8156 -9053 8190 -9019
rect 8238 -9053 8272 -9019
rect 8310 -9053 8344 -9019
rect 8392 -9053 8426 -9019
rect 8464 -9053 8498 -9019
rect 8546 -9053 8580 -9019
rect 8618 -9053 8652 -9019
rect 8700 -9053 8734 -9019
rect 8772 -9053 8806 -9019
rect 8854 -9053 8888 -9019
rect 8926 -9053 8960 -9019
rect 9008 -9053 9042 -9019
rect 9080 -9053 9114 -9019
rect 9162 -9053 9196 -9019
rect 9234 -9053 9268 -9019
rect 9316 -9053 9350 -9019
rect 9388 -9053 9422 -9019
rect 9470 -9053 9504 -9019
rect 9542 -9053 9576 -9019
rect 9624 -9053 9658 -9019
rect 9696 -9053 9730 -9019
rect 9778 -9053 9812 -9019
rect 9850 -9053 9884 -9019
rect 9932 -9053 9966 -9019
rect 10004 -9053 10038 -9019
rect 10086 -9053 10120 -9019
rect 10158 -9053 10192 -9019
rect 10240 -9053 10274 -9019
rect 10312 -9053 10346 -9019
rect 10394 -9053 10428 -9019
rect 10466 -9053 10500 -9019
rect 10548 -9053 10582 -9019
rect 10620 -9053 10654 -9019
rect 10702 -9053 10736 -9019
rect 10774 -9053 10808 -9019
rect 10856 -9053 10890 -9019
rect 10928 -9053 10962 -9019
rect 11010 -9053 11044 -9019
rect 11082 -9053 11116 -9019
rect 11164 -9053 11198 -9019
rect 11236 -9053 11270 -9019
rect 11318 -9053 11352 -9019
rect 11390 -9053 11424 -9019
rect 11472 -9053 11506 -9019
rect 11544 -9053 11578 -9019
rect 11626 -9053 11660 -9019
rect 11698 -9053 11732 -9019
rect 11780 -9053 11814 -9019
rect 11852 -9053 11886 -9019
rect 11934 -9053 11968 -9019
rect 12006 -9053 12040 -9019
rect 4080 -9127 4114 -9093
rect 4152 -9127 4186 -9093
rect 4234 -9127 4268 -9093
rect 4306 -9127 4340 -9093
rect 4388 -9127 4422 -9093
rect 4460 -9127 4494 -9093
rect 4542 -9127 4576 -9093
rect 4614 -9127 4648 -9093
rect 4696 -9127 4730 -9093
rect 4768 -9127 4802 -9093
rect 4850 -9127 4884 -9093
rect 4922 -9127 4956 -9093
rect 5004 -9127 5038 -9093
rect 5076 -9127 5110 -9093
rect 5158 -9127 5192 -9093
rect 5230 -9127 5264 -9093
rect 5312 -9127 5346 -9093
rect 5384 -9127 5418 -9093
rect 5466 -9127 5500 -9093
rect 5538 -9127 5572 -9093
rect 5620 -9127 5654 -9093
rect 5692 -9127 5726 -9093
rect 5774 -9127 5808 -9093
rect 5846 -9127 5880 -9093
rect 5928 -9127 5962 -9093
rect 6000 -9127 6034 -9093
rect 6082 -9127 6116 -9093
rect 6154 -9127 6188 -9093
rect 6236 -9127 6270 -9093
rect 6308 -9127 6342 -9093
rect 6390 -9127 6424 -9093
rect 6462 -9127 6496 -9093
rect 6544 -9127 6578 -9093
rect 6616 -9127 6650 -9093
rect 6698 -9127 6732 -9093
rect 6770 -9127 6804 -9093
rect 6852 -9127 6886 -9093
rect 6924 -9127 6958 -9093
rect 7006 -9127 7040 -9093
rect 7078 -9127 7112 -9093
rect 7160 -9127 7194 -9093
rect 7232 -9127 7266 -9093
rect 7314 -9127 7348 -9093
rect 7386 -9127 7420 -9093
rect 7468 -9127 7502 -9093
rect 7540 -9127 7574 -9093
rect 7622 -9127 7656 -9093
rect 7694 -9127 7728 -9093
rect 7776 -9127 7810 -9093
rect 7848 -9127 7882 -9093
rect 7930 -9127 7964 -9093
rect 8002 -9127 8036 -9093
rect 8084 -9127 8118 -9093
rect 8156 -9127 8190 -9093
rect 8238 -9127 8272 -9093
rect 8310 -9127 8344 -9093
rect 8392 -9127 8426 -9093
rect 8464 -9127 8498 -9093
rect 8546 -9127 8580 -9093
rect 8618 -9127 8652 -9093
rect 8700 -9127 8734 -9093
rect 8772 -9127 8806 -9093
rect 8854 -9127 8888 -9093
rect 8926 -9127 8960 -9093
rect 9008 -9127 9042 -9093
rect 9080 -9127 9114 -9093
rect 9162 -9127 9196 -9093
rect 9234 -9127 9268 -9093
rect 9316 -9127 9350 -9093
rect 9388 -9127 9422 -9093
rect 9470 -9127 9504 -9093
rect 9542 -9127 9576 -9093
rect 9624 -9127 9658 -9093
rect 9696 -9127 9730 -9093
rect 9778 -9127 9812 -9093
rect 9850 -9127 9884 -9093
rect 9932 -9127 9966 -9093
rect 10004 -9127 10038 -9093
rect 10086 -9127 10120 -9093
rect 10158 -9127 10192 -9093
rect 10240 -9127 10274 -9093
rect 10312 -9127 10346 -9093
rect 10394 -9127 10428 -9093
rect 10466 -9127 10500 -9093
rect 10548 -9127 10582 -9093
rect 10620 -9127 10654 -9093
rect 10702 -9127 10736 -9093
rect 10774 -9127 10808 -9093
rect 10856 -9127 10890 -9093
rect 10928 -9127 10962 -9093
rect 11010 -9127 11044 -9093
rect 11082 -9127 11116 -9093
rect 11164 -9127 11198 -9093
rect 11236 -9127 11270 -9093
rect 11318 -9127 11352 -9093
rect 11390 -9127 11424 -9093
rect 11472 -9127 11506 -9093
rect 11544 -9127 11578 -9093
rect 11626 -9127 11660 -9093
rect 11698 -9127 11732 -9093
rect 11780 -9127 11814 -9093
rect 11852 -9127 11886 -9093
rect 11934 -9127 11968 -9093
rect 12006 -9127 12040 -9093
rect 4080 -9201 4114 -9167
rect 4152 -9201 4186 -9167
rect 4234 -9201 4268 -9167
rect 4306 -9201 4340 -9167
rect 4388 -9201 4422 -9167
rect 4460 -9201 4494 -9167
rect 4542 -9201 4576 -9167
rect 4614 -9201 4648 -9167
rect 4696 -9201 4730 -9167
rect 4768 -9201 4802 -9167
rect 4850 -9201 4884 -9167
rect 4922 -9201 4956 -9167
rect 5004 -9201 5038 -9167
rect 5076 -9201 5110 -9167
rect 5158 -9201 5192 -9167
rect 5230 -9201 5264 -9167
rect 5312 -9201 5346 -9167
rect 5384 -9201 5418 -9167
rect 5466 -9201 5500 -9167
rect 5538 -9201 5572 -9167
rect 5620 -9201 5654 -9167
rect 5692 -9201 5726 -9167
rect 5774 -9201 5808 -9167
rect 5846 -9201 5880 -9167
rect 5928 -9201 5962 -9167
rect 6000 -9201 6034 -9167
rect 6082 -9201 6116 -9167
rect 6154 -9201 6188 -9167
rect 6236 -9201 6270 -9167
rect 6308 -9201 6342 -9167
rect 6390 -9201 6424 -9167
rect 6462 -9201 6496 -9167
rect 6544 -9201 6578 -9167
rect 6616 -9201 6650 -9167
rect 6698 -9201 6732 -9167
rect 6770 -9201 6804 -9167
rect 6852 -9201 6886 -9167
rect 6924 -9201 6958 -9167
rect 7006 -9201 7040 -9167
rect 7078 -9201 7112 -9167
rect 7160 -9201 7194 -9167
rect 7232 -9201 7266 -9167
rect 7314 -9201 7348 -9167
rect 7386 -9201 7420 -9167
rect 7468 -9201 7502 -9167
rect 7540 -9201 7574 -9167
rect 7622 -9201 7656 -9167
rect 7694 -9201 7728 -9167
rect 7776 -9201 7810 -9167
rect 7848 -9201 7882 -9167
rect 7930 -9201 7964 -9167
rect 8002 -9201 8036 -9167
rect 8084 -9201 8118 -9167
rect 8156 -9201 8190 -9167
rect 8238 -9201 8272 -9167
rect 8310 -9201 8344 -9167
rect 8392 -9201 8426 -9167
rect 8464 -9201 8498 -9167
rect 8546 -9201 8580 -9167
rect 8618 -9201 8652 -9167
rect 8700 -9201 8734 -9167
rect 8772 -9201 8806 -9167
rect 8854 -9201 8888 -9167
rect 8926 -9201 8960 -9167
rect 9008 -9201 9042 -9167
rect 9080 -9201 9114 -9167
rect 9162 -9201 9196 -9167
rect 9234 -9201 9268 -9167
rect 9316 -9201 9350 -9167
rect 9388 -9201 9422 -9167
rect 9470 -9201 9504 -9167
rect 9542 -9201 9576 -9167
rect 9624 -9201 9658 -9167
rect 9696 -9201 9730 -9167
rect 9778 -9201 9812 -9167
rect 9850 -9201 9884 -9167
rect 9932 -9201 9966 -9167
rect 10004 -9201 10038 -9167
rect 10086 -9201 10120 -9167
rect 10158 -9201 10192 -9167
rect 10240 -9201 10274 -9167
rect 10312 -9201 10346 -9167
rect 10394 -9201 10428 -9167
rect 10466 -9201 10500 -9167
rect 10548 -9201 10582 -9167
rect 10620 -9201 10654 -9167
rect 10702 -9201 10736 -9167
rect 10774 -9201 10808 -9167
rect 10856 -9201 10890 -9167
rect 10928 -9201 10962 -9167
rect 11010 -9201 11044 -9167
rect 11082 -9201 11116 -9167
rect 11164 -9201 11198 -9167
rect 11236 -9201 11270 -9167
rect 11318 -9201 11352 -9167
rect 11390 -9201 11424 -9167
rect 11472 -9201 11506 -9167
rect 11544 -9201 11578 -9167
rect 11626 -9201 11660 -9167
rect 11698 -9201 11732 -9167
rect 11780 -9201 11814 -9167
rect 11852 -9201 11886 -9167
rect 11934 -9201 11968 -9167
rect 12006 -9201 12040 -9167
rect 4080 -9275 4114 -9241
rect 4152 -9275 4186 -9241
rect 4234 -9275 4268 -9241
rect 4306 -9275 4340 -9241
rect 4388 -9275 4422 -9241
rect 4460 -9275 4494 -9241
rect 4542 -9275 4576 -9241
rect 4614 -9275 4648 -9241
rect 4696 -9275 4730 -9241
rect 4768 -9275 4802 -9241
rect 4850 -9275 4884 -9241
rect 4922 -9275 4956 -9241
rect 5004 -9275 5038 -9241
rect 5076 -9275 5110 -9241
rect 5158 -9275 5192 -9241
rect 5230 -9275 5264 -9241
rect 5312 -9275 5346 -9241
rect 5384 -9275 5418 -9241
rect 5466 -9275 5500 -9241
rect 5538 -9275 5572 -9241
rect 5620 -9275 5654 -9241
rect 5692 -9275 5726 -9241
rect 5774 -9275 5808 -9241
rect 5846 -9275 5880 -9241
rect 5928 -9275 5962 -9241
rect 6000 -9275 6034 -9241
rect 6082 -9275 6116 -9241
rect 6154 -9275 6188 -9241
rect 6236 -9275 6270 -9241
rect 6308 -9275 6342 -9241
rect 6390 -9275 6424 -9241
rect 6462 -9275 6496 -9241
rect 6544 -9275 6578 -9241
rect 6616 -9275 6650 -9241
rect 6698 -9275 6732 -9241
rect 6770 -9275 6804 -9241
rect 6852 -9275 6886 -9241
rect 6924 -9275 6958 -9241
rect 7006 -9275 7040 -9241
rect 7078 -9275 7112 -9241
rect 7160 -9275 7194 -9241
rect 7232 -9275 7266 -9241
rect 7314 -9275 7348 -9241
rect 7386 -9275 7420 -9241
rect 7468 -9275 7502 -9241
rect 7540 -9275 7574 -9241
rect 7622 -9275 7656 -9241
rect 7694 -9275 7728 -9241
rect 7776 -9275 7810 -9241
rect 7848 -9275 7882 -9241
rect 7930 -9275 7964 -9241
rect 8002 -9275 8036 -9241
rect 8084 -9275 8118 -9241
rect 8156 -9275 8190 -9241
rect 8238 -9275 8272 -9241
rect 8310 -9275 8344 -9241
rect 8392 -9275 8426 -9241
rect 8464 -9275 8498 -9241
rect 8546 -9275 8580 -9241
rect 8618 -9275 8652 -9241
rect 8700 -9275 8734 -9241
rect 8772 -9275 8806 -9241
rect 8854 -9275 8888 -9241
rect 8926 -9275 8960 -9241
rect 9008 -9275 9042 -9241
rect 9080 -9275 9114 -9241
rect 9162 -9275 9196 -9241
rect 9234 -9275 9268 -9241
rect 9316 -9275 9350 -9241
rect 9388 -9275 9422 -9241
rect 9470 -9275 9504 -9241
rect 9542 -9275 9576 -9241
rect 9624 -9275 9658 -9241
rect 9696 -9275 9730 -9241
rect 9778 -9275 9812 -9241
rect 9850 -9275 9884 -9241
rect 9932 -9275 9966 -9241
rect 10004 -9275 10038 -9241
rect 10086 -9275 10120 -9241
rect 10158 -9275 10192 -9241
rect 10240 -9275 10274 -9241
rect 10312 -9275 10346 -9241
rect 10394 -9275 10428 -9241
rect 10466 -9275 10500 -9241
rect 10548 -9275 10582 -9241
rect 10620 -9275 10654 -9241
rect 10702 -9275 10736 -9241
rect 10774 -9275 10808 -9241
rect 10856 -9275 10890 -9241
rect 10928 -9275 10962 -9241
rect 11010 -9275 11044 -9241
rect 11082 -9275 11116 -9241
rect 11164 -9275 11198 -9241
rect 11236 -9275 11270 -9241
rect 11318 -9275 11352 -9241
rect 11390 -9275 11424 -9241
rect 11472 -9275 11506 -9241
rect 11544 -9275 11578 -9241
rect 11626 -9275 11660 -9241
rect 11698 -9275 11732 -9241
rect 11780 -9275 11814 -9241
rect 11852 -9275 11886 -9241
rect 11934 -9275 11968 -9241
rect 12006 -9275 12040 -9241
rect 4080 -9349 4114 -9315
rect 4152 -9349 4186 -9315
rect 4234 -9349 4268 -9315
rect 4306 -9349 4340 -9315
rect 4388 -9349 4422 -9315
rect 4460 -9349 4494 -9315
rect 4542 -9349 4576 -9315
rect 4614 -9349 4648 -9315
rect 4696 -9349 4730 -9315
rect 4768 -9349 4802 -9315
rect 4850 -9349 4884 -9315
rect 4922 -9349 4956 -9315
rect 5004 -9349 5038 -9315
rect 5076 -9349 5110 -9315
rect 5158 -9349 5192 -9315
rect 5230 -9349 5264 -9315
rect 5312 -9349 5346 -9315
rect 5384 -9349 5418 -9315
rect 5466 -9349 5500 -9315
rect 5538 -9349 5572 -9315
rect 5620 -9349 5654 -9315
rect 5692 -9349 5726 -9315
rect 5774 -9349 5808 -9315
rect 5846 -9349 5880 -9315
rect 5928 -9349 5962 -9315
rect 6000 -9349 6034 -9315
rect 6082 -9349 6116 -9315
rect 6154 -9349 6188 -9315
rect 6236 -9349 6270 -9315
rect 6308 -9349 6342 -9315
rect 6390 -9349 6424 -9315
rect 6462 -9349 6496 -9315
rect 6544 -9349 6578 -9315
rect 6616 -9349 6650 -9315
rect 6698 -9349 6732 -9315
rect 6770 -9349 6804 -9315
rect 6852 -9349 6886 -9315
rect 6924 -9349 6958 -9315
rect 7006 -9349 7040 -9315
rect 7078 -9349 7112 -9315
rect 7160 -9349 7194 -9315
rect 7232 -9349 7266 -9315
rect 7314 -9349 7348 -9315
rect 7386 -9349 7420 -9315
rect 7468 -9349 7502 -9315
rect 7540 -9349 7574 -9315
rect 7622 -9349 7656 -9315
rect 7694 -9349 7728 -9315
rect 7776 -9349 7810 -9315
rect 7848 -9349 7882 -9315
rect 7930 -9349 7964 -9315
rect 8002 -9349 8036 -9315
rect 8084 -9349 8118 -9315
rect 8156 -9349 8190 -9315
rect 8238 -9349 8272 -9315
rect 8310 -9349 8344 -9315
rect 8392 -9349 8426 -9315
rect 8464 -9349 8498 -9315
rect 8546 -9349 8580 -9315
rect 8618 -9349 8652 -9315
rect 8700 -9349 8734 -9315
rect 8772 -9349 8806 -9315
rect 8854 -9349 8888 -9315
rect 8926 -9349 8960 -9315
rect 9008 -9349 9042 -9315
rect 9080 -9349 9114 -9315
rect 9162 -9349 9196 -9315
rect 9234 -9349 9268 -9315
rect 9316 -9349 9350 -9315
rect 9388 -9349 9422 -9315
rect 9470 -9349 9504 -9315
rect 9542 -9349 9576 -9315
rect 9624 -9349 9658 -9315
rect 9696 -9349 9730 -9315
rect 9778 -9349 9812 -9315
rect 9850 -9349 9884 -9315
rect 9932 -9349 9966 -9315
rect 10004 -9349 10038 -9315
rect 10086 -9349 10120 -9315
rect 10158 -9349 10192 -9315
rect 10240 -9349 10274 -9315
rect 10312 -9349 10346 -9315
rect 10394 -9349 10428 -9315
rect 10466 -9349 10500 -9315
rect 10548 -9349 10582 -9315
rect 10620 -9349 10654 -9315
rect 10702 -9349 10736 -9315
rect 10774 -9349 10808 -9315
rect 10856 -9349 10890 -9315
rect 10928 -9349 10962 -9315
rect 11010 -9349 11044 -9315
rect 11082 -9349 11116 -9315
rect 11164 -9349 11198 -9315
rect 11236 -9349 11270 -9315
rect 11318 -9349 11352 -9315
rect 11390 -9349 11424 -9315
rect 11472 -9349 11506 -9315
rect 11544 -9349 11578 -9315
rect 11626 -9349 11660 -9315
rect 11698 -9349 11732 -9315
rect 11780 -9349 11814 -9315
rect 11852 -9349 11886 -9315
rect 11934 -9349 11968 -9315
rect 12006 -9349 12040 -9315
rect 4080 -9423 4114 -9389
rect 4152 -9423 4186 -9389
rect 4234 -9423 4268 -9389
rect 4306 -9423 4340 -9389
rect 4388 -9423 4422 -9389
rect 4460 -9423 4494 -9389
rect 4542 -9423 4576 -9389
rect 4614 -9423 4648 -9389
rect 4696 -9423 4730 -9389
rect 4768 -9423 4802 -9389
rect 4850 -9423 4884 -9389
rect 4922 -9423 4956 -9389
rect 5004 -9423 5038 -9389
rect 5076 -9423 5110 -9389
rect 5158 -9423 5192 -9389
rect 5230 -9423 5264 -9389
rect 5312 -9423 5346 -9389
rect 5384 -9423 5418 -9389
rect 5466 -9423 5500 -9389
rect 5538 -9423 5572 -9389
rect 5620 -9423 5654 -9389
rect 5692 -9423 5726 -9389
rect 5774 -9423 5808 -9389
rect 5846 -9423 5880 -9389
rect 5928 -9423 5962 -9389
rect 6000 -9423 6034 -9389
rect 6082 -9423 6116 -9389
rect 6154 -9423 6188 -9389
rect 6236 -9423 6270 -9389
rect 6308 -9423 6342 -9389
rect 6390 -9423 6424 -9389
rect 6462 -9423 6496 -9389
rect 6544 -9423 6578 -9389
rect 6616 -9423 6650 -9389
rect 6698 -9423 6732 -9389
rect 6770 -9423 6804 -9389
rect 6852 -9423 6886 -9389
rect 6924 -9423 6958 -9389
rect 7006 -9423 7040 -9389
rect 7078 -9423 7112 -9389
rect 7160 -9423 7194 -9389
rect 7232 -9423 7266 -9389
rect 7314 -9423 7348 -9389
rect 7386 -9423 7420 -9389
rect 7468 -9423 7502 -9389
rect 7540 -9423 7574 -9389
rect 7622 -9423 7656 -9389
rect 7694 -9423 7728 -9389
rect 7776 -9423 7810 -9389
rect 7848 -9423 7882 -9389
rect 7930 -9423 7964 -9389
rect 8002 -9423 8036 -9389
rect 8084 -9423 8118 -9389
rect 8156 -9423 8190 -9389
rect 8238 -9423 8272 -9389
rect 8310 -9423 8344 -9389
rect 8392 -9423 8426 -9389
rect 8464 -9423 8498 -9389
rect 8546 -9423 8580 -9389
rect 8618 -9423 8652 -9389
rect 8700 -9423 8734 -9389
rect 8772 -9423 8806 -9389
rect 8854 -9423 8888 -9389
rect 8926 -9423 8960 -9389
rect 9008 -9423 9042 -9389
rect 9080 -9423 9114 -9389
rect 9162 -9423 9196 -9389
rect 9234 -9423 9268 -9389
rect 9316 -9423 9350 -9389
rect 9388 -9423 9422 -9389
rect 9470 -9423 9504 -9389
rect 9542 -9423 9576 -9389
rect 9624 -9423 9658 -9389
rect 9696 -9423 9730 -9389
rect 9778 -9423 9812 -9389
rect 9850 -9423 9884 -9389
rect 9932 -9423 9966 -9389
rect 10004 -9423 10038 -9389
rect 10086 -9423 10120 -9389
rect 10158 -9423 10192 -9389
rect 10240 -9423 10274 -9389
rect 10312 -9423 10346 -9389
rect 10394 -9423 10428 -9389
rect 10466 -9423 10500 -9389
rect 10548 -9423 10582 -9389
rect 10620 -9423 10654 -9389
rect 10702 -9423 10736 -9389
rect 10774 -9423 10808 -9389
rect 10856 -9423 10890 -9389
rect 10928 -9423 10962 -9389
rect 11010 -9423 11044 -9389
rect 11082 -9423 11116 -9389
rect 11164 -9423 11198 -9389
rect 11236 -9423 11270 -9389
rect 11318 -9423 11352 -9389
rect 11390 -9423 11424 -9389
rect 11472 -9423 11506 -9389
rect 11544 -9423 11578 -9389
rect 11626 -9423 11660 -9389
rect 11698 -9423 11732 -9389
rect 11780 -9423 11814 -9389
rect 11852 -9423 11886 -9389
rect 11934 -9423 11968 -9389
rect 12006 -9423 12040 -9389
rect 4060 -9712 4094 -9678
rect 4134 -9712 4168 -9678
rect 4208 -9712 4242 -9678
rect 4282 -9712 4316 -9678
rect 4356 -9712 4390 -9678
rect 4430 -9712 4464 -9678
rect 4504 -9712 4538 -9678
rect 4578 -9712 4612 -9678
rect 4652 -9712 4686 -9678
rect 4726 -9712 4760 -9678
rect 4800 -9712 4834 -9678
rect 4874 -9712 4908 -9678
rect 4948 -9712 4982 -9678
rect 5022 -9712 5056 -9678
rect 5096 -9712 5130 -9678
rect 5170 -9712 5204 -9678
rect 5244 -9712 5278 -9678
rect 5318 -9712 5352 -9678
rect 5392 -9712 5426 -9678
rect 5466 -9712 5500 -9678
rect 5540 -9712 5574 -9678
rect 5614 -9712 5648 -9678
rect 5688 -9712 5722 -9678
rect 5762 -9712 5796 -9678
rect 5836 -9712 5870 -9678
rect 5910 -9712 5944 -9678
rect 5984 -9712 6018 -9678
rect 6058 -9712 6092 -9678
rect 6132 -9712 6166 -9678
rect 6206 -9712 6240 -9678
rect 6280 -9712 6314 -9678
rect 6354 -9712 6388 -9678
rect 6428 -9712 6462 -9678
rect 6502 -9712 6536 -9678
rect 6576 -9712 6610 -9678
rect 6650 -9712 6684 -9678
rect 6724 -9712 6758 -9678
rect 6798 -9712 6832 -9678
rect 6872 -9712 6906 -9678
rect 6946 -9712 6980 -9678
rect 7020 -9712 7054 -9678
rect 7094 -9712 7128 -9678
rect 7168 -9712 7202 -9678
rect 7242 -9712 7276 -9678
rect 7316 -9712 7350 -9678
rect 7390 -9712 7424 -9678
rect 7464 -9712 7498 -9678
rect 7538 -9712 7572 -9678
rect 7612 -9712 7646 -9678
rect 7686 -9712 7720 -9678
rect 7760 -9712 7794 -9678
rect 7834 -9712 7868 -9678
rect 7908 -9712 7942 -9678
rect 7982 -9712 8016 -9678
rect 8056 -9712 8090 -9678
rect 8130 -9712 8164 -9678
rect 8204 -9712 8238 -9678
rect 8278 -9712 8312 -9678
rect 8352 -9712 8386 -9678
rect 8426 -9712 8460 -9678
rect 8500 -9712 8534 -9678
rect 8574 -9712 8608 -9678
rect 8648 -9712 8682 -9678
rect 8722 -9712 8756 -9678
rect 8796 -9712 8830 -9678
rect 8870 -9712 8904 -9678
rect 8944 -9712 8978 -9678
rect 9018 -9712 9052 -9678
rect 9092 -9712 9126 -9678
rect 9166 -9712 9200 -9678
rect 9240 -9712 9274 -9678
rect 9314 -9712 9348 -9678
rect 9388 -9712 9422 -9678
rect 9462 -9712 9496 -9678
rect 9536 -9712 9570 -9678
rect 9610 -9712 9644 -9678
rect 9684 -9712 9718 -9678
rect 9758 -9712 9792 -9678
rect 9832 -9712 9866 -9678
rect 9906 -9712 9940 -9678
rect 9980 -9712 10014 -9678
rect 10054 -9712 10088 -9678
rect 10128 -9712 10162 -9678
rect 10202 -9712 10236 -9678
rect 10276 -9712 10310 -9678
rect 10350 -9712 10384 -9678
rect 10424 -9712 10458 -9678
rect 10498 -9712 10532 -9678
rect 10572 -9712 10606 -9678
rect 10646 -9712 10680 -9678
rect 10720 -9712 10754 -9678
rect 10794 -9712 10828 -9678
rect 10868 -9712 10902 -9678
rect 10942 -9712 10976 -9678
rect 11016 -9712 11050 -9678
rect 11090 -9712 11124 -9678
rect 11164 -9712 11198 -9678
rect 11238 -9712 11272 -9678
rect 11312 -9712 11346 -9678
rect 11386 -9712 11420 -9678
rect 11460 -9712 11494 -9678
rect 11534 -9712 11568 -9678
rect 11608 -9712 11642 -9678
rect 11682 -9712 11716 -9678
rect 11756 -9712 11790 -9678
rect 11830 -9712 11864 -9678
rect 11904 -9712 11938 -9678
rect 11978 -9712 12012 -9678
rect 12052 -9712 12086 -9678
rect 12126 -9712 12160 -9678
rect 12200 -9712 12234 -9678
rect 12274 -9712 12308 -9678
rect 12348 -9712 12382 -9678
rect 12422 -9712 12456 -9678
rect 12496 -9712 12530 -9678
rect 12570 -9712 12604 -9678
rect 12644 -9712 12678 -9678
rect 12718 -9712 12752 -9678
rect 12792 -9712 12826 -9678
rect 12866 -9712 12900 -9678
rect 12940 -9712 12974 -9678
rect 13014 -9712 13048 -9678
rect 13088 -9712 13122 -9678
rect 13162 -9712 13196 -9678
rect 13236 -9712 13270 -9678
rect 13310 -9712 13344 -9678
rect 13384 -9712 13418 -9678
rect 13458 -9712 13492 -9678
rect 13532 -9712 13566 -9678
rect 13606 -9712 13640 -9678
rect 13680 -9712 13714 -9678
rect 13754 -9712 13788 -9678
rect 13828 -9712 13862 -9678
rect 13902 -9712 13936 -9678
rect 13976 -9712 14010 -9678
rect 14050 -9712 14084 -9678
rect 14124 -9712 14158 -9678
rect 14198 -9712 14232 -9678
rect 14272 -9712 14306 -9678
rect 14346 -9712 14380 -9678
rect 14420 -9712 14454 -9678
rect 14494 -9712 14528 -9678
rect 14568 -9712 14602 -9678
rect 14642 -9712 14676 -9678
rect 14716 -9712 14750 -9678
rect 14790 -9712 14824 -9678
rect 14864 -9712 14898 -9678
rect 14938 -9712 14972 -9678
rect 15012 -9712 15046 -9678
rect 15086 -9712 15120 -9678
rect 15160 -9712 15194 -9678
rect 15234 -9712 15268 -9678
rect 15308 -9712 15342 -9678
rect 15382 -9712 15416 -9678
rect 15456 -9712 15490 -9678
rect 15530 -9712 15564 -9678
rect 15604 -9712 15638 -9678
rect 15678 -9712 15712 -9678
rect 15752 -9712 15786 -9678
rect 15826 -9712 15860 -9678
rect 15900 -9712 15934 -9678
rect 15974 -9712 16008 -9678
rect 16048 -9712 16082 -9678
rect 16122 -9712 16156 -9678
rect 16196 -9712 16230 -9678
rect 16270 -9712 16304 -9678
rect 16344 -9712 16378 -9678
rect 16418 -9712 16452 -9678
rect 16492 -9712 16526 -9678
rect 16566 -9712 16600 -9678
rect 16640 -9712 16674 -9678
rect 16714 -9712 16748 -9678
rect 16788 -9712 16822 -9678
rect 16862 -9712 16896 -9678
rect 16936 -9712 16970 -9678
rect 17010 -9712 17044 -9678
rect 17084 -9712 17118 -9678
rect 17158 -9712 17192 -9678
rect 17232 -9712 17266 -9678
rect 17306 -9712 17340 -9678
rect 17380 -9712 17414 -9678
rect 17454 -9712 17488 -9678
rect 17528 -9712 17562 -9678
rect 17602 -9712 17636 -9678
rect 17676 -9712 17710 -9678
rect 17750 -9712 17784 -9678
rect 17824 -9712 17858 -9678
rect 17898 -9712 17932 -9678
rect 17972 -9712 18006 -9678
rect 18046 -9712 18080 -9678
rect 18120 -9712 18154 -9678
rect 18194 -9712 18228 -9678
rect 18268 -9712 18302 -9678
rect 18342 -9712 18376 -9678
rect 18416 -9712 18450 -9678
rect 18490 -9712 18524 -9678
rect 18564 -9712 18598 -9678
rect 18638 -9712 18672 -9678
rect 18712 -9712 18746 -9678
rect 18786 -9712 18820 -9678
rect 18860 -9712 18894 -9678
rect 18934 -9712 18968 -9678
rect 19008 -9712 19042 -9678
rect 19082 -9712 19116 -9678
rect 19156 -9712 19190 -9678
rect 19230 -9712 19264 -9678
rect 19304 -9712 19338 -9678
rect 19378 -9712 19412 -9678
rect 19452 -9712 19486 -9678
rect 19526 -9712 19560 -9678
rect 19600 -9712 19634 -9678
rect 19674 -9712 19708 -9678
rect 19748 -9712 19782 -9678
rect 19822 -9712 19856 -9678
rect 19896 -9712 19930 -9678
rect 19970 -9712 20004 -9678
rect 20044 -9712 20078 -9678
rect 20118 -9712 20152 -9678
rect 20192 -9712 20226 -9678
rect 20266 -9712 20300 -9678
rect 20340 -9712 20374 -9678
rect 20414 -9712 20448 -9678
rect 20488 -9712 20522 -9678
rect 20562 -9712 20596 -9678
rect 20636 -9712 20670 -9678
rect 20710 -9712 20744 -9678
rect 20784 -9712 20818 -9678
rect 20858 -9712 20892 -9678
rect 20932 -9712 20966 -9678
rect 21006 -9712 21040 -9678
rect 21080 -9712 21114 -9678
rect 21154 -9712 21188 -9678
rect 21228 -9712 21262 -9678
rect 21302 -9712 21336 -9678
rect 21376 -9712 21410 -9678
rect 21450 -9712 21484 -9678
rect 21524 -9712 21558 -9678
rect 21598 -9712 21632 -9678
rect 21672 -9712 21706 -9678
rect 21746 -9712 21780 -9678
rect 21820 -9712 21854 -9678
rect 21894 -9712 21928 -9678
rect 21968 -9712 22002 -9678
rect 22042 -9712 22076 -9678
rect 22116 -9712 22150 -9678
rect 22190 -9712 22224 -9678
rect 22264 -9712 22298 -9678
rect 22338 -9712 22372 -9678
rect 22412 -9712 22446 -9678
rect 22486 -9712 22520 -9678
rect 22560 -9712 22594 -9678
rect 22634 -9712 22668 -9678
rect 22708 -9712 22742 -9678
rect 22782 -9712 22816 -9678
rect 22856 -9712 22890 -9678
rect 22930 -9712 22964 -9678
rect 23004 -9712 23038 -9678
rect 23078 -9712 23112 -9678
rect 23152 -9712 23186 -9678
rect 23226 -9712 23260 -9678
rect 23300 -9712 23334 -9678
rect 23374 -9712 23408 -9678
rect 23448 -9712 23482 -9678
rect 23522 -9712 23556 -9678
rect 23596 -9712 23630 -9678
rect 23670 -9712 23704 -9678
rect 23744 -9712 23778 -9678
rect 23818 -9712 23852 -9678
rect 23892 -9712 23926 -9678
rect 23966 -9712 24000 -9678
rect 24040 -9712 24074 -9678
rect 24114 -9712 24148 -9678
rect 24188 -9712 24222 -9678
rect 24262 -9712 24296 -9678
rect 24336 -9712 24370 -9678
rect 24410 -9712 24444 -9678
rect 24484 -9712 24518 -9678
rect 24558 -9712 24592 -9678
rect 24632 -9712 24666 -9678
rect 24706 -9712 24740 -9678
rect 24780 -9712 24814 -9678
rect 24854 -9712 24888 -9678
rect 24928 -9712 24962 -9678
rect 25002 -9712 25036 -9678
rect 25076 -9712 25110 -9678
rect 25150 -9712 25184 -9678
rect 4060 -9786 4094 -9752
rect 4134 -9786 4168 -9752
rect 4208 -9786 4242 -9752
rect 4282 -9786 4316 -9752
rect 4356 -9786 4390 -9752
rect 4430 -9786 4464 -9752
rect 4504 -9786 4538 -9752
rect 4578 -9786 4612 -9752
rect 4652 -9786 4686 -9752
rect 4726 -9786 4760 -9752
rect 4800 -9786 4834 -9752
rect 4874 -9786 4908 -9752
rect 4948 -9786 4982 -9752
rect 5022 -9786 5056 -9752
rect 5096 -9786 5130 -9752
rect 5170 -9786 5204 -9752
rect 5244 -9786 5278 -9752
rect 5318 -9786 5352 -9752
rect 5392 -9786 5426 -9752
rect 5466 -9786 5500 -9752
rect 5540 -9786 5574 -9752
rect 5614 -9786 5648 -9752
rect 5688 -9786 5722 -9752
rect 5762 -9786 5796 -9752
rect 5836 -9786 5870 -9752
rect 5910 -9786 5944 -9752
rect 5984 -9786 6018 -9752
rect 6058 -9786 6092 -9752
rect 6132 -9786 6166 -9752
rect 6206 -9786 6240 -9752
rect 6280 -9786 6314 -9752
rect 6354 -9786 6388 -9752
rect 6428 -9786 6462 -9752
rect 6502 -9786 6536 -9752
rect 6576 -9786 6610 -9752
rect 6650 -9786 6684 -9752
rect 6724 -9786 6758 -9752
rect 6798 -9786 6832 -9752
rect 6872 -9786 6906 -9752
rect 6946 -9786 6980 -9752
rect 7020 -9786 7054 -9752
rect 7094 -9786 7128 -9752
rect 7168 -9786 7202 -9752
rect 7242 -9786 7276 -9752
rect 7316 -9786 7350 -9752
rect 7390 -9786 7424 -9752
rect 7464 -9786 7498 -9752
rect 7538 -9786 7572 -9752
rect 7612 -9786 7646 -9752
rect 7686 -9786 7720 -9752
rect 7760 -9786 7794 -9752
rect 7834 -9786 7868 -9752
rect 7908 -9786 7942 -9752
rect 7982 -9786 8016 -9752
rect 8056 -9786 8090 -9752
rect 8130 -9786 8164 -9752
rect 8204 -9786 8238 -9752
rect 8278 -9786 8312 -9752
rect 8352 -9786 8386 -9752
rect 8426 -9786 8460 -9752
rect 8500 -9786 8534 -9752
rect 8574 -9786 8608 -9752
rect 8648 -9786 8682 -9752
rect 8722 -9786 8756 -9752
rect 8796 -9786 8830 -9752
rect 8870 -9786 8904 -9752
rect 8944 -9786 8978 -9752
rect 9018 -9786 9052 -9752
rect 9092 -9786 9126 -9752
rect 9166 -9786 9200 -9752
rect 9240 -9786 9274 -9752
rect 9314 -9786 9348 -9752
rect 9388 -9786 9422 -9752
rect 9462 -9786 9496 -9752
rect 9536 -9786 9570 -9752
rect 9610 -9786 9644 -9752
rect 9684 -9786 9718 -9752
rect 9758 -9786 9792 -9752
rect 9832 -9786 9866 -9752
rect 9906 -9786 9940 -9752
rect 9980 -9786 10014 -9752
rect 10054 -9786 10088 -9752
rect 10128 -9786 10162 -9752
rect 10202 -9786 10236 -9752
rect 10276 -9786 10310 -9752
rect 10350 -9786 10384 -9752
rect 10424 -9786 10458 -9752
rect 10498 -9786 10532 -9752
rect 10572 -9786 10606 -9752
rect 10646 -9786 10680 -9752
rect 10720 -9786 10754 -9752
rect 10794 -9786 10828 -9752
rect 10868 -9786 10902 -9752
rect 10942 -9786 10976 -9752
rect 11016 -9786 11050 -9752
rect 11090 -9786 11124 -9752
rect 11164 -9786 11198 -9752
rect 11238 -9786 11272 -9752
rect 11312 -9786 11346 -9752
rect 11386 -9786 11420 -9752
rect 11460 -9786 11494 -9752
rect 11534 -9786 11568 -9752
rect 11608 -9786 11642 -9752
rect 11682 -9786 11716 -9752
rect 11756 -9786 11790 -9752
rect 11830 -9786 11864 -9752
rect 11904 -9786 11938 -9752
rect 11978 -9786 12012 -9752
rect 12052 -9786 12086 -9752
rect 12126 -9786 12160 -9752
rect 12200 -9786 12234 -9752
rect 12274 -9786 12308 -9752
rect 12348 -9786 12382 -9752
rect 12422 -9786 12456 -9752
rect 12496 -9786 12530 -9752
rect 12570 -9786 12604 -9752
rect 12644 -9786 12678 -9752
rect 12718 -9786 12752 -9752
rect 12792 -9786 12826 -9752
rect 12866 -9786 12900 -9752
rect 12940 -9786 12974 -9752
rect 13014 -9786 13048 -9752
rect 13088 -9786 13122 -9752
rect 13162 -9786 13196 -9752
rect 13236 -9786 13270 -9752
rect 13310 -9786 13344 -9752
rect 13384 -9786 13418 -9752
rect 13458 -9786 13492 -9752
rect 13532 -9786 13566 -9752
rect 13606 -9786 13640 -9752
rect 13680 -9786 13714 -9752
rect 13754 -9786 13788 -9752
rect 13828 -9786 13862 -9752
rect 13902 -9786 13936 -9752
rect 13976 -9786 14010 -9752
rect 14050 -9786 14084 -9752
rect 14124 -9786 14158 -9752
rect 14198 -9786 14232 -9752
rect 14272 -9786 14306 -9752
rect 14346 -9786 14380 -9752
rect 14420 -9786 14454 -9752
rect 14494 -9786 14528 -9752
rect 14568 -9786 14602 -9752
rect 14642 -9786 14676 -9752
rect 14716 -9786 14750 -9752
rect 14790 -9786 14824 -9752
rect 14864 -9786 14898 -9752
rect 14938 -9786 14972 -9752
rect 15012 -9786 15046 -9752
rect 15086 -9786 15120 -9752
rect 15160 -9786 15194 -9752
rect 15234 -9786 15268 -9752
rect 15308 -9786 15342 -9752
rect 15382 -9786 15416 -9752
rect 15456 -9786 15490 -9752
rect 15530 -9786 15564 -9752
rect 15604 -9786 15638 -9752
rect 15678 -9786 15712 -9752
rect 15752 -9786 15786 -9752
rect 15826 -9786 15860 -9752
rect 15900 -9786 15934 -9752
rect 15974 -9786 16008 -9752
rect 16048 -9786 16082 -9752
rect 16122 -9786 16156 -9752
rect 16196 -9786 16230 -9752
rect 16270 -9786 16304 -9752
rect 16344 -9786 16378 -9752
rect 16418 -9786 16452 -9752
rect 16492 -9786 16526 -9752
rect 16566 -9786 16600 -9752
rect 16640 -9786 16674 -9752
rect 16714 -9786 16748 -9752
rect 16788 -9786 16822 -9752
rect 16862 -9786 16896 -9752
rect 16936 -9786 16970 -9752
rect 17010 -9786 17044 -9752
rect 17084 -9786 17118 -9752
rect 17158 -9786 17192 -9752
rect 17232 -9786 17266 -9752
rect 17306 -9786 17340 -9752
rect 17380 -9786 17414 -9752
rect 17454 -9786 17488 -9752
rect 17528 -9786 17562 -9752
rect 17602 -9786 17636 -9752
rect 17676 -9786 17710 -9752
rect 17750 -9786 17784 -9752
rect 17824 -9786 17858 -9752
rect 17898 -9786 17932 -9752
rect 17972 -9786 18006 -9752
rect 18046 -9786 18080 -9752
rect 18120 -9786 18154 -9752
rect 18194 -9786 18228 -9752
rect 18268 -9786 18302 -9752
rect 18342 -9786 18376 -9752
rect 18416 -9786 18450 -9752
rect 18490 -9786 18524 -9752
rect 18564 -9786 18598 -9752
rect 18638 -9786 18672 -9752
rect 18712 -9786 18746 -9752
rect 18786 -9786 18820 -9752
rect 18860 -9786 18894 -9752
rect 18934 -9786 18968 -9752
rect 19008 -9786 19042 -9752
rect 19082 -9786 19116 -9752
rect 19156 -9786 19190 -9752
rect 19230 -9786 19264 -9752
rect 19304 -9786 19338 -9752
rect 19378 -9786 19412 -9752
rect 19452 -9786 19486 -9752
rect 19526 -9786 19560 -9752
rect 19600 -9786 19634 -9752
rect 19674 -9786 19708 -9752
rect 19748 -9786 19782 -9752
rect 19822 -9786 19856 -9752
rect 19896 -9786 19930 -9752
rect 19970 -9786 20004 -9752
rect 20044 -9786 20078 -9752
rect 20118 -9786 20152 -9752
rect 20192 -9786 20226 -9752
rect 20266 -9786 20300 -9752
rect 20340 -9786 20374 -9752
rect 20414 -9786 20448 -9752
rect 20488 -9786 20522 -9752
rect 20562 -9786 20596 -9752
rect 20636 -9786 20670 -9752
rect 20710 -9786 20744 -9752
rect 20784 -9786 20818 -9752
rect 20858 -9786 20892 -9752
rect 20932 -9786 20966 -9752
rect 21006 -9786 21040 -9752
rect 21080 -9786 21114 -9752
rect 21154 -9786 21188 -9752
rect 21228 -9786 21262 -9752
rect 21302 -9786 21336 -9752
rect 21376 -9786 21410 -9752
rect 21450 -9786 21484 -9752
rect 21524 -9786 21558 -9752
rect 21598 -9786 21632 -9752
rect 21672 -9786 21706 -9752
rect 21746 -9786 21780 -9752
rect 21820 -9786 21854 -9752
rect 21894 -9786 21928 -9752
rect 21968 -9786 22002 -9752
rect 22042 -9786 22076 -9752
rect 22116 -9786 22150 -9752
rect 22190 -9786 22224 -9752
rect 22264 -9786 22298 -9752
rect 22338 -9786 22372 -9752
rect 22412 -9786 22446 -9752
rect 22486 -9786 22520 -9752
rect 22560 -9786 22594 -9752
rect 22634 -9786 22668 -9752
rect 22708 -9786 22742 -9752
rect 22782 -9786 22816 -9752
rect 22856 -9786 22890 -9752
rect 22930 -9786 22964 -9752
rect 23004 -9786 23038 -9752
rect 23078 -9786 23112 -9752
rect 23152 -9786 23186 -9752
rect 23226 -9786 23260 -9752
rect 23300 -9786 23334 -9752
rect 23374 -9786 23408 -9752
rect 23448 -9786 23482 -9752
rect 23522 -9786 23556 -9752
rect 23596 -9786 23630 -9752
rect 23670 -9786 23704 -9752
rect 23744 -9786 23778 -9752
rect 23818 -9786 23852 -9752
rect 23892 -9786 23926 -9752
rect 23966 -9786 24000 -9752
rect 24040 -9786 24074 -9752
rect 24114 -9786 24148 -9752
rect 24188 -9786 24222 -9752
rect 24262 -9786 24296 -9752
rect 24336 -9786 24370 -9752
rect 24410 -9786 24444 -9752
rect 24484 -9786 24518 -9752
rect 24558 -9786 24592 -9752
rect 24632 -9786 24666 -9752
rect 24706 -9786 24740 -9752
rect 24780 -9786 24814 -9752
rect 24854 -9786 24888 -9752
rect 24928 -9786 24962 -9752
rect 25002 -9786 25036 -9752
rect 25076 -9786 25110 -9752
rect 25150 -9786 25184 -9752
rect 4060 -9860 4094 -9826
rect 4134 -9860 4168 -9826
rect 4208 -9860 4242 -9826
rect 4282 -9860 4316 -9826
rect 4356 -9860 4390 -9826
rect 4430 -9860 4464 -9826
rect 4504 -9860 4538 -9826
rect 4578 -9860 4612 -9826
rect 4652 -9860 4686 -9826
rect 4726 -9860 4760 -9826
rect 4800 -9860 4834 -9826
rect 4874 -9860 4908 -9826
rect 4948 -9860 4982 -9826
rect 5022 -9860 5056 -9826
rect 5096 -9860 5130 -9826
rect 5170 -9860 5204 -9826
rect 5244 -9860 5278 -9826
rect 5318 -9860 5352 -9826
rect 5392 -9860 5426 -9826
rect 5466 -9860 5500 -9826
rect 5540 -9860 5574 -9826
rect 5614 -9860 5648 -9826
rect 5688 -9860 5722 -9826
rect 5762 -9860 5796 -9826
rect 5836 -9860 5870 -9826
rect 5910 -9860 5944 -9826
rect 5984 -9860 6018 -9826
rect 6058 -9860 6092 -9826
rect 6132 -9860 6166 -9826
rect 6206 -9860 6240 -9826
rect 6280 -9860 6314 -9826
rect 6354 -9860 6388 -9826
rect 6428 -9860 6462 -9826
rect 6502 -9860 6536 -9826
rect 6576 -9860 6610 -9826
rect 6650 -9860 6684 -9826
rect 6724 -9860 6758 -9826
rect 6798 -9860 6832 -9826
rect 6872 -9860 6906 -9826
rect 6946 -9860 6980 -9826
rect 7020 -9860 7054 -9826
rect 7094 -9860 7128 -9826
rect 7168 -9860 7202 -9826
rect 7242 -9860 7276 -9826
rect 7316 -9860 7350 -9826
rect 7390 -9860 7424 -9826
rect 7464 -9860 7498 -9826
rect 7538 -9860 7572 -9826
rect 7612 -9860 7646 -9826
rect 7686 -9860 7720 -9826
rect 7760 -9860 7794 -9826
rect 7834 -9860 7868 -9826
rect 7908 -9860 7942 -9826
rect 7982 -9860 8016 -9826
rect 8056 -9860 8090 -9826
rect 8130 -9860 8164 -9826
rect 8204 -9860 8238 -9826
rect 8278 -9860 8312 -9826
rect 8352 -9860 8386 -9826
rect 8426 -9860 8460 -9826
rect 8500 -9860 8534 -9826
rect 8574 -9860 8608 -9826
rect 8648 -9860 8682 -9826
rect 8722 -9860 8756 -9826
rect 8796 -9860 8830 -9826
rect 8870 -9860 8904 -9826
rect 8944 -9860 8978 -9826
rect 9018 -9860 9052 -9826
rect 9092 -9860 9126 -9826
rect 9166 -9860 9200 -9826
rect 9240 -9860 9274 -9826
rect 9314 -9860 9348 -9826
rect 9388 -9860 9422 -9826
rect 9462 -9860 9496 -9826
rect 9536 -9860 9570 -9826
rect 9610 -9860 9644 -9826
rect 9684 -9860 9718 -9826
rect 9758 -9860 9792 -9826
rect 9832 -9860 9866 -9826
rect 9906 -9860 9940 -9826
rect 9980 -9860 10014 -9826
rect 10054 -9860 10088 -9826
rect 10128 -9860 10162 -9826
rect 10202 -9860 10236 -9826
rect 10276 -9860 10310 -9826
rect 10350 -9860 10384 -9826
rect 10424 -9860 10458 -9826
rect 10498 -9860 10532 -9826
rect 10572 -9860 10606 -9826
rect 10646 -9860 10680 -9826
rect 10720 -9860 10754 -9826
rect 10794 -9860 10828 -9826
rect 10868 -9860 10902 -9826
rect 10942 -9860 10976 -9826
rect 11016 -9860 11050 -9826
rect 11090 -9860 11124 -9826
rect 11164 -9860 11198 -9826
rect 11238 -9860 11272 -9826
rect 11312 -9860 11346 -9826
rect 11386 -9860 11420 -9826
rect 11460 -9860 11494 -9826
rect 11534 -9860 11568 -9826
rect 11608 -9860 11642 -9826
rect 11682 -9860 11716 -9826
rect 11756 -9860 11790 -9826
rect 11830 -9860 11864 -9826
rect 11904 -9860 11938 -9826
rect 11978 -9860 12012 -9826
rect 12052 -9860 12086 -9826
rect 12126 -9860 12160 -9826
rect 12200 -9860 12234 -9826
rect 12274 -9860 12308 -9826
rect 12348 -9860 12382 -9826
rect 12422 -9860 12456 -9826
rect 12496 -9860 12530 -9826
rect 12570 -9860 12604 -9826
rect 12644 -9860 12678 -9826
rect 12718 -9860 12752 -9826
rect 12792 -9860 12826 -9826
rect 12866 -9860 12900 -9826
rect 12940 -9860 12974 -9826
rect 13014 -9860 13048 -9826
rect 13088 -9860 13122 -9826
rect 13162 -9860 13196 -9826
rect 13236 -9860 13270 -9826
rect 13310 -9860 13344 -9826
rect 13384 -9860 13418 -9826
rect 13458 -9860 13492 -9826
rect 13532 -9860 13566 -9826
rect 13606 -9860 13640 -9826
rect 13680 -9860 13714 -9826
rect 13754 -9860 13788 -9826
rect 13828 -9860 13862 -9826
rect 13902 -9860 13936 -9826
rect 13976 -9860 14010 -9826
rect 14050 -9860 14084 -9826
rect 14124 -9860 14158 -9826
rect 14198 -9860 14232 -9826
rect 14272 -9860 14306 -9826
rect 14346 -9860 14380 -9826
rect 14420 -9860 14454 -9826
rect 14494 -9860 14528 -9826
rect 14568 -9860 14602 -9826
rect 14642 -9860 14676 -9826
rect 14716 -9860 14750 -9826
rect 14790 -9860 14824 -9826
rect 14864 -9860 14898 -9826
rect 14938 -9860 14972 -9826
rect 15012 -9860 15046 -9826
rect 15086 -9860 15120 -9826
rect 15160 -9860 15194 -9826
rect 15234 -9860 15268 -9826
rect 15308 -9860 15342 -9826
rect 15382 -9860 15416 -9826
rect 15456 -9860 15490 -9826
rect 15530 -9860 15564 -9826
rect 15604 -9860 15638 -9826
rect 15678 -9860 15712 -9826
rect 15752 -9860 15786 -9826
rect 15826 -9860 15860 -9826
rect 15900 -9860 15934 -9826
rect 15974 -9860 16008 -9826
rect 16048 -9860 16082 -9826
rect 16122 -9860 16156 -9826
rect 16196 -9860 16230 -9826
rect 16270 -9860 16304 -9826
rect 16344 -9860 16378 -9826
rect 16418 -9860 16452 -9826
rect 16492 -9860 16526 -9826
rect 16566 -9860 16600 -9826
rect 16640 -9860 16674 -9826
rect 16714 -9860 16748 -9826
rect 16788 -9860 16822 -9826
rect 16862 -9860 16896 -9826
rect 16936 -9860 16970 -9826
rect 17010 -9860 17044 -9826
rect 17084 -9860 17118 -9826
rect 17158 -9860 17192 -9826
rect 17232 -9860 17266 -9826
rect 17306 -9860 17340 -9826
rect 17380 -9860 17414 -9826
rect 17454 -9860 17488 -9826
rect 17528 -9860 17562 -9826
rect 17602 -9860 17636 -9826
rect 17676 -9860 17710 -9826
rect 17750 -9860 17784 -9826
rect 17824 -9860 17858 -9826
rect 17898 -9860 17932 -9826
rect 17972 -9860 18006 -9826
rect 18046 -9860 18080 -9826
rect 18120 -9860 18154 -9826
rect 18194 -9860 18228 -9826
rect 18268 -9860 18302 -9826
rect 18342 -9860 18376 -9826
rect 18416 -9860 18450 -9826
rect 18490 -9860 18524 -9826
rect 18564 -9860 18598 -9826
rect 18638 -9860 18672 -9826
rect 18712 -9860 18746 -9826
rect 18786 -9860 18820 -9826
rect 18860 -9860 18894 -9826
rect 18934 -9860 18968 -9826
rect 19008 -9860 19042 -9826
rect 19082 -9860 19116 -9826
rect 19156 -9860 19190 -9826
rect 19230 -9860 19264 -9826
rect 19304 -9860 19338 -9826
rect 19378 -9860 19412 -9826
rect 19452 -9860 19486 -9826
rect 19526 -9860 19560 -9826
rect 19600 -9860 19634 -9826
rect 19674 -9860 19708 -9826
rect 19748 -9860 19782 -9826
rect 19822 -9860 19856 -9826
rect 19896 -9860 19930 -9826
rect 19970 -9860 20004 -9826
rect 20044 -9860 20078 -9826
rect 20118 -9860 20152 -9826
rect 20192 -9860 20226 -9826
rect 20266 -9860 20300 -9826
rect 20340 -9860 20374 -9826
rect 20414 -9860 20448 -9826
rect 20488 -9860 20522 -9826
rect 20562 -9860 20596 -9826
rect 20636 -9860 20670 -9826
rect 20710 -9860 20744 -9826
rect 20784 -9860 20818 -9826
rect 20858 -9860 20892 -9826
rect 20932 -9860 20966 -9826
rect 21006 -9860 21040 -9826
rect 21080 -9860 21114 -9826
rect 21154 -9860 21188 -9826
rect 21228 -9860 21262 -9826
rect 21302 -9860 21336 -9826
rect 21376 -9860 21410 -9826
rect 21450 -9860 21484 -9826
rect 21524 -9860 21558 -9826
rect 21598 -9860 21632 -9826
rect 21672 -9860 21706 -9826
rect 21746 -9860 21780 -9826
rect 21820 -9860 21854 -9826
rect 21894 -9860 21928 -9826
rect 21968 -9860 22002 -9826
rect 22042 -9860 22076 -9826
rect 22116 -9860 22150 -9826
rect 22190 -9860 22224 -9826
rect 22264 -9860 22298 -9826
rect 22338 -9860 22372 -9826
rect 22412 -9860 22446 -9826
rect 22486 -9860 22520 -9826
rect 22560 -9860 22594 -9826
rect 22634 -9860 22668 -9826
rect 22708 -9860 22742 -9826
rect 22782 -9860 22816 -9826
rect 22856 -9860 22890 -9826
rect 22930 -9860 22964 -9826
rect 23004 -9860 23038 -9826
rect 23078 -9860 23112 -9826
rect 23152 -9860 23186 -9826
rect 23226 -9860 23260 -9826
rect 23300 -9860 23334 -9826
rect 23374 -9860 23408 -9826
rect 23448 -9860 23482 -9826
rect 23522 -9860 23556 -9826
rect 23596 -9860 23630 -9826
rect 23670 -9860 23704 -9826
rect 23744 -9860 23778 -9826
rect 23818 -9860 23852 -9826
rect 23892 -9860 23926 -9826
rect 23966 -9860 24000 -9826
rect 24040 -9860 24074 -9826
rect 24114 -9860 24148 -9826
rect 24188 -9860 24222 -9826
rect 24262 -9860 24296 -9826
rect 24336 -9860 24370 -9826
rect 24410 -9860 24444 -9826
rect 24484 -9860 24518 -9826
rect 24558 -9860 24592 -9826
rect 24632 -9860 24666 -9826
rect 24706 -9860 24740 -9826
rect 24780 -9860 24814 -9826
rect 24854 -9860 24888 -9826
rect 24928 -9860 24962 -9826
rect 25002 -9860 25036 -9826
rect 25076 -9860 25110 -9826
rect 25150 -9860 25184 -9826
rect 4060 -9934 4094 -9900
rect 4134 -9934 4168 -9900
rect 4208 -9934 4242 -9900
rect 4282 -9934 4316 -9900
rect 4356 -9934 4390 -9900
rect 4430 -9934 4464 -9900
rect 4504 -9934 4538 -9900
rect 4578 -9934 4612 -9900
rect 4652 -9934 4686 -9900
rect 4726 -9934 4760 -9900
rect 4800 -9934 4834 -9900
rect 4874 -9934 4908 -9900
rect 4948 -9934 4982 -9900
rect 5022 -9934 5056 -9900
rect 5096 -9934 5130 -9900
rect 5170 -9934 5204 -9900
rect 5244 -9934 5278 -9900
rect 5318 -9934 5352 -9900
rect 5392 -9934 5426 -9900
rect 5466 -9934 5500 -9900
rect 5540 -9934 5574 -9900
rect 5614 -9934 5648 -9900
rect 5688 -9934 5722 -9900
rect 5762 -9934 5796 -9900
rect 5836 -9934 5870 -9900
rect 5910 -9934 5944 -9900
rect 5984 -9934 6018 -9900
rect 6058 -9934 6092 -9900
rect 6132 -9934 6166 -9900
rect 6206 -9934 6240 -9900
rect 6280 -9934 6314 -9900
rect 6354 -9934 6388 -9900
rect 6428 -9934 6462 -9900
rect 6502 -9934 6536 -9900
rect 6576 -9934 6610 -9900
rect 6650 -9934 6684 -9900
rect 6724 -9934 6758 -9900
rect 6798 -9934 6832 -9900
rect 6872 -9934 6906 -9900
rect 6946 -9934 6980 -9900
rect 7020 -9934 7054 -9900
rect 7094 -9934 7128 -9900
rect 7168 -9934 7202 -9900
rect 7242 -9934 7276 -9900
rect 7316 -9934 7350 -9900
rect 7390 -9934 7424 -9900
rect 7464 -9934 7498 -9900
rect 7538 -9934 7572 -9900
rect 7612 -9934 7646 -9900
rect 7686 -9934 7720 -9900
rect 7760 -9934 7794 -9900
rect 7834 -9934 7868 -9900
rect 7908 -9934 7942 -9900
rect 7982 -9934 8016 -9900
rect 8056 -9934 8090 -9900
rect 8130 -9934 8164 -9900
rect 8204 -9934 8238 -9900
rect 8278 -9934 8312 -9900
rect 8352 -9934 8386 -9900
rect 8426 -9934 8460 -9900
rect 8500 -9934 8534 -9900
rect 8574 -9934 8608 -9900
rect 8648 -9934 8682 -9900
rect 8722 -9934 8756 -9900
rect 8796 -9934 8830 -9900
rect 8870 -9934 8904 -9900
rect 8944 -9934 8978 -9900
rect 9018 -9934 9052 -9900
rect 9092 -9934 9126 -9900
rect 9166 -9934 9200 -9900
rect 9240 -9934 9274 -9900
rect 9314 -9934 9348 -9900
rect 9388 -9934 9422 -9900
rect 9462 -9934 9496 -9900
rect 9536 -9934 9570 -9900
rect 9610 -9934 9644 -9900
rect 9684 -9934 9718 -9900
rect 9758 -9934 9792 -9900
rect 9832 -9934 9866 -9900
rect 9906 -9934 9940 -9900
rect 9980 -9934 10014 -9900
rect 10054 -9934 10088 -9900
rect 10128 -9934 10162 -9900
rect 10202 -9934 10236 -9900
rect 10276 -9934 10310 -9900
rect 10350 -9934 10384 -9900
rect 10424 -9934 10458 -9900
rect 10498 -9934 10532 -9900
rect 10572 -9934 10606 -9900
rect 10646 -9934 10680 -9900
rect 10720 -9934 10754 -9900
rect 10794 -9934 10828 -9900
rect 10868 -9934 10902 -9900
rect 10942 -9934 10976 -9900
rect 11016 -9934 11050 -9900
rect 11090 -9934 11124 -9900
rect 11164 -9934 11198 -9900
rect 11238 -9934 11272 -9900
rect 11312 -9934 11346 -9900
rect 11386 -9934 11420 -9900
rect 11460 -9934 11494 -9900
rect 11534 -9934 11568 -9900
rect 11608 -9934 11642 -9900
rect 11682 -9934 11716 -9900
rect 11756 -9934 11790 -9900
rect 11830 -9934 11864 -9900
rect 11904 -9934 11938 -9900
rect 11978 -9934 12012 -9900
rect 12052 -9934 12086 -9900
rect 12126 -9934 12160 -9900
rect 12200 -9934 12234 -9900
rect 12274 -9934 12308 -9900
rect 12348 -9934 12382 -9900
rect 12422 -9934 12456 -9900
rect 12496 -9934 12530 -9900
rect 12570 -9934 12604 -9900
rect 12644 -9934 12678 -9900
rect 12718 -9934 12752 -9900
rect 12792 -9934 12826 -9900
rect 12866 -9934 12900 -9900
rect 12940 -9934 12974 -9900
rect 13014 -9934 13048 -9900
rect 13088 -9934 13122 -9900
rect 13162 -9934 13196 -9900
rect 13236 -9934 13270 -9900
rect 13310 -9934 13344 -9900
rect 13384 -9934 13418 -9900
rect 13458 -9934 13492 -9900
rect 13532 -9934 13566 -9900
rect 13606 -9934 13640 -9900
rect 13680 -9934 13714 -9900
rect 13754 -9934 13788 -9900
rect 13828 -9934 13862 -9900
rect 13902 -9934 13936 -9900
rect 13976 -9934 14010 -9900
rect 14050 -9934 14084 -9900
rect 14124 -9934 14158 -9900
rect 14198 -9934 14232 -9900
rect 14272 -9934 14306 -9900
rect 14346 -9934 14380 -9900
rect 14420 -9934 14454 -9900
rect 14494 -9934 14528 -9900
rect 14568 -9934 14602 -9900
rect 14642 -9934 14676 -9900
rect 14716 -9934 14750 -9900
rect 14790 -9934 14824 -9900
rect 14864 -9934 14898 -9900
rect 14938 -9934 14972 -9900
rect 15012 -9934 15046 -9900
rect 15086 -9934 15120 -9900
rect 15160 -9934 15194 -9900
rect 15234 -9934 15268 -9900
rect 15308 -9934 15342 -9900
rect 15382 -9934 15416 -9900
rect 15456 -9934 15490 -9900
rect 15530 -9934 15564 -9900
rect 15604 -9934 15638 -9900
rect 15678 -9934 15712 -9900
rect 15752 -9934 15786 -9900
rect 15826 -9934 15860 -9900
rect 15900 -9934 15934 -9900
rect 15974 -9934 16008 -9900
rect 16048 -9934 16082 -9900
rect 16122 -9934 16156 -9900
rect 16196 -9934 16230 -9900
rect 16270 -9934 16304 -9900
rect 16344 -9934 16378 -9900
rect 16418 -9934 16452 -9900
rect 16492 -9934 16526 -9900
rect 16566 -9934 16600 -9900
rect 16640 -9934 16674 -9900
rect 16714 -9934 16748 -9900
rect 16788 -9934 16822 -9900
rect 16862 -9934 16896 -9900
rect 16936 -9934 16970 -9900
rect 17010 -9934 17044 -9900
rect 17084 -9934 17118 -9900
rect 17158 -9934 17192 -9900
rect 17232 -9934 17266 -9900
rect 17306 -9934 17340 -9900
rect 17380 -9934 17414 -9900
rect 17454 -9934 17488 -9900
rect 17528 -9934 17562 -9900
rect 17602 -9934 17636 -9900
rect 17676 -9934 17710 -9900
rect 17750 -9934 17784 -9900
rect 17824 -9934 17858 -9900
rect 17898 -9934 17932 -9900
rect 17972 -9934 18006 -9900
rect 18046 -9934 18080 -9900
rect 18120 -9934 18154 -9900
rect 18194 -9934 18228 -9900
rect 18268 -9934 18302 -9900
rect 18342 -9934 18376 -9900
rect 18416 -9934 18450 -9900
rect 18490 -9934 18524 -9900
rect 18564 -9934 18598 -9900
rect 18638 -9934 18672 -9900
rect 18712 -9934 18746 -9900
rect 18786 -9934 18820 -9900
rect 18860 -9934 18894 -9900
rect 18934 -9934 18968 -9900
rect 19008 -9934 19042 -9900
rect 19082 -9934 19116 -9900
rect 19156 -9934 19190 -9900
rect 19230 -9934 19264 -9900
rect 19304 -9934 19338 -9900
rect 19378 -9934 19412 -9900
rect 19452 -9934 19486 -9900
rect 19526 -9934 19560 -9900
rect 19600 -9934 19634 -9900
rect 19674 -9934 19708 -9900
rect 19748 -9934 19782 -9900
rect 19822 -9934 19856 -9900
rect 19896 -9934 19930 -9900
rect 19970 -9934 20004 -9900
rect 20044 -9934 20078 -9900
rect 20118 -9934 20152 -9900
rect 20192 -9934 20226 -9900
rect 20266 -9934 20300 -9900
rect 20340 -9934 20374 -9900
rect 20414 -9934 20448 -9900
rect 20488 -9934 20522 -9900
rect 20562 -9934 20596 -9900
rect 20636 -9934 20670 -9900
rect 20710 -9934 20744 -9900
rect 20784 -9934 20818 -9900
rect 20858 -9934 20892 -9900
rect 20932 -9934 20966 -9900
rect 21006 -9934 21040 -9900
rect 21080 -9934 21114 -9900
rect 21154 -9934 21188 -9900
rect 21228 -9934 21262 -9900
rect 21302 -9934 21336 -9900
rect 21376 -9934 21410 -9900
rect 21450 -9934 21484 -9900
rect 21524 -9934 21558 -9900
rect 21598 -9934 21632 -9900
rect 21672 -9934 21706 -9900
rect 21746 -9934 21780 -9900
rect 21820 -9934 21854 -9900
rect 21894 -9934 21928 -9900
rect 21968 -9934 22002 -9900
rect 22042 -9934 22076 -9900
rect 22116 -9934 22150 -9900
rect 22190 -9934 22224 -9900
rect 22264 -9934 22298 -9900
rect 22338 -9934 22372 -9900
rect 22412 -9934 22446 -9900
rect 22486 -9934 22520 -9900
rect 22560 -9934 22594 -9900
rect 22634 -9934 22668 -9900
rect 22708 -9934 22742 -9900
rect 22782 -9934 22816 -9900
rect 22856 -9934 22890 -9900
rect 22930 -9934 22964 -9900
rect 23004 -9934 23038 -9900
rect 23078 -9934 23112 -9900
rect 23152 -9934 23186 -9900
rect 23226 -9934 23260 -9900
rect 23300 -9934 23334 -9900
rect 23374 -9934 23408 -9900
rect 23448 -9934 23482 -9900
rect 23522 -9934 23556 -9900
rect 23596 -9934 23630 -9900
rect 23670 -9934 23704 -9900
rect 23744 -9934 23778 -9900
rect 23818 -9934 23852 -9900
rect 23892 -9934 23926 -9900
rect 23966 -9934 24000 -9900
rect 24040 -9934 24074 -9900
rect 24114 -9934 24148 -9900
rect 24188 -9934 24222 -9900
rect 24262 -9934 24296 -9900
rect 24336 -9934 24370 -9900
rect 24410 -9934 24444 -9900
rect 24484 -9934 24518 -9900
rect 24558 -9934 24592 -9900
rect 24632 -9934 24666 -9900
rect 24706 -9934 24740 -9900
rect 24780 -9934 24814 -9900
rect 24854 -9934 24888 -9900
rect 24928 -9934 24962 -9900
rect 25002 -9934 25036 -9900
rect 25076 -9934 25110 -9900
rect 25150 -9934 25184 -9900
<< nsubdiffcont >>
rect 4792 3118 10762 3152
rect 12482 3117 18452 3151
rect 18621 3117 24591 3151
rect 4792 3030 10762 3064
rect 12482 3029 18452 3063
rect 18621 3029 24591 3063
rect 4792 2942 10762 2976
rect 12482 2941 18452 2975
rect 18621 2941 24591 2975
rect 4792 1427 10762 1461
rect 4792 1339 10762 1373
rect 4696 -333 4730 1277
rect 10824 -333 10858 1277
rect 4792 -429 10762 -395
rect 4792 -517 10762 -483
rect 4792 -605 10762 -571
rect 4792 -711 10762 -677
rect 4696 -2383 4730 -773
rect 10824 -2383 10858 -773
rect 4792 -2479 10762 -2445
rect 4792 -2567 10762 -2533
rect 4792 -2655 10762 -2621
rect 4792 -2761 10762 -2727
rect 4696 -4433 4730 -2823
rect 10824 -4433 10858 -2823
rect 4792 -4529 10762 -4495
rect 4792 -4617 10762 -4583
rect 4792 -4705 10762 -4671
rect 4792 -6667 10762 -6633
rect 4792 -6755 10762 -6721
<< poly >>
rect 7795 2040 7861 2054
rect 7795 2006 7811 2040
rect 7845 2006 7861 2040
rect 7795 1990 7861 2006
rect 7913 2040 7979 2054
rect 7913 2006 7929 2040
rect 7963 2006 7979 2040
rect 7913 1990 7979 2006
rect 8031 2040 8097 2054
rect 8031 2006 8047 2040
rect 8081 2006 8097 2040
rect 8031 1990 8097 2006
rect 8149 2040 8215 2054
rect 8149 2006 8165 2040
rect 8199 2006 8215 2040
rect 8149 1990 8215 2006
rect 8267 2040 8333 2054
rect 8267 2006 8283 2040
rect 8317 2006 8333 2040
rect 8267 1990 8333 2006
rect 8385 2040 8451 2054
rect 8385 2006 8401 2040
rect 8435 2006 8451 2040
rect 8385 1990 8451 2006
rect 8503 2040 8569 2054
rect 8503 2006 8519 2040
rect 8553 2006 8569 2040
rect 8503 1990 8569 2006
rect 8849 2040 8915 2054
rect 8849 2006 8865 2040
rect 8899 2006 8915 2040
rect 8849 1990 8915 2006
rect 8967 2040 9033 2054
rect 8967 2006 8983 2040
rect 9017 2006 9033 2040
rect 8967 1990 9033 2006
rect 9085 2040 9151 2054
rect 9085 2006 9101 2040
rect 9135 2006 9151 2040
rect 9085 1990 9151 2006
rect 9203 2040 9269 2054
rect 9203 2006 9219 2040
rect 9253 2006 9269 2040
rect 9203 1990 9269 2006
rect 9321 2040 9387 2054
rect 9321 2006 9337 2040
rect 9371 2006 9387 2040
rect 9321 1990 9387 2006
rect 9439 2040 9505 2054
rect 9439 2006 9455 2040
rect 9489 2006 9505 2040
rect 9439 1990 9505 2006
rect 9557 2040 9623 2054
rect 9557 2006 9573 2040
rect 9607 2006 9623 2040
rect 9557 1990 9623 2006
rect 9675 2040 9741 2054
rect 9675 2006 9691 2040
rect 9725 2006 9741 2040
rect 9675 1990 9741 2006
rect 9793 2040 9859 2054
rect 9793 2006 9809 2040
rect 9843 2006 9859 2040
rect 9793 1990 9859 2006
rect 9911 2040 9977 2054
rect 9911 2006 9927 2040
rect 9961 2006 9977 2040
rect 9911 1990 9977 2006
rect 10029 2040 10095 2054
rect 10029 2006 10045 2040
rect 10079 2006 10095 2040
rect 10029 1990 10095 2006
rect 10147 2040 10213 2054
rect 10147 2006 10163 2040
rect 10197 2006 10213 2040
rect 10147 1990 10213 2006
rect 10265 2040 10331 2054
rect 10265 2006 10281 2040
rect 10315 2006 10331 2040
rect 10265 1990 10331 2006
rect 10383 2040 10449 2054
rect 10383 2006 10399 2040
rect 10433 2006 10449 2040
rect 10383 1990 10449 2006
rect 10501 2040 10567 2054
rect 10501 2006 10517 2040
rect 10551 2006 10567 2040
rect 10501 1990 10567 2006
rect 12665 2039 12723 2045
rect 12665 2005 12677 2039
rect 12711 2005 12723 2039
rect 12665 1989 12723 2005
rect 12779 2039 12845 2055
rect 12779 2005 12795 2039
rect 12829 2005 12845 2039
rect 12779 1989 12845 2005
rect 12897 2039 12963 2055
rect 12897 2005 12913 2039
rect 12947 2005 12963 2039
rect 12897 1989 12963 2005
rect 13015 2039 13081 2055
rect 13015 2005 13031 2039
rect 13065 2005 13081 2039
rect 13015 1989 13081 2005
rect 13133 2039 13199 2055
rect 13133 2005 13149 2039
rect 13183 2005 13199 2039
rect 13133 1989 13199 2005
rect 13251 2039 13317 2055
rect 13251 2005 13267 2039
rect 13301 2005 13317 2039
rect 13251 1989 13317 2005
rect 13369 2039 13435 2055
rect 13369 2005 13385 2039
rect 13419 2005 13435 2039
rect 13369 1989 13435 2005
rect 13487 2039 13553 2055
rect 13487 2005 13503 2039
rect 13537 2005 13553 2039
rect 13487 1989 13553 2005
rect 13605 2039 13671 2055
rect 13605 2005 13621 2039
rect 13655 2005 13671 2039
rect 13605 1989 13671 2005
rect 13723 2039 13789 2055
rect 13723 2005 13739 2039
rect 13773 2005 13789 2039
rect 13723 1989 13789 2005
rect 13841 2039 13907 2055
rect 13841 2005 13857 2039
rect 13891 2005 13907 2039
rect 13841 1989 13907 2005
rect 13959 2039 14025 2055
rect 13959 2005 13975 2039
rect 14009 2005 14025 2039
rect 13959 1989 14025 2005
rect 14077 2039 14143 2055
rect 14077 2005 14093 2039
rect 14127 2005 14143 2039
rect 14077 1989 14143 2005
rect 14195 2039 14261 2055
rect 14195 2005 14211 2039
rect 14245 2005 14261 2039
rect 14195 1989 14261 2005
rect 14313 2039 14379 2055
rect 14313 2005 14329 2039
rect 14363 2005 14379 2039
rect 14313 1989 14379 2005
rect 14431 2039 14497 2055
rect 14431 2005 14447 2039
rect 14481 2005 14497 2039
rect 14431 1989 14497 2005
rect 14549 2039 14615 2055
rect 14549 2005 14565 2039
rect 14599 2005 14615 2039
rect 14549 1989 14615 2005
rect 14667 2039 14733 2055
rect 14667 2005 14683 2039
rect 14717 2005 14733 2039
rect 14667 1989 14733 2005
rect 14785 2039 14851 2055
rect 14785 2005 14801 2039
rect 14835 2005 14851 2039
rect 14785 1989 14851 2005
rect 14903 2039 14969 2055
rect 14903 2005 14919 2039
rect 14953 2005 14969 2039
rect 14903 1989 14969 2005
rect 15021 2039 15087 2055
rect 15021 2005 15037 2039
rect 15071 2005 15087 2039
rect 15021 1989 15087 2005
rect 15139 2039 15205 2055
rect 15139 2005 15155 2039
rect 15189 2005 15205 2039
rect 15139 1989 15205 2005
rect 15257 2039 15323 2055
rect 15257 2005 15273 2039
rect 15307 2005 15323 2039
rect 15257 1989 15323 2005
rect 15375 2039 15441 2055
rect 15375 2005 15391 2039
rect 15425 2005 15441 2039
rect 15375 1989 15441 2005
rect 16788 2039 16846 2045
rect 16788 2005 16800 2039
rect 16834 2005 16846 2039
rect 16788 1989 16846 2005
rect 16902 2039 16968 2055
rect 16902 2005 16918 2039
rect 16952 2005 16968 2039
rect 16902 1989 16968 2005
rect 17020 2039 17086 2055
rect 17020 2005 17036 2039
rect 17070 2005 17086 2039
rect 17020 1989 17086 2005
rect 17138 2039 17204 2055
rect 17138 2005 17154 2039
rect 17188 2005 17204 2039
rect 17138 1989 17204 2005
rect 17256 2039 17322 2055
rect 17256 2005 17272 2039
rect 17306 2005 17322 2039
rect 17256 1989 17322 2005
rect 17374 2039 17440 2055
rect 17374 2005 17390 2039
rect 17424 2005 17440 2039
rect 17374 1989 17440 2005
rect 17492 2039 17558 2055
rect 17492 2005 17508 2039
rect 17542 2005 17558 2039
rect 17492 1989 17558 2005
rect 17610 2039 17676 2055
rect 17610 2005 17626 2039
rect 17660 2005 17676 2039
rect 17610 1989 17676 2005
rect 17728 2039 17794 2055
rect 17728 2005 17744 2039
rect 17778 2005 17794 2039
rect 17728 1989 17794 2005
rect 17846 2039 17912 2055
rect 17846 2005 17862 2039
rect 17896 2005 17912 2039
rect 17846 1989 17912 2005
rect 17964 2039 18030 2055
rect 17964 2005 17980 2039
rect 18014 2005 18030 2039
rect 17964 1989 18030 2005
rect 18082 2039 18148 2055
rect 18082 2005 18098 2039
rect 18132 2005 18148 2039
rect 18082 1989 18148 2005
rect 18200 2039 18266 2055
rect 18200 2005 18216 2039
rect 18250 2005 18266 2039
rect 18200 1989 18266 2005
rect 18318 2039 18384 2055
rect 18318 2005 18334 2039
rect 18368 2005 18384 2039
rect 18318 1989 18384 2005
rect 18436 2039 18502 2055
rect 18436 2005 18452 2039
rect 18486 2005 18502 2039
rect 18436 1989 18502 2005
rect 18554 2039 18620 2055
rect 18554 2005 18570 2039
rect 18604 2005 18620 2039
rect 18554 1989 18620 2005
rect 18672 2039 18738 2055
rect 18672 2005 18688 2039
rect 18722 2005 18738 2039
rect 18672 1989 18738 2005
rect 18790 2039 18856 2055
rect 18790 2005 18806 2039
rect 18840 2005 18856 2039
rect 18790 1989 18856 2005
rect 18908 2039 18974 2055
rect 18908 2005 18924 2039
rect 18958 2005 18974 2039
rect 18908 1989 18974 2005
rect 19026 2039 19092 2055
rect 19026 2005 19042 2039
rect 19076 2005 19092 2039
rect 19026 1989 19092 2005
rect 19144 2039 19210 2055
rect 19144 2005 19160 2039
rect 19194 2005 19210 2039
rect 19144 1989 19210 2005
rect 19262 2039 19328 2055
rect 19262 2005 19278 2039
rect 19312 2005 19328 2039
rect 19262 1989 19328 2005
rect 19380 2039 19446 2055
rect 19380 2005 19396 2039
rect 19430 2005 19446 2039
rect 19380 1989 19446 2005
rect 19498 2039 19564 2055
rect 19498 2005 19514 2039
rect 19548 2005 19564 2039
rect 19498 1989 19564 2005
rect 20911 2039 20969 2045
rect 20911 2005 20923 2039
rect 20957 2005 20969 2039
rect 20911 1989 20969 2005
rect 21025 2039 21091 2055
rect 21025 2005 21041 2039
rect 21075 2005 21091 2039
rect 21025 1989 21091 2005
rect 21143 2039 21209 2055
rect 21143 2005 21159 2039
rect 21193 2005 21209 2039
rect 21143 1989 21209 2005
rect 21261 2039 21327 2055
rect 21261 2005 21277 2039
rect 21311 2005 21327 2039
rect 21261 1989 21327 2005
rect 21379 2039 21445 2055
rect 21379 2005 21395 2039
rect 21429 2005 21445 2039
rect 21379 1989 21445 2005
rect 21497 2039 21563 2055
rect 21497 2005 21513 2039
rect 21547 2005 21563 2039
rect 21497 1989 21563 2005
rect 21615 2039 21681 2055
rect 21615 2005 21631 2039
rect 21665 2005 21681 2039
rect 21615 1989 21681 2005
rect 21733 2039 21799 2055
rect 21733 2005 21749 2039
rect 21783 2005 21799 2039
rect 21733 1989 21799 2005
rect 21851 2039 21917 2055
rect 21851 2005 21867 2039
rect 21901 2005 21917 2039
rect 21851 1989 21917 2005
rect 21969 2039 22035 2055
rect 21969 2005 21985 2039
rect 22019 2005 22035 2039
rect 21969 1989 22035 2005
rect 22087 2039 22153 2055
rect 22087 2005 22103 2039
rect 22137 2005 22153 2039
rect 22087 1989 22153 2005
rect 22205 2039 22271 2055
rect 22205 2005 22221 2039
rect 22255 2005 22271 2039
rect 22205 1989 22271 2005
rect 22323 2039 22389 2055
rect 22323 2005 22339 2039
rect 22373 2005 22389 2039
rect 22323 1989 22389 2005
rect 22441 2039 22507 2055
rect 22441 2005 22457 2039
rect 22491 2005 22507 2039
rect 22441 1989 22507 2005
rect 22559 2039 22625 2055
rect 22559 2005 22575 2039
rect 22609 2005 22625 2039
rect 22559 1989 22625 2005
rect 22677 2039 22743 2055
rect 22677 2005 22693 2039
rect 22727 2005 22743 2039
rect 22677 1989 22743 2005
rect 22795 2039 22861 2055
rect 22795 2005 22811 2039
rect 22845 2005 22861 2039
rect 22795 1989 22861 2005
rect 22913 2039 22979 2055
rect 22913 2005 22929 2039
rect 22963 2005 22979 2039
rect 22913 1989 22979 2005
rect 23031 2039 23097 2055
rect 23031 2005 23047 2039
rect 23081 2005 23097 2039
rect 23031 1989 23097 2005
rect 23149 2039 23215 2055
rect 23149 2005 23165 2039
rect 23199 2005 23215 2039
rect 23149 1989 23215 2005
rect 23267 2039 23333 2055
rect 23267 2005 23283 2039
rect 23317 2005 23333 2039
rect 23267 1989 23333 2005
rect 23385 2039 23451 2055
rect 23385 2005 23401 2039
rect 23435 2005 23451 2039
rect 23385 1989 23451 2005
rect 23503 2039 23569 2055
rect 23503 2005 23519 2039
rect 23553 2005 23569 2039
rect 23503 1989 23569 2005
rect 23621 2039 23687 2055
rect 23621 2005 23637 2039
rect 23671 2005 23687 2039
rect 23621 1989 23687 2005
rect 12665 1931 12723 1947
rect 12665 1897 12677 1931
rect 12711 1897 12723 1931
rect 12665 1891 12723 1897
rect 12779 1931 12845 1947
rect 12779 1897 12795 1931
rect 12829 1897 12845 1931
rect 12779 1881 12845 1897
rect 12897 1931 12963 1947
rect 12897 1897 12913 1931
rect 12947 1897 12963 1931
rect 12897 1881 12963 1897
rect 13015 1931 13081 1947
rect 13015 1897 13031 1931
rect 13065 1897 13081 1931
rect 13015 1881 13081 1897
rect 13133 1931 13199 1947
rect 13133 1897 13149 1931
rect 13183 1897 13199 1931
rect 13133 1881 13199 1897
rect 13251 1931 13317 1947
rect 13251 1897 13267 1931
rect 13301 1897 13317 1931
rect 13251 1881 13317 1897
rect 13369 1931 13435 1947
rect 13369 1897 13385 1931
rect 13419 1897 13435 1931
rect 13369 1881 13435 1897
rect 13487 1931 13553 1947
rect 13487 1897 13503 1931
rect 13537 1897 13553 1931
rect 13487 1881 13553 1897
rect 13605 1931 13671 1947
rect 13605 1897 13621 1931
rect 13655 1897 13671 1931
rect 13605 1881 13671 1897
rect 13723 1931 13789 1947
rect 13723 1897 13739 1931
rect 13773 1897 13789 1931
rect 13723 1881 13789 1897
rect 13841 1931 13907 1947
rect 13841 1897 13857 1931
rect 13891 1897 13907 1931
rect 13841 1881 13907 1897
rect 13959 1931 14025 1947
rect 13959 1897 13975 1931
rect 14009 1897 14025 1931
rect 13959 1881 14025 1897
rect 14077 1931 14143 1947
rect 14077 1897 14093 1931
rect 14127 1897 14143 1931
rect 14077 1881 14143 1897
rect 14195 1931 14261 1947
rect 14195 1897 14211 1931
rect 14245 1897 14261 1931
rect 14195 1881 14261 1897
rect 14313 1931 14379 1947
rect 14313 1897 14329 1931
rect 14363 1897 14379 1931
rect 14313 1881 14379 1897
rect 14431 1931 14497 1947
rect 14431 1897 14447 1931
rect 14481 1897 14497 1931
rect 14431 1881 14497 1897
rect 14549 1931 14615 1947
rect 14549 1897 14565 1931
rect 14599 1897 14615 1931
rect 14549 1881 14615 1897
rect 14667 1931 14733 1947
rect 14667 1897 14683 1931
rect 14717 1897 14733 1931
rect 14667 1881 14733 1897
rect 14785 1931 14851 1947
rect 14785 1897 14801 1931
rect 14835 1897 14851 1931
rect 14785 1881 14851 1897
rect 14903 1931 14969 1947
rect 14903 1897 14919 1931
rect 14953 1897 14969 1931
rect 14903 1881 14969 1897
rect 15021 1931 15087 1947
rect 15021 1897 15037 1931
rect 15071 1897 15087 1931
rect 15021 1881 15087 1897
rect 15139 1931 15205 1947
rect 15139 1897 15155 1931
rect 15189 1897 15205 1931
rect 15139 1881 15205 1897
rect 15257 1931 15323 1947
rect 15257 1897 15273 1931
rect 15307 1897 15323 1931
rect 15257 1881 15323 1897
rect 15375 1931 15441 1947
rect 15375 1897 15391 1931
rect 15425 1897 15441 1931
rect 15375 1881 15441 1897
rect 16788 1931 16846 1947
rect 16788 1897 16800 1931
rect 16834 1897 16846 1931
rect 16788 1891 16846 1897
rect 16902 1931 16968 1947
rect 16902 1897 16918 1931
rect 16952 1897 16968 1931
rect 16902 1881 16968 1897
rect 17020 1931 17086 1947
rect 17020 1897 17036 1931
rect 17070 1897 17086 1931
rect 17020 1881 17086 1897
rect 17138 1931 17204 1947
rect 17138 1897 17154 1931
rect 17188 1897 17204 1931
rect 17138 1881 17204 1897
rect 17256 1931 17322 1947
rect 17256 1897 17272 1931
rect 17306 1897 17322 1931
rect 17256 1881 17322 1897
rect 17374 1931 17440 1947
rect 17374 1897 17390 1931
rect 17424 1897 17440 1931
rect 17374 1881 17440 1897
rect 17492 1931 17558 1947
rect 17492 1897 17508 1931
rect 17542 1897 17558 1931
rect 17492 1881 17558 1897
rect 17610 1931 17676 1947
rect 17610 1897 17626 1931
rect 17660 1897 17676 1931
rect 17610 1881 17676 1897
rect 17728 1931 17794 1947
rect 17728 1897 17744 1931
rect 17778 1897 17794 1931
rect 17728 1881 17794 1897
rect 17846 1931 17912 1947
rect 17846 1897 17862 1931
rect 17896 1897 17912 1931
rect 17846 1881 17912 1897
rect 17964 1931 18030 1947
rect 17964 1897 17980 1931
rect 18014 1897 18030 1931
rect 17964 1881 18030 1897
rect 18082 1931 18148 1947
rect 18082 1897 18098 1931
rect 18132 1897 18148 1931
rect 18082 1881 18148 1897
rect 18200 1931 18266 1947
rect 18200 1897 18216 1931
rect 18250 1897 18266 1931
rect 18200 1881 18266 1897
rect 18318 1931 18384 1947
rect 18318 1897 18334 1931
rect 18368 1897 18384 1931
rect 18318 1881 18384 1897
rect 18436 1931 18502 1947
rect 18436 1897 18452 1931
rect 18486 1897 18502 1931
rect 18436 1881 18502 1897
rect 18554 1931 18620 1947
rect 18554 1897 18570 1931
rect 18604 1897 18620 1931
rect 18554 1881 18620 1897
rect 18672 1931 18738 1947
rect 18672 1897 18688 1931
rect 18722 1897 18738 1931
rect 18672 1881 18738 1897
rect 18790 1931 18856 1947
rect 18790 1897 18806 1931
rect 18840 1897 18856 1931
rect 18790 1881 18856 1897
rect 18908 1931 18974 1947
rect 18908 1897 18924 1931
rect 18958 1897 18974 1931
rect 18908 1881 18974 1897
rect 19026 1931 19092 1947
rect 19026 1897 19042 1931
rect 19076 1897 19092 1931
rect 19026 1881 19092 1897
rect 19144 1931 19210 1947
rect 19144 1897 19160 1931
rect 19194 1897 19210 1931
rect 19144 1881 19210 1897
rect 19262 1931 19328 1947
rect 19262 1897 19278 1931
rect 19312 1897 19328 1931
rect 19262 1881 19328 1897
rect 19380 1931 19446 1947
rect 19380 1897 19396 1931
rect 19430 1897 19446 1931
rect 19380 1881 19446 1897
rect 19498 1931 19564 1947
rect 19498 1897 19514 1931
rect 19548 1897 19564 1931
rect 19498 1881 19564 1897
rect 20911 1931 20969 1947
rect 20911 1897 20923 1931
rect 20957 1897 20969 1931
rect 20911 1891 20969 1897
rect 21025 1931 21091 1947
rect 21025 1897 21041 1931
rect 21075 1897 21091 1931
rect 21025 1881 21091 1897
rect 21143 1931 21209 1947
rect 21143 1897 21159 1931
rect 21193 1897 21209 1931
rect 21143 1881 21209 1897
rect 21261 1931 21327 1947
rect 21261 1897 21277 1931
rect 21311 1897 21327 1931
rect 21261 1881 21327 1897
rect 21379 1931 21445 1947
rect 21379 1897 21395 1931
rect 21429 1897 21445 1931
rect 21379 1881 21445 1897
rect 21497 1931 21563 1947
rect 21497 1897 21513 1931
rect 21547 1897 21563 1931
rect 21497 1881 21563 1897
rect 21615 1931 21681 1947
rect 21615 1897 21631 1931
rect 21665 1897 21681 1931
rect 21615 1881 21681 1897
rect 21733 1931 21799 1947
rect 21733 1897 21749 1931
rect 21783 1897 21799 1931
rect 21733 1881 21799 1897
rect 21851 1931 21917 1947
rect 21851 1897 21867 1931
rect 21901 1897 21917 1931
rect 21851 1881 21917 1897
rect 21969 1931 22035 1947
rect 21969 1897 21985 1931
rect 22019 1897 22035 1931
rect 21969 1881 22035 1897
rect 22087 1931 22153 1947
rect 22087 1897 22103 1931
rect 22137 1897 22153 1931
rect 22087 1881 22153 1897
rect 22205 1931 22271 1947
rect 22205 1897 22221 1931
rect 22255 1897 22271 1931
rect 22205 1881 22271 1897
rect 22323 1931 22389 1947
rect 22323 1897 22339 1931
rect 22373 1897 22389 1931
rect 22323 1881 22389 1897
rect 22441 1931 22507 1947
rect 22441 1897 22457 1931
rect 22491 1897 22507 1931
rect 22441 1881 22507 1897
rect 22559 1931 22625 1947
rect 22559 1897 22575 1931
rect 22609 1897 22625 1931
rect 22559 1881 22625 1897
rect 22677 1931 22743 1947
rect 22677 1897 22693 1931
rect 22727 1897 22743 1931
rect 22677 1881 22743 1897
rect 22795 1931 22861 1947
rect 22795 1897 22811 1931
rect 22845 1897 22861 1931
rect 22795 1881 22861 1897
rect 22913 1931 22979 1947
rect 22913 1897 22929 1931
rect 22963 1897 22979 1931
rect 22913 1881 22979 1897
rect 23031 1931 23097 1947
rect 23031 1897 23047 1931
rect 23081 1897 23097 1931
rect 23031 1881 23097 1897
rect 23149 1931 23215 1947
rect 23149 1897 23165 1931
rect 23199 1897 23215 1931
rect 23149 1881 23215 1897
rect 23267 1931 23333 1947
rect 23267 1897 23283 1931
rect 23317 1897 23333 1931
rect 23267 1881 23333 1897
rect 23385 1931 23451 1947
rect 23385 1897 23401 1931
rect 23435 1897 23451 1931
rect 23385 1881 23451 1897
rect 23503 1931 23569 1947
rect 23503 1897 23519 1931
rect 23553 1897 23569 1931
rect 23503 1881 23569 1897
rect 23621 1931 23687 1947
rect 23621 1897 23637 1931
rect 23671 1897 23687 1931
rect 23621 1881 23687 1897
rect 4853 1221 4919 1287
rect 4971 1221 5037 1287
rect 5089 1221 5155 1287
rect 5207 1221 5273 1287
rect 5325 1221 5391 1287
rect 5443 1221 5509 1287
rect 5561 1221 5627 1287
rect 5679 1221 5745 1287
rect 5797 1221 5863 1287
rect 5915 1221 5981 1287
rect 6033 1221 6099 1287
rect 6151 1221 6217 1287
rect 6269 1221 6335 1287
rect 6387 1221 6453 1287
rect 6505 1221 6571 1287
rect 6623 1221 6689 1287
rect 6741 1221 6807 1287
rect 6859 1221 6925 1287
rect 6977 1221 7043 1287
rect 7095 1221 7161 1287
rect 7213 1221 7279 1287
rect 7331 1221 7397 1287
rect 7449 1221 7515 1287
rect 7567 1221 7633 1287
rect 7685 1221 7751 1287
rect 7803 1221 7869 1287
rect 7921 1221 7987 1287
rect 8039 1221 8105 1287
rect 8157 1221 8223 1287
rect 8275 1221 8341 1287
rect 8393 1221 8459 1287
rect 8511 1221 8577 1287
rect 8629 1221 8695 1287
rect 8747 1221 8813 1287
rect 8865 1221 8931 1287
rect 8983 1221 9049 1287
rect 9101 1221 9167 1287
rect 9219 1221 9285 1287
rect 9337 1221 9403 1287
rect 9455 1221 9521 1287
rect 9573 1221 9639 1287
rect 9691 1221 9757 1287
rect 9809 1221 9875 1287
rect 9927 1221 9993 1287
rect 10045 1221 10111 1287
rect 10163 1221 10229 1287
rect 10281 1221 10347 1287
rect 10399 1221 10465 1287
rect 10517 1221 10583 1287
rect 10635 1221 10701 1287
rect 4856 1190 4916 1221
rect 4974 1190 5034 1221
rect 5092 1190 5152 1221
rect 5210 1190 5270 1221
rect 5328 1190 5388 1221
rect 5446 1190 5506 1221
rect 5564 1190 5624 1221
rect 5682 1190 5742 1221
rect 5800 1190 5860 1221
rect 5918 1190 5978 1221
rect 6036 1190 6096 1221
rect 6154 1190 6214 1221
rect 6272 1190 6332 1221
rect 6390 1190 6450 1221
rect 6508 1190 6568 1221
rect 6626 1190 6686 1221
rect 6744 1190 6804 1221
rect 6862 1190 6922 1221
rect 6980 1190 7040 1221
rect 7098 1190 7158 1221
rect 7216 1190 7276 1221
rect 7334 1190 7394 1221
rect 7452 1190 7512 1221
rect 7570 1190 7630 1221
rect 7688 1190 7748 1221
rect 7806 1190 7866 1221
rect 7924 1190 7984 1221
rect 8042 1190 8102 1221
rect 8160 1190 8220 1221
rect 8278 1190 8338 1221
rect 8396 1190 8456 1221
rect 8514 1190 8574 1221
rect 8632 1190 8692 1221
rect 8750 1190 8810 1221
rect 8868 1190 8928 1221
rect 8986 1190 9046 1221
rect 9104 1190 9164 1221
rect 9222 1190 9282 1221
rect 9340 1190 9400 1221
rect 9458 1190 9518 1221
rect 9576 1190 9636 1221
rect 9694 1190 9754 1221
rect 9812 1190 9872 1221
rect 9930 1190 9990 1221
rect 10048 1190 10108 1221
rect 10166 1190 10226 1221
rect 10284 1190 10344 1221
rect 10402 1190 10462 1221
rect 10520 1190 10580 1221
rect 10638 1190 10698 1221
rect 4856 559 4916 590
rect 4974 559 5034 590
rect 5092 559 5152 590
rect 5210 559 5270 590
rect 5328 559 5388 590
rect 5446 559 5506 590
rect 5564 559 5624 590
rect 5682 559 5742 590
rect 5800 559 5860 590
rect 5918 559 5978 590
rect 6036 559 6096 590
rect 6154 559 6214 590
rect 6272 559 6332 590
rect 6390 559 6450 590
rect 6508 559 6568 590
rect 6626 559 6686 590
rect 6744 559 6804 590
rect 6862 559 6922 590
rect 6980 559 7040 590
rect 7098 559 7158 590
rect 7216 559 7276 590
rect 7334 559 7394 590
rect 7452 559 7512 590
rect 7570 559 7630 590
rect 7688 559 7748 590
rect 7806 559 7866 590
rect 7924 559 7984 590
rect 8042 559 8102 590
rect 8160 559 8220 590
rect 8278 559 8338 590
rect 8396 559 8456 590
rect 8514 559 8574 590
rect 8632 559 8692 590
rect 8750 559 8810 590
rect 8868 559 8928 590
rect 8986 559 9046 590
rect 9104 559 9164 590
rect 9222 559 9282 590
rect 9340 559 9400 590
rect 9458 559 9518 590
rect 9576 559 9636 590
rect 9694 559 9754 590
rect 9812 559 9872 590
rect 9930 559 9990 590
rect 10048 559 10108 590
rect 10166 559 10226 590
rect 10284 559 10344 590
rect 10402 559 10462 590
rect 10520 559 10580 590
rect 10638 559 10698 590
rect 4853 543 4919 559
rect 4853 509 4869 543
rect 4903 509 4919 543
rect 4853 435 4919 509
rect 4853 401 4869 435
rect 4903 401 4919 435
rect 4853 385 4919 401
rect 4971 543 5037 559
rect 4971 509 4987 543
rect 5021 509 5037 543
rect 4971 435 5037 509
rect 4971 401 4987 435
rect 5021 401 5037 435
rect 4971 385 5037 401
rect 5089 543 5155 559
rect 5089 509 5105 543
rect 5139 509 5155 543
rect 5089 435 5155 509
rect 5089 401 5105 435
rect 5139 401 5155 435
rect 5089 385 5155 401
rect 5207 543 5273 559
rect 5207 509 5223 543
rect 5257 509 5273 543
rect 5207 435 5273 509
rect 5207 401 5223 435
rect 5257 401 5273 435
rect 5207 385 5273 401
rect 5325 543 5391 559
rect 5325 509 5341 543
rect 5375 509 5391 543
rect 5325 435 5391 509
rect 5325 401 5341 435
rect 5375 401 5391 435
rect 5325 385 5391 401
rect 5443 543 5509 559
rect 5443 509 5459 543
rect 5493 509 5509 543
rect 5443 435 5509 509
rect 5443 401 5459 435
rect 5493 401 5509 435
rect 5443 385 5509 401
rect 5561 543 5627 559
rect 5561 509 5577 543
rect 5611 509 5627 543
rect 5561 435 5627 509
rect 5561 401 5577 435
rect 5611 401 5627 435
rect 5561 385 5627 401
rect 5679 543 5745 559
rect 5679 509 5695 543
rect 5729 509 5745 543
rect 5679 435 5745 509
rect 5679 401 5695 435
rect 5729 401 5745 435
rect 5679 385 5745 401
rect 5797 543 5863 559
rect 5797 509 5813 543
rect 5847 509 5863 543
rect 5797 435 5863 509
rect 5797 401 5813 435
rect 5847 401 5863 435
rect 5797 385 5863 401
rect 5915 543 5981 559
rect 5915 509 5931 543
rect 5965 509 5981 543
rect 5915 435 5981 509
rect 5915 401 5931 435
rect 5965 401 5981 435
rect 5915 385 5981 401
rect 6033 543 6099 559
rect 6033 509 6049 543
rect 6083 509 6099 543
rect 6033 435 6099 509
rect 6033 401 6049 435
rect 6083 401 6099 435
rect 6033 385 6099 401
rect 6151 543 6217 559
rect 6151 509 6167 543
rect 6201 509 6217 543
rect 6151 435 6217 509
rect 6151 401 6167 435
rect 6201 401 6217 435
rect 6151 385 6217 401
rect 6269 543 6335 559
rect 6269 509 6285 543
rect 6319 509 6335 543
rect 6269 435 6335 509
rect 6269 401 6285 435
rect 6319 401 6335 435
rect 6269 385 6335 401
rect 6387 543 6453 559
rect 6387 509 6403 543
rect 6437 509 6453 543
rect 6387 435 6453 509
rect 6387 401 6403 435
rect 6437 401 6453 435
rect 6387 385 6453 401
rect 6505 543 6571 559
rect 6505 509 6521 543
rect 6555 509 6571 543
rect 6505 435 6571 509
rect 6505 401 6521 435
rect 6555 401 6571 435
rect 6505 385 6571 401
rect 6623 543 6689 559
rect 6623 509 6639 543
rect 6673 509 6689 543
rect 6623 435 6689 509
rect 6623 401 6639 435
rect 6673 401 6689 435
rect 6623 385 6689 401
rect 6741 543 6807 559
rect 6741 509 6757 543
rect 6791 509 6807 543
rect 6741 435 6807 509
rect 6741 401 6757 435
rect 6791 401 6807 435
rect 6741 385 6807 401
rect 6859 543 6925 559
rect 6859 509 6875 543
rect 6909 509 6925 543
rect 6859 435 6925 509
rect 6859 401 6875 435
rect 6909 401 6925 435
rect 6859 385 6925 401
rect 6977 543 7043 559
rect 6977 509 6993 543
rect 7027 509 7043 543
rect 6977 435 7043 509
rect 6977 401 6993 435
rect 7027 401 7043 435
rect 6977 385 7043 401
rect 7095 543 7161 559
rect 7095 509 7111 543
rect 7145 509 7161 543
rect 7095 435 7161 509
rect 7095 401 7111 435
rect 7145 401 7161 435
rect 7095 385 7161 401
rect 7213 543 7279 559
rect 7213 509 7229 543
rect 7263 509 7279 543
rect 7213 435 7279 509
rect 7213 401 7229 435
rect 7263 401 7279 435
rect 7213 385 7279 401
rect 7331 543 7397 559
rect 7331 509 7347 543
rect 7381 509 7397 543
rect 7331 435 7397 509
rect 7331 401 7347 435
rect 7381 401 7397 435
rect 7331 385 7397 401
rect 7449 543 7515 559
rect 7449 509 7465 543
rect 7499 509 7515 543
rect 7449 435 7515 509
rect 7449 401 7465 435
rect 7499 401 7515 435
rect 7449 385 7515 401
rect 7567 543 7633 559
rect 7567 509 7583 543
rect 7617 509 7633 543
rect 7567 435 7633 509
rect 7567 401 7583 435
rect 7617 401 7633 435
rect 7567 385 7633 401
rect 7685 543 7751 559
rect 7685 509 7701 543
rect 7735 509 7751 543
rect 7685 435 7751 509
rect 7685 401 7701 435
rect 7735 401 7751 435
rect 7685 385 7751 401
rect 7803 543 7869 559
rect 7803 509 7819 543
rect 7853 509 7869 543
rect 7803 435 7869 509
rect 7803 401 7819 435
rect 7853 401 7869 435
rect 7803 385 7869 401
rect 7921 543 7987 559
rect 7921 509 7937 543
rect 7971 509 7987 543
rect 7921 435 7987 509
rect 7921 401 7937 435
rect 7971 401 7987 435
rect 7921 385 7987 401
rect 8039 543 8105 559
rect 8039 509 8055 543
rect 8089 509 8105 543
rect 8039 435 8105 509
rect 8039 401 8055 435
rect 8089 401 8105 435
rect 8039 385 8105 401
rect 8157 543 8223 559
rect 8157 509 8173 543
rect 8207 509 8223 543
rect 8157 435 8223 509
rect 8157 401 8173 435
rect 8207 401 8223 435
rect 8157 385 8223 401
rect 8275 543 8341 559
rect 8275 509 8291 543
rect 8325 509 8341 543
rect 8275 435 8341 509
rect 8275 401 8291 435
rect 8325 401 8341 435
rect 8275 385 8341 401
rect 8393 543 8459 559
rect 8393 509 8409 543
rect 8443 509 8459 543
rect 8393 435 8459 509
rect 8393 401 8409 435
rect 8443 401 8459 435
rect 8393 385 8459 401
rect 8511 543 8577 559
rect 8511 509 8527 543
rect 8561 509 8577 543
rect 8511 435 8577 509
rect 8511 401 8527 435
rect 8561 401 8577 435
rect 8511 385 8577 401
rect 8629 543 8695 559
rect 8629 509 8645 543
rect 8679 509 8695 543
rect 8629 435 8695 509
rect 8629 401 8645 435
rect 8679 401 8695 435
rect 8629 385 8695 401
rect 8747 543 8813 559
rect 8747 509 8763 543
rect 8797 509 8813 543
rect 8747 435 8813 509
rect 8747 401 8763 435
rect 8797 401 8813 435
rect 8747 385 8813 401
rect 8865 543 8931 559
rect 8865 509 8881 543
rect 8915 509 8931 543
rect 8865 435 8931 509
rect 8865 401 8881 435
rect 8915 401 8931 435
rect 8865 385 8931 401
rect 8983 543 9049 559
rect 8983 509 8999 543
rect 9033 509 9049 543
rect 8983 435 9049 509
rect 8983 401 8999 435
rect 9033 401 9049 435
rect 8983 385 9049 401
rect 9101 543 9167 559
rect 9101 509 9117 543
rect 9151 509 9167 543
rect 9101 435 9167 509
rect 9101 401 9117 435
rect 9151 401 9167 435
rect 9101 385 9167 401
rect 9219 543 9285 559
rect 9219 509 9235 543
rect 9269 509 9285 543
rect 9219 435 9285 509
rect 9219 401 9235 435
rect 9269 401 9285 435
rect 9219 385 9285 401
rect 9337 543 9403 559
rect 9337 509 9353 543
rect 9387 509 9403 543
rect 9337 435 9403 509
rect 9337 401 9353 435
rect 9387 401 9403 435
rect 9337 385 9403 401
rect 9455 543 9521 559
rect 9455 509 9471 543
rect 9505 509 9521 543
rect 9455 435 9521 509
rect 9455 401 9471 435
rect 9505 401 9521 435
rect 9455 385 9521 401
rect 9573 543 9639 559
rect 9573 509 9589 543
rect 9623 509 9639 543
rect 9573 435 9639 509
rect 9573 401 9589 435
rect 9623 401 9639 435
rect 9573 385 9639 401
rect 9691 543 9757 559
rect 9691 509 9707 543
rect 9741 509 9757 543
rect 9691 435 9757 509
rect 9691 401 9707 435
rect 9741 401 9757 435
rect 9691 385 9757 401
rect 9809 543 9875 559
rect 9809 509 9825 543
rect 9859 509 9875 543
rect 9809 435 9875 509
rect 9809 401 9825 435
rect 9859 401 9875 435
rect 9809 385 9875 401
rect 9927 543 9993 559
rect 9927 509 9943 543
rect 9977 509 9993 543
rect 9927 435 9993 509
rect 9927 401 9943 435
rect 9977 401 9993 435
rect 9927 385 9993 401
rect 10045 543 10111 559
rect 10045 509 10061 543
rect 10095 509 10111 543
rect 10045 435 10111 509
rect 10045 401 10061 435
rect 10095 401 10111 435
rect 10045 385 10111 401
rect 10163 543 10229 559
rect 10163 509 10179 543
rect 10213 509 10229 543
rect 10163 435 10229 509
rect 10163 401 10179 435
rect 10213 401 10229 435
rect 10163 385 10229 401
rect 10281 543 10347 559
rect 10281 509 10297 543
rect 10331 509 10347 543
rect 10281 435 10347 509
rect 10281 401 10297 435
rect 10331 401 10347 435
rect 10281 385 10347 401
rect 10399 543 10465 559
rect 10399 509 10415 543
rect 10449 509 10465 543
rect 10399 435 10465 509
rect 10399 401 10415 435
rect 10449 401 10465 435
rect 10399 385 10465 401
rect 10517 543 10583 559
rect 10517 509 10533 543
rect 10567 509 10583 543
rect 10517 435 10583 509
rect 10517 401 10533 435
rect 10567 401 10583 435
rect 10517 385 10583 401
rect 10635 543 10701 559
rect 10635 509 10651 543
rect 10685 509 10701 543
rect 10635 435 10701 509
rect 10635 401 10651 435
rect 10685 401 10701 435
rect 10635 385 10701 401
rect 4856 354 4916 385
rect 4974 354 5034 385
rect 5092 354 5152 385
rect 5210 354 5270 385
rect 5328 354 5388 385
rect 5446 354 5506 385
rect 5564 354 5624 385
rect 5682 354 5742 385
rect 5800 354 5860 385
rect 5918 354 5978 385
rect 6036 354 6096 385
rect 6154 354 6214 385
rect 6272 354 6332 385
rect 6390 354 6450 385
rect 6508 354 6568 385
rect 6626 354 6686 385
rect 6744 354 6804 385
rect 6862 354 6922 385
rect 6980 354 7040 385
rect 7098 354 7158 385
rect 7216 354 7276 385
rect 7334 354 7394 385
rect 7452 354 7512 385
rect 7570 354 7630 385
rect 7688 354 7748 385
rect 7806 354 7866 385
rect 7924 354 7984 385
rect 8042 354 8102 385
rect 8160 354 8220 385
rect 8278 354 8338 385
rect 8396 354 8456 385
rect 8514 354 8574 385
rect 8632 354 8692 385
rect 8750 354 8810 385
rect 8868 354 8928 385
rect 8986 354 9046 385
rect 9104 354 9164 385
rect 9222 354 9282 385
rect 9340 354 9400 385
rect 9458 354 9518 385
rect 9576 354 9636 385
rect 9694 354 9754 385
rect 9812 354 9872 385
rect 9930 354 9990 385
rect 10048 354 10108 385
rect 10166 354 10226 385
rect 10284 354 10344 385
rect 10402 354 10462 385
rect 10520 354 10580 385
rect 10638 354 10698 385
rect 4856 -277 4916 -246
rect 4974 -277 5034 -246
rect 5092 -277 5152 -246
rect 5210 -277 5270 -246
rect 5328 -277 5388 -246
rect 5446 -277 5506 -246
rect 5564 -277 5624 -246
rect 5682 -277 5742 -246
rect 5800 -277 5860 -246
rect 5918 -277 5978 -246
rect 6036 -277 6096 -246
rect 6154 -277 6214 -246
rect 6272 -277 6332 -246
rect 6390 -277 6450 -246
rect 6508 -277 6568 -246
rect 6626 -277 6686 -246
rect 6744 -277 6804 -246
rect 6862 -277 6922 -246
rect 6980 -277 7040 -246
rect 7098 -277 7158 -246
rect 7216 -277 7276 -246
rect 7334 -277 7394 -246
rect 7452 -277 7512 -246
rect 7570 -277 7630 -246
rect 7688 -277 7748 -246
rect 7806 -277 7866 -246
rect 7924 -277 7984 -246
rect 8042 -277 8102 -246
rect 8160 -277 8220 -246
rect 8278 -277 8338 -246
rect 8396 -277 8456 -246
rect 8514 -277 8574 -246
rect 8632 -277 8692 -246
rect 8750 -277 8810 -246
rect 8868 -277 8928 -246
rect 8986 -277 9046 -246
rect 9104 -277 9164 -246
rect 9222 -277 9282 -246
rect 9340 -277 9400 -246
rect 9458 -277 9518 -246
rect 9576 -277 9636 -246
rect 9694 -277 9754 -246
rect 9812 -277 9872 -246
rect 9930 -277 9990 -246
rect 10048 -277 10108 -246
rect 10166 -277 10226 -246
rect 10284 -277 10344 -246
rect 10402 -277 10462 -246
rect 10520 -277 10580 -246
rect 10638 -277 10698 -246
rect 4853 -343 4919 -277
rect 4971 -343 5037 -277
rect 5089 -343 5155 -277
rect 5207 -343 5273 -277
rect 5325 -343 5391 -277
rect 5443 -343 5509 -277
rect 5561 -343 5627 -277
rect 5679 -343 5745 -277
rect 5797 -343 5863 -277
rect 5915 -343 5981 -277
rect 6033 -343 6099 -277
rect 6151 -343 6217 -277
rect 6269 -343 6335 -277
rect 6387 -343 6453 -277
rect 6505 -343 6571 -277
rect 6623 -343 6689 -277
rect 6741 -343 6807 -277
rect 6859 -343 6925 -277
rect 6977 -343 7043 -277
rect 7095 -343 7161 -277
rect 7213 -343 7279 -277
rect 7331 -343 7397 -277
rect 7449 -343 7515 -277
rect 7567 -343 7633 -277
rect 7685 -343 7751 -277
rect 7803 -343 7869 -277
rect 7921 -343 7987 -277
rect 8039 -343 8105 -277
rect 8157 -343 8223 -277
rect 8275 -343 8341 -277
rect 8393 -343 8459 -277
rect 8511 -343 8577 -277
rect 8629 -343 8695 -277
rect 8747 -343 8813 -277
rect 8865 -343 8931 -277
rect 8983 -343 9049 -277
rect 9101 -343 9167 -277
rect 9219 -343 9285 -277
rect 9337 -343 9403 -277
rect 9455 -343 9521 -277
rect 9573 -343 9639 -277
rect 9691 -343 9757 -277
rect 9809 -343 9875 -277
rect 9927 -343 9993 -277
rect 10045 -343 10111 -277
rect 10163 -343 10229 -277
rect 10281 -343 10347 -277
rect 10399 -343 10465 -277
rect 10517 -343 10583 -277
rect 10635 -343 10701 -277
rect 4853 -829 4919 -763
rect 4971 -829 5037 -763
rect 5089 -829 5155 -763
rect 5207 -829 5273 -763
rect 5325 -829 5391 -763
rect 5443 -829 5509 -763
rect 5561 -829 5627 -763
rect 5679 -829 5745 -763
rect 5797 -829 5863 -763
rect 5915 -829 5981 -763
rect 6033 -829 6099 -763
rect 6151 -829 6217 -763
rect 6269 -829 6335 -763
rect 6387 -829 6453 -763
rect 6505 -829 6571 -763
rect 6623 -829 6689 -763
rect 6741 -829 6807 -763
rect 6859 -829 6925 -763
rect 6977 -829 7043 -763
rect 7095 -829 7161 -763
rect 7213 -829 7279 -763
rect 7331 -829 7397 -763
rect 7449 -829 7515 -763
rect 7567 -829 7633 -763
rect 7685 -829 7751 -763
rect 7803 -829 7869 -763
rect 7921 -829 7987 -763
rect 8039 -829 8105 -763
rect 8157 -829 8223 -763
rect 8275 -829 8341 -763
rect 8393 -829 8459 -763
rect 8511 -829 8577 -763
rect 8629 -829 8695 -763
rect 8747 -829 8813 -763
rect 8865 -829 8931 -763
rect 8983 -829 9049 -763
rect 9101 -829 9167 -763
rect 9219 -829 9285 -763
rect 9337 -829 9403 -763
rect 9455 -829 9521 -763
rect 9573 -829 9639 -763
rect 9691 -829 9757 -763
rect 9809 -829 9875 -763
rect 9927 -829 9993 -763
rect 10045 -829 10111 -763
rect 10163 -829 10229 -763
rect 10281 -829 10347 -763
rect 10399 -829 10465 -763
rect 10517 -829 10583 -763
rect 10635 -829 10701 -763
rect 4856 -860 4916 -829
rect 4974 -860 5034 -829
rect 5092 -860 5152 -829
rect 5210 -860 5270 -829
rect 5328 -860 5388 -829
rect 5446 -860 5506 -829
rect 5564 -860 5624 -829
rect 5682 -860 5742 -829
rect 5800 -860 5860 -829
rect 5918 -860 5978 -829
rect 6036 -860 6096 -829
rect 6154 -860 6214 -829
rect 6272 -860 6332 -829
rect 6390 -860 6450 -829
rect 6508 -860 6568 -829
rect 6626 -860 6686 -829
rect 6744 -860 6804 -829
rect 6862 -860 6922 -829
rect 6980 -860 7040 -829
rect 7098 -860 7158 -829
rect 7216 -860 7276 -829
rect 7334 -860 7394 -829
rect 7452 -860 7512 -829
rect 7570 -860 7630 -829
rect 7688 -860 7748 -829
rect 7806 -860 7866 -829
rect 7924 -860 7984 -829
rect 8042 -860 8102 -829
rect 8160 -860 8220 -829
rect 8278 -860 8338 -829
rect 8396 -860 8456 -829
rect 8514 -860 8574 -829
rect 8632 -860 8692 -829
rect 8750 -860 8810 -829
rect 8868 -860 8928 -829
rect 8986 -860 9046 -829
rect 9104 -860 9164 -829
rect 9222 -860 9282 -829
rect 9340 -860 9400 -829
rect 9458 -860 9518 -829
rect 9576 -860 9636 -829
rect 9694 -860 9754 -829
rect 9812 -860 9872 -829
rect 9930 -860 9990 -829
rect 10048 -860 10108 -829
rect 10166 -860 10226 -829
rect 10284 -860 10344 -829
rect 10402 -860 10462 -829
rect 10520 -860 10580 -829
rect 10638 -860 10698 -829
rect 4856 -1491 4916 -1460
rect 4974 -1491 5034 -1460
rect 5092 -1491 5152 -1460
rect 5210 -1491 5270 -1460
rect 5328 -1491 5388 -1460
rect 5446 -1491 5506 -1460
rect 5564 -1491 5624 -1460
rect 5682 -1491 5742 -1460
rect 5800 -1491 5860 -1460
rect 5918 -1491 5978 -1460
rect 6036 -1491 6096 -1460
rect 6154 -1491 6214 -1460
rect 6272 -1491 6332 -1460
rect 6390 -1491 6450 -1460
rect 6508 -1491 6568 -1460
rect 6626 -1491 6686 -1460
rect 6744 -1491 6804 -1460
rect 6862 -1491 6922 -1460
rect 6980 -1491 7040 -1460
rect 7098 -1491 7158 -1460
rect 7216 -1491 7276 -1460
rect 7334 -1491 7394 -1460
rect 7452 -1491 7512 -1460
rect 7570 -1491 7630 -1460
rect 7688 -1491 7748 -1460
rect 7806 -1491 7866 -1460
rect 7924 -1491 7984 -1460
rect 8042 -1491 8102 -1460
rect 8160 -1491 8220 -1460
rect 8278 -1491 8338 -1460
rect 8396 -1491 8456 -1460
rect 8514 -1491 8574 -1460
rect 8632 -1491 8692 -1460
rect 8750 -1491 8810 -1460
rect 8868 -1491 8928 -1460
rect 8986 -1491 9046 -1460
rect 9104 -1491 9164 -1460
rect 9222 -1491 9282 -1460
rect 9340 -1491 9400 -1460
rect 9458 -1491 9518 -1460
rect 9576 -1491 9636 -1460
rect 9694 -1491 9754 -1460
rect 9812 -1491 9872 -1460
rect 9930 -1491 9990 -1460
rect 10048 -1491 10108 -1460
rect 10166 -1491 10226 -1460
rect 10284 -1491 10344 -1460
rect 10402 -1491 10462 -1460
rect 10520 -1491 10580 -1460
rect 10638 -1491 10698 -1460
rect 4853 -1507 4919 -1491
rect 4853 -1541 4869 -1507
rect 4903 -1541 4919 -1507
rect 4853 -1615 4919 -1541
rect 4853 -1649 4869 -1615
rect 4903 -1649 4919 -1615
rect 4853 -1665 4919 -1649
rect 4971 -1507 5037 -1491
rect 4971 -1541 4987 -1507
rect 5021 -1541 5037 -1507
rect 4971 -1615 5037 -1541
rect 4971 -1649 4987 -1615
rect 5021 -1649 5037 -1615
rect 4971 -1665 5037 -1649
rect 5089 -1507 5155 -1491
rect 5089 -1541 5105 -1507
rect 5139 -1541 5155 -1507
rect 5089 -1615 5155 -1541
rect 5089 -1649 5105 -1615
rect 5139 -1649 5155 -1615
rect 5089 -1665 5155 -1649
rect 5207 -1507 5273 -1491
rect 5207 -1541 5223 -1507
rect 5257 -1541 5273 -1507
rect 5207 -1615 5273 -1541
rect 5207 -1649 5223 -1615
rect 5257 -1649 5273 -1615
rect 5207 -1665 5273 -1649
rect 5325 -1507 5391 -1491
rect 5325 -1541 5341 -1507
rect 5375 -1541 5391 -1507
rect 5325 -1615 5391 -1541
rect 5325 -1649 5341 -1615
rect 5375 -1649 5391 -1615
rect 5325 -1665 5391 -1649
rect 5443 -1507 5509 -1491
rect 5443 -1541 5459 -1507
rect 5493 -1541 5509 -1507
rect 5443 -1615 5509 -1541
rect 5443 -1649 5459 -1615
rect 5493 -1649 5509 -1615
rect 5443 -1665 5509 -1649
rect 5561 -1507 5627 -1491
rect 5561 -1541 5577 -1507
rect 5611 -1541 5627 -1507
rect 5561 -1615 5627 -1541
rect 5561 -1649 5577 -1615
rect 5611 -1649 5627 -1615
rect 5561 -1665 5627 -1649
rect 5679 -1507 5745 -1491
rect 5679 -1541 5695 -1507
rect 5729 -1541 5745 -1507
rect 5679 -1615 5745 -1541
rect 5679 -1649 5695 -1615
rect 5729 -1649 5745 -1615
rect 5679 -1665 5745 -1649
rect 5797 -1507 5863 -1491
rect 5797 -1541 5813 -1507
rect 5847 -1541 5863 -1507
rect 5797 -1615 5863 -1541
rect 5797 -1649 5813 -1615
rect 5847 -1649 5863 -1615
rect 5797 -1665 5863 -1649
rect 5915 -1507 5981 -1491
rect 5915 -1541 5931 -1507
rect 5965 -1541 5981 -1507
rect 5915 -1615 5981 -1541
rect 5915 -1649 5931 -1615
rect 5965 -1649 5981 -1615
rect 5915 -1665 5981 -1649
rect 6033 -1507 6099 -1491
rect 6033 -1541 6049 -1507
rect 6083 -1541 6099 -1507
rect 6033 -1615 6099 -1541
rect 6033 -1649 6049 -1615
rect 6083 -1649 6099 -1615
rect 6033 -1665 6099 -1649
rect 6151 -1507 6217 -1491
rect 6151 -1541 6167 -1507
rect 6201 -1541 6217 -1507
rect 6151 -1615 6217 -1541
rect 6151 -1649 6167 -1615
rect 6201 -1649 6217 -1615
rect 6151 -1665 6217 -1649
rect 6269 -1507 6335 -1491
rect 6269 -1541 6285 -1507
rect 6319 -1541 6335 -1507
rect 6269 -1615 6335 -1541
rect 6269 -1649 6285 -1615
rect 6319 -1649 6335 -1615
rect 6269 -1665 6335 -1649
rect 6387 -1507 6453 -1491
rect 6387 -1541 6403 -1507
rect 6437 -1541 6453 -1507
rect 6387 -1615 6453 -1541
rect 6387 -1649 6403 -1615
rect 6437 -1649 6453 -1615
rect 6387 -1665 6453 -1649
rect 6505 -1507 6571 -1491
rect 6505 -1541 6521 -1507
rect 6555 -1541 6571 -1507
rect 6505 -1615 6571 -1541
rect 6505 -1649 6521 -1615
rect 6555 -1649 6571 -1615
rect 6505 -1665 6571 -1649
rect 6623 -1507 6689 -1491
rect 6623 -1541 6639 -1507
rect 6673 -1541 6689 -1507
rect 6623 -1615 6689 -1541
rect 6623 -1649 6639 -1615
rect 6673 -1649 6689 -1615
rect 6623 -1665 6689 -1649
rect 6741 -1507 6807 -1491
rect 6741 -1541 6757 -1507
rect 6791 -1541 6807 -1507
rect 6741 -1615 6807 -1541
rect 6741 -1649 6757 -1615
rect 6791 -1649 6807 -1615
rect 6741 -1665 6807 -1649
rect 6859 -1507 6925 -1491
rect 6859 -1541 6875 -1507
rect 6909 -1541 6925 -1507
rect 6859 -1615 6925 -1541
rect 6859 -1649 6875 -1615
rect 6909 -1649 6925 -1615
rect 6859 -1665 6925 -1649
rect 6977 -1507 7043 -1491
rect 6977 -1541 6993 -1507
rect 7027 -1541 7043 -1507
rect 6977 -1615 7043 -1541
rect 6977 -1649 6993 -1615
rect 7027 -1649 7043 -1615
rect 6977 -1665 7043 -1649
rect 7095 -1507 7161 -1491
rect 7095 -1541 7111 -1507
rect 7145 -1541 7161 -1507
rect 7095 -1615 7161 -1541
rect 7095 -1649 7111 -1615
rect 7145 -1649 7161 -1615
rect 7095 -1665 7161 -1649
rect 7213 -1507 7279 -1491
rect 7213 -1541 7229 -1507
rect 7263 -1541 7279 -1507
rect 7213 -1615 7279 -1541
rect 7213 -1649 7229 -1615
rect 7263 -1649 7279 -1615
rect 7213 -1665 7279 -1649
rect 7331 -1507 7397 -1491
rect 7331 -1541 7347 -1507
rect 7381 -1541 7397 -1507
rect 7331 -1615 7397 -1541
rect 7331 -1649 7347 -1615
rect 7381 -1649 7397 -1615
rect 7331 -1665 7397 -1649
rect 7449 -1507 7515 -1491
rect 7449 -1541 7465 -1507
rect 7499 -1541 7515 -1507
rect 7449 -1615 7515 -1541
rect 7449 -1649 7465 -1615
rect 7499 -1649 7515 -1615
rect 7449 -1665 7515 -1649
rect 7567 -1507 7633 -1491
rect 7567 -1541 7583 -1507
rect 7617 -1541 7633 -1507
rect 7567 -1615 7633 -1541
rect 7567 -1649 7583 -1615
rect 7617 -1649 7633 -1615
rect 7567 -1665 7633 -1649
rect 7685 -1507 7751 -1491
rect 7685 -1541 7701 -1507
rect 7735 -1541 7751 -1507
rect 7685 -1615 7751 -1541
rect 7685 -1649 7701 -1615
rect 7735 -1649 7751 -1615
rect 7685 -1665 7751 -1649
rect 7803 -1507 7869 -1491
rect 7803 -1541 7819 -1507
rect 7853 -1541 7869 -1507
rect 7803 -1615 7869 -1541
rect 7803 -1649 7819 -1615
rect 7853 -1649 7869 -1615
rect 7803 -1665 7869 -1649
rect 7921 -1507 7987 -1491
rect 7921 -1541 7937 -1507
rect 7971 -1541 7987 -1507
rect 7921 -1615 7987 -1541
rect 7921 -1649 7937 -1615
rect 7971 -1649 7987 -1615
rect 7921 -1665 7987 -1649
rect 8039 -1507 8105 -1491
rect 8039 -1541 8055 -1507
rect 8089 -1541 8105 -1507
rect 8039 -1615 8105 -1541
rect 8039 -1649 8055 -1615
rect 8089 -1649 8105 -1615
rect 8039 -1665 8105 -1649
rect 8157 -1507 8223 -1491
rect 8157 -1541 8173 -1507
rect 8207 -1541 8223 -1507
rect 8157 -1615 8223 -1541
rect 8157 -1649 8173 -1615
rect 8207 -1649 8223 -1615
rect 8157 -1665 8223 -1649
rect 8275 -1507 8341 -1491
rect 8275 -1541 8291 -1507
rect 8325 -1541 8341 -1507
rect 8275 -1615 8341 -1541
rect 8275 -1649 8291 -1615
rect 8325 -1649 8341 -1615
rect 8275 -1665 8341 -1649
rect 8393 -1507 8459 -1491
rect 8393 -1541 8409 -1507
rect 8443 -1541 8459 -1507
rect 8393 -1615 8459 -1541
rect 8393 -1649 8409 -1615
rect 8443 -1649 8459 -1615
rect 8393 -1665 8459 -1649
rect 8511 -1507 8577 -1491
rect 8511 -1541 8527 -1507
rect 8561 -1541 8577 -1507
rect 8511 -1615 8577 -1541
rect 8511 -1649 8527 -1615
rect 8561 -1649 8577 -1615
rect 8511 -1665 8577 -1649
rect 8629 -1507 8695 -1491
rect 8629 -1541 8645 -1507
rect 8679 -1541 8695 -1507
rect 8629 -1615 8695 -1541
rect 8629 -1649 8645 -1615
rect 8679 -1649 8695 -1615
rect 8629 -1665 8695 -1649
rect 8747 -1507 8813 -1491
rect 8747 -1541 8763 -1507
rect 8797 -1541 8813 -1507
rect 8747 -1615 8813 -1541
rect 8747 -1649 8763 -1615
rect 8797 -1649 8813 -1615
rect 8747 -1665 8813 -1649
rect 8865 -1507 8931 -1491
rect 8865 -1541 8881 -1507
rect 8915 -1541 8931 -1507
rect 8865 -1615 8931 -1541
rect 8865 -1649 8881 -1615
rect 8915 -1649 8931 -1615
rect 8865 -1665 8931 -1649
rect 8983 -1507 9049 -1491
rect 8983 -1541 8999 -1507
rect 9033 -1541 9049 -1507
rect 8983 -1615 9049 -1541
rect 8983 -1649 8999 -1615
rect 9033 -1649 9049 -1615
rect 8983 -1665 9049 -1649
rect 9101 -1507 9167 -1491
rect 9101 -1541 9117 -1507
rect 9151 -1541 9167 -1507
rect 9101 -1615 9167 -1541
rect 9101 -1649 9117 -1615
rect 9151 -1649 9167 -1615
rect 9101 -1665 9167 -1649
rect 9219 -1507 9285 -1491
rect 9219 -1541 9235 -1507
rect 9269 -1541 9285 -1507
rect 9219 -1615 9285 -1541
rect 9219 -1649 9235 -1615
rect 9269 -1649 9285 -1615
rect 9219 -1665 9285 -1649
rect 9337 -1507 9403 -1491
rect 9337 -1541 9353 -1507
rect 9387 -1541 9403 -1507
rect 9337 -1615 9403 -1541
rect 9337 -1649 9353 -1615
rect 9387 -1649 9403 -1615
rect 9337 -1665 9403 -1649
rect 9455 -1507 9521 -1491
rect 9455 -1541 9471 -1507
rect 9505 -1541 9521 -1507
rect 9455 -1615 9521 -1541
rect 9455 -1649 9471 -1615
rect 9505 -1649 9521 -1615
rect 9455 -1665 9521 -1649
rect 9573 -1507 9639 -1491
rect 9573 -1541 9589 -1507
rect 9623 -1541 9639 -1507
rect 9573 -1615 9639 -1541
rect 9573 -1649 9589 -1615
rect 9623 -1649 9639 -1615
rect 9573 -1665 9639 -1649
rect 9691 -1507 9757 -1491
rect 9691 -1541 9707 -1507
rect 9741 -1541 9757 -1507
rect 9691 -1615 9757 -1541
rect 9691 -1649 9707 -1615
rect 9741 -1649 9757 -1615
rect 9691 -1665 9757 -1649
rect 9809 -1507 9875 -1491
rect 9809 -1541 9825 -1507
rect 9859 -1541 9875 -1507
rect 9809 -1615 9875 -1541
rect 9809 -1649 9825 -1615
rect 9859 -1649 9875 -1615
rect 9809 -1665 9875 -1649
rect 9927 -1507 9993 -1491
rect 9927 -1541 9943 -1507
rect 9977 -1541 9993 -1507
rect 9927 -1615 9993 -1541
rect 9927 -1649 9943 -1615
rect 9977 -1649 9993 -1615
rect 9927 -1665 9993 -1649
rect 10045 -1507 10111 -1491
rect 10045 -1541 10061 -1507
rect 10095 -1541 10111 -1507
rect 10045 -1615 10111 -1541
rect 10045 -1649 10061 -1615
rect 10095 -1649 10111 -1615
rect 10045 -1665 10111 -1649
rect 10163 -1507 10229 -1491
rect 10163 -1541 10179 -1507
rect 10213 -1541 10229 -1507
rect 10163 -1615 10229 -1541
rect 10163 -1649 10179 -1615
rect 10213 -1649 10229 -1615
rect 10163 -1665 10229 -1649
rect 10281 -1507 10347 -1491
rect 10281 -1541 10297 -1507
rect 10331 -1541 10347 -1507
rect 10281 -1615 10347 -1541
rect 10281 -1649 10297 -1615
rect 10331 -1649 10347 -1615
rect 10281 -1665 10347 -1649
rect 10399 -1507 10465 -1491
rect 10399 -1541 10415 -1507
rect 10449 -1541 10465 -1507
rect 10399 -1615 10465 -1541
rect 10399 -1649 10415 -1615
rect 10449 -1649 10465 -1615
rect 10399 -1665 10465 -1649
rect 10517 -1507 10583 -1491
rect 10517 -1541 10533 -1507
rect 10567 -1541 10583 -1507
rect 10517 -1615 10583 -1541
rect 10517 -1649 10533 -1615
rect 10567 -1649 10583 -1615
rect 10517 -1665 10583 -1649
rect 10635 -1507 10701 -1491
rect 10635 -1541 10651 -1507
rect 10685 -1541 10701 -1507
rect 10635 -1615 10701 -1541
rect 10635 -1649 10651 -1615
rect 10685 -1649 10701 -1615
rect 10635 -1665 10701 -1649
rect 4856 -1696 4916 -1665
rect 4974 -1696 5034 -1665
rect 5092 -1696 5152 -1665
rect 5210 -1696 5270 -1665
rect 5328 -1696 5388 -1665
rect 5446 -1696 5506 -1665
rect 5564 -1696 5624 -1665
rect 5682 -1696 5742 -1665
rect 5800 -1696 5860 -1665
rect 5918 -1696 5978 -1665
rect 6036 -1696 6096 -1665
rect 6154 -1696 6214 -1665
rect 6272 -1696 6332 -1665
rect 6390 -1696 6450 -1665
rect 6508 -1696 6568 -1665
rect 6626 -1696 6686 -1665
rect 6744 -1696 6804 -1665
rect 6862 -1696 6922 -1665
rect 6980 -1696 7040 -1665
rect 7098 -1696 7158 -1665
rect 7216 -1696 7276 -1665
rect 7334 -1696 7394 -1665
rect 7452 -1696 7512 -1665
rect 7570 -1696 7630 -1665
rect 7688 -1696 7748 -1665
rect 7806 -1696 7866 -1665
rect 7924 -1696 7984 -1665
rect 8042 -1696 8102 -1665
rect 8160 -1696 8220 -1665
rect 8278 -1696 8338 -1665
rect 8396 -1696 8456 -1665
rect 8514 -1696 8574 -1665
rect 8632 -1696 8692 -1665
rect 8750 -1696 8810 -1665
rect 8868 -1696 8928 -1665
rect 8986 -1696 9046 -1665
rect 9104 -1696 9164 -1665
rect 9222 -1696 9282 -1665
rect 9340 -1696 9400 -1665
rect 9458 -1696 9518 -1665
rect 9576 -1696 9636 -1665
rect 9694 -1696 9754 -1665
rect 9812 -1696 9872 -1665
rect 9930 -1696 9990 -1665
rect 10048 -1696 10108 -1665
rect 10166 -1696 10226 -1665
rect 10284 -1696 10344 -1665
rect 10402 -1696 10462 -1665
rect 10520 -1696 10580 -1665
rect 10638 -1696 10698 -1665
rect 4856 -2327 4916 -2296
rect 4974 -2327 5034 -2296
rect 5092 -2327 5152 -2296
rect 5210 -2327 5270 -2296
rect 5328 -2327 5388 -2296
rect 5446 -2327 5506 -2296
rect 5564 -2327 5624 -2296
rect 5682 -2327 5742 -2296
rect 5800 -2327 5860 -2296
rect 5918 -2327 5978 -2296
rect 6036 -2327 6096 -2296
rect 6154 -2327 6214 -2296
rect 6272 -2327 6332 -2296
rect 6390 -2327 6450 -2296
rect 6508 -2327 6568 -2296
rect 6626 -2327 6686 -2296
rect 6744 -2327 6804 -2296
rect 6862 -2327 6922 -2296
rect 6980 -2327 7040 -2296
rect 7098 -2327 7158 -2296
rect 7216 -2327 7276 -2296
rect 7334 -2327 7394 -2296
rect 7452 -2327 7512 -2296
rect 7570 -2327 7630 -2296
rect 7688 -2327 7748 -2296
rect 7806 -2327 7866 -2296
rect 7924 -2327 7984 -2296
rect 8042 -2327 8102 -2296
rect 8160 -2327 8220 -2296
rect 8278 -2327 8338 -2296
rect 8396 -2327 8456 -2296
rect 8514 -2327 8574 -2296
rect 8632 -2327 8692 -2296
rect 8750 -2327 8810 -2296
rect 8868 -2327 8928 -2296
rect 8986 -2327 9046 -2296
rect 9104 -2327 9164 -2296
rect 9222 -2327 9282 -2296
rect 9340 -2327 9400 -2296
rect 9458 -2327 9518 -2296
rect 9576 -2327 9636 -2296
rect 9694 -2327 9754 -2296
rect 9812 -2327 9872 -2296
rect 9930 -2327 9990 -2296
rect 10048 -2327 10108 -2296
rect 10166 -2327 10226 -2296
rect 10284 -2327 10344 -2296
rect 10402 -2327 10462 -2296
rect 10520 -2327 10580 -2296
rect 10638 -2327 10698 -2296
rect 4853 -2393 4919 -2327
rect 4971 -2393 5037 -2327
rect 5089 -2393 5155 -2327
rect 5207 -2393 5273 -2327
rect 5325 -2393 5391 -2327
rect 5443 -2393 5509 -2327
rect 5561 -2393 5627 -2327
rect 5679 -2393 5745 -2327
rect 5797 -2393 5863 -2327
rect 5915 -2393 5981 -2327
rect 6033 -2393 6099 -2327
rect 6151 -2393 6217 -2327
rect 6269 -2393 6335 -2327
rect 6387 -2393 6453 -2327
rect 6505 -2393 6571 -2327
rect 6623 -2393 6689 -2327
rect 6741 -2393 6807 -2327
rect 6859 -2393 6925 -2327
rect 6977 -2393 7043 -2327
rect 7095 -2393 7161 -2327
rect 7213 -2393 7279 -2327
rect 7331 -2393 7397 -2327
rect 7449 -2393 7515 -2327
rect 7567 -2393 7633 -2327
rect 7685 -2393 7751 -2327
rect 7803 -2393 7869 -2327
rect 7921 -2393 7987 -2327
rect 8039 -2393 8105 -2327
rect 8157 -2393 8223 -2327
rect 8275 -2393 8341 -2327
rect 8393 -2393 8459 -2327
rect 8511 -2393 8577 -2327
rect 8629 -2393 8695 -2327
rect 8747 -2393 8813 -2327
rect 8865 -2393 8931 -2327
rect 8983 -2393 9049 -2327
rect 9101 -2393 9167 -2327
rect 9219 -2393 9285 -2327
rect 9337 -2393 9403 -2327
rect 9455 -2393 9521 -2327
rect 9573 -2393 9639 -2327
rect 9691 -2393 9757 -2327
rect 9809 -2393 9875 -2327
rect 9927 -2393 9993 -2327
rect 10045 -2393 10111 -2327
rect 10163 -2393 10229 -2327
rect 10281 -2393 10347 -2327
rect 10399 -2393 10465 -2327
rect 10517 -2393 10583 -2327
rect 10635 -2393 10701 -2327
rect 4853 -2879 4919 -2813
rect 4971 -2879 5037 -2813
rect 5089 -2879 5155 -2813
rect 5207 -2879 5273 -2813
rect 5325 -2879 5391 -2813
rect 5443 -2879 5509 -2813
rect 5561 -2879 5627 -2813
rect 5679 -2879 5745 -2813
rect 5797 -2879 5863 -2813
rect 5915 -2879 5981 -2813
rect 6033 -2879 6099 -2813
rect 6151 -2879 6217 -2813
rect 6269 -2879 6335 -2813
rect 6387 -2879 6453 -2813
rect 6505 -2879 6571 -2813
rect 6623 -2879 6689 -2813
rect 6741 -2879 6807 -2813
rect 6859 -2879 6925 -2813
rect 6977 -2879 7043 -2813
rect 7095 -2879 7161 -2813
rect 7213 -2879 7279 -2813
rect 7331 -2879 7397 -2813
rect 7449 -2879 7515 -2813
rect 7567 -2879 7633 -2813
rect 7685 -2879 7751 -2813
rect 7803 -2879 7869 -2813
rect 7921 -2879 7987 -2813
rect 8039 -2879 8105 -2813
rect 8157 -2879 8223 -2813
rect 8275 -2879 8341 -2813
rect 8393 -2879 8459 -2813
rect 8511 -2879 8577 -2813
rect 8629 -2879 8695 -2813
rect 8747 -2879 8813 -2813
rect 8865 -2879 8931 -2813
rect 8983 -2879 9049 -2813
rect 9101 -2879 9167 -2813
rect 9219 -2879 9285 -2813
rect 9337 -2879 9403 -2813
rect 9455 -2879 9521 -2813
rect 9573 -2879 9639 -2813
rect 9691 -2879 9757 -2813
rect 9809 -2879 9875 -2813
rect 9927 -2879 9993 -2813
rect 10045 -2879 10111 -2813
rect 10163 -2879 10229 -2813
rect 10281 -2879 10347 -2813
rect 10399 -2879 10465 -2813
rect 10517 -2879 10583 -2813
rect 10635 -2879 10701 -2813
rect 4856 -2910 4916 -2879
rect 4974 -2910 5034 -2879
rect 5092 -2910 5152 -2879
rect 5210 -2910 5270 -2879
rect 5328 -2910 5388 -2879
rect 5446 -2910 5506 -2879
rect 5564 -2910 5624 -2879
rect 5682 -2910 5742 -2879
rect 5800 -2910 5860 -2879
rect 5918 -2910 5978 -2879
rect 6036 -2910 6096 -2879
rect 6154 -2910 6214 -2879
rect 6272 -2910 6332 -2879
rect 6390 -2910 6450 -2879
rect 6508 -2910 6568 -2879
rect 6626 -2910 6686 -2879
rect 6744 -2910 6804 -2879
rect 6862 -2910 6922 -2879
rect 6980 -2910 7040 -2879
rect 7098 -2910 7158 -2879
rect 7216 -2910 7276 -2879
rect 7334 -2910 7394 -2879
rect 7452 -2910 7512 -2879
rect 7570 -2910 7630 -2879
rect 7688 -2910 7748 -2879
rect 7806 -2910 7866 -2879
rect 7924 -2910 7984 -2879
rect 8042 -2910 8102 -2879
rect 8160 -2910 8220 -2879
rect 8278 -2910 8338 -2879
rect 8396 -2910 8456 -2879
rect 8514 -2910 8574 -2879
rect 8632 -2910 8692 -2879
rect 8750 -2910 8810 -2879
rect 8868 -2910 8928 -2879
rect 8986 -2910 9046 -2879
rect 9104 -2910 9164 -2879
rect 9222 -2910 9282 -2879
rect 9340 -2910 9400 -2879
rect 9458 -2910 9518 -2879
rect 9576 -2910 9636 -2879
rect 9694 -2910 9754 -2879
rect 9812 -2910 9872 -2879
rect 9930 -2910 9990 -2879
rect 10048 -2910 10108 -2879
rect 10166 -2910 10226 -2879
rect 10284 -2910 10344 -2879
rect 10402 -2910 10462 -2879
rect 10520 -2910 10580 -2879
rect 10638 -2910 10698 -2879
rect 4856 -3541 4916 -3510
rect 4974 -3541 5034 -3510
rect 5092 -3541 5152 -3510
rect 5210 -3541 5270 -3510
rect 5328 -3541 5388 -3510
rect 5446 -3541 5506 -3510
rect 5564 -3541 5624 -3510
rect 5682 -3541 5742 -3510
rect 5800 -3541 5860 -3510
rect 5918 -3541 5978 -3510
rect 6036 -3541 6096 -3510
rect 6154 -3541 6214 -3510
rect 6272 -3541 6332 -3510
rect 6390 -3541 6450 -3510
rect 6508 -3541 6568 -3510
rect 6626 -3541 6686 -3510
rect 6744 -3541 6804 -3510
rect 6862 -3541 6922 -3510
rect 6980 -3541 7040 -3510
rect 7098 -3541 7158 -3510
rect 7216 -3541 7276 -3510
rect 7334 -3541 7394 -3510
rect 7452 -3541 7512 -3510
rect 7570 -3541 7630 -3510
rect 7688 -3541 7748 -3510
rect 7806 -3541 7866 -3510
rect 7924 -3541 7984 -3510
rect 8042 -3541 8102 -3510
rect 8160 -3541 8220 -3510
rect 8278 -3541 8338 -3510
rect 8396 -3541 8456 -3510
rect 8514 -3541 8574 -3510
rect 8632 -3541 8692 -3510
rect 8750 -3541 8810 -3510
rect 8868 -3541 8928 -3510
rect 8986 -3541 9046 -3510
rect 9104 -3541 9164 -3510
rect 9222 -3541 9282 -3510
rect 9340 -3541 9400 -3510
rect 9458 -3541 9518 -3510
rect 9576 -3541 9636 -3510
rect 9694 -3541 9754 -3510
rect 9812 -3541 9872 -3510
rect 9930 -3541 9990 -3510
rect 10048 -3541 10108 -3510
rect 10166 -3541 10226 -3510
rect 10284 -3541 10344 -3510
rect 10402 -3541 10462 -3510
rect 10520 -3541 10580 -3510
rect 10638 -3541 10698 -3510
rect 4853 -3557 4919 -3541
rect 4853 -3591 4869 -3557
rect 4903 -3591 4919 -3557
rect 4853 -3665 4919 -3591
rect 4853 -3699 4869 -3665
rect 4903 -3699 4919 -3665
rect 4853 -3715 4919 -3699
rect 4971 -3557 5037 -3541
rect 4971 -3591 4987 -3557
rect 5021 -3591 5037 -3557
rect 4971 -3665 5037 -3591
rect 4971 -3699 4987 -3665
rect 5021 -3699 5037 -3665
rect 4971 -3715 5037 -3699
rect 5089 -3557 5155 -3541
rect 5089 -3591 5105 -3557
rect 5139 -3591 5155 -3557
rect 5089 -3665 5155 -3591
rect 5089 -3699 5105 -3665
rect 5139 -3699 5155 -3665
rect 5089 -3715 5155 -3699
rect 5207 -3557 5273 -3541
rect 5207 -3591 5223 -3557
rect 5257 -3591 5273 -3557
rect 5207 -3665 5273 -3591
rect 5207 -3699 5223 -3665
rect 5257 -3699 5273 -3665
rect 5207 -3715 5273 -3699
rect 5325 -3557 5391 -3541
rect 5325 -3591 5341 -3557
rect 5375 -3591 5391 -3557
rect 5325 -3665 5391 -3591
rect 5325 -3699 5341 -3665
rect 5375 -3699 5391 -3665
rect 5325 -3715 5391 -3699
rect 5443 -3557 5509 -3541
rect 5443 -3591 5459 -3557
rect 5493 -3591 5509 -3557
rect 5443 -3665 5509 -3591
rect 5443 -3699 5459 -3665
rect 5493 -3699 5509 -3665
rect 5443 -3715 5509 -3699
rect 5561 -3557 5627 -3541
rect 5561 -3591 5577 -3557
rect 5611 -3591 5627 -3557
rect 5561 -3665 5627 -3591
rect 5561 -3699 5577 -3665
rect 5611 -3699 5627 -3665
rect 5561 -3715 5627 -3699
rect 5679 -3557 5745 -3541
rect 5679 -3591 5695 -3557
rect 5729 -3591 5745 -3557
rect 5679 -3665 5745 -3591
rect 5679 -3699 5695 -3665
rect 5729 -3699 5745 -3665
rect 5679 -3715 5745 -3699
rect 5797 -3557 5863 -3541
rect 5797 -3591 5813 -3557
rect 5847 -3591 5863 -3557
rect 5797 -3665 5863 -3591
rect 5797 -3699 5813 -3665
rect 5847 -3699 5863 -3665
rect 5797 -3715 5863 -3699
rect 5915 -3557 5981 -3541
rect 5915 -3591 5931 -3557
rect 5965 -3591 5981 -3557
rect 5915 -3665 5981 -3591
rect 5915 -3699 5931 -3665
rect 5965 -3699 5981 -3665
rect 5915 -3715 5981 -3699
rect 6033 -3557 6099 -3541
rect 6033 -3591 6049 -3557
rect 6083 -3591 6099 -3557
rect 6033 -3665 6099 -3591
rect 6033 -3699 6049 -3665
rect 6083 -3699 6099 -3665
rect 6033 -3715 6099 -3699
rect 6151 -3557 6217 -3541
rect 6151 -3591 6167 -3557
rect 6201 -3591 6217 -3557
rect 6151 -3665 6217 -3591
rect 6151 -3699 6167 -3665
rect 6201 -3699 6217 -3665
rect 6151 -3715 6217 -3699
rect 6269 -3557 6335 -3541
rect 6269 -3591 6285 -3557
rect 6319 -3591 6335 -3557
rect 6269 -3665 6335 -3591
rect 6269 -3699 6285 -3665
rect 6319 -3699 6335 -3665
rect 6269 -3715 6335 -3699
rect 6387 -3557 6453 -3541
rect 6387 -3591 6403 -3557
rect 6437 -3591 6453 -3557
rect 6387 -3665 6453 -3591
rect 6387 -3699 6403 -3665
rect 6437 -3699 6453 -3665
rect 6387 -3715 6453 -3699
rect 6505 -3557 6571 -3541
rect 6505 -3591 6521 -3557
rect 6555 -3591 6571 -3557
rect 6505 -3665 6571 -3591
rect 6505 -3699 6521 -3665
rect 6555 -3699 6571 -3665
rect 6505 -3715 6571 -3699
rect 6623 -3557 6689 -3541
rect 6623 -3591 6639 -3557
rect 6673 -3591 6689 -3557
rect 6623 -3665 6689 -3591
rect 6623 -3699 6639 -3665
rect 6673 -3699 6689 -3665
rect 6623 -3715 6689 -3699
rect 6741 -3557 6807 -3541
rect 6741 -3591 6757 -3557
rect 6791 -3591 6807 -3557
rect 6741 -3665 6807 -3591
rect 6741 -3699 6757 -3665
rect 6791 -3699 6807 -3665
rect 6741 -3715 6807 -3699
rect 6859 -3557 6925 -3541
rect 6859 -3591 6875 -3557
rect 6909 -3591 6925 -3557
rect 6859 -3665 6925 -3591
rect 6859 -3699 6875 -3665
rect 6909 -3699 6925 -3665
rect 6859 -3715 6925 -3699
rect 6977 -3557 7043 -3541
rect 6977 -3591 6993 -3557
rect 7027 -3591 7043 -3557
rect 6977 -3665 7043 -3591
rect 6977 -3699 6993 -3665
rect 7027 -3699 7043 -3665
rect 6977 -3715 7043 -3699
rect 7095 -3557 7161 -3541
rect 7095 -3591 7111 -3557
rect 7145 -3591 7161 -3557
rect 7095 -3665 7161 -3591
rect 7095 -3699 7111 -3665
rect 7145 -3699 7161 -3665
rect 7095 -3715 7161 -3699
rect 7213 -3557 7279 -3541
rect 7213 -3591 7229 -3557
rect 7263 -3591 7279 -3557
rect 7213 -3665 7279 -3591
rect 7213 -3699 7229 -3665
rect 7263 -3699 7279 -3665
rect 7213 -3715 7279 -3699
rect 7331 -3557 7397 -3541
rect 7331 -3591 7347 -3557
rect 7381 -3591 7397 -3557
rect 7331 -3665 7397 -3591
rect 7331 -3699 7347 -3665
rect 7381 -3699 7397 -3665
rect 7331 -3715 7397 -3699
rect 7449 -3557 7515 -3541
rect 7449 -3591 7465 -3557
rect 7499 -3591 7515 -3557
rect 7449 -3665 7515 -3591
rect 7449 -3699 7465 -3665
rect 7499 -3699 7515 -3665
rect 7449 -3715 7515 -3699
rect 7567 -3557 7633 -3541
rect 7567 -3591 7583 -3557
rect 7617 -3591 7633 -3557
rect 7567 -3665 7633 -3591
rect 7567 -3699 7583 -3665
rect 7617 -3699 7633 -3665
rect 7567 -3715 7633 -3699
rect 7685 -3557 7751 -3541
rect 7685 -3591 7701 -3557
rect 7735 -3591 7751 -3557
rect 7685 -3665 7751 -3591
rect 7685 -3699 7701 -3665
rect 7735 -3699 7751 -3665
rect 7685 -3715 7751 -3699
rect 7803 -3557 7869 -3541
rect 7803 -3591 7819 -3557
rect 7853 -3591 7869 -3557
rect 7803 -3665 7869 -3591
rect 7803 -3699 7819 -3665
rect 7853 -3699 7869 -3665
rect 7803 -3715 7869 -3699
rect 7921 -3557 7987 -3541
rect 7921 -3591 7937 -3557
rect 7971 -3591 7987 -3557
rect 7921 -3665 7987 -3591
rect 7921 -3699 7937 -3665
rect 7971 -3699 7987 -3665
rect 7921 -3715 7987 -3699
rect 8039 -3557 8105 -3541
rect 8039 -3591 8055 -3557
rect 8089 -3591 8105 -3557
rect 8039 -3665 8105 -3591
rect 8039 -3699 8055 -3665
rect 8089 -3699 8105 -3665
rect 8039 -3715 8105 -3699
rect 8157 -3557 8223 -3541
rect 8157 -3591 8173 -3557
rect 8207 -3591 8223 -3557
rect 8157 -3665 8223 -3591
rect 8157 -3699 8173 -3665
rect 8207 -3699 8223 -3665
rect 8157 -3715 8223 -3699
rect 8275 -3557 8341 -3541
rect 8275 -3591 8291 -3557
rect 8325 -3591 8341 -3557
rect 8275 -3665 8341 -3591
rect 8275 -3699 8291 -3665
rect 8325 -3699 8341 -3665
rect 8275 -3715 8341 -3699
rect 8393 -3557 8459 -3541
rect 8393 -3591 8409 -3557
rect 8443 -3591 8459 -3557
rect 8393 -3665 8459 -3591
rect 8393 -3699 8409 -3665
rect 8443 -3699 8459 -3665
rect 8393 -3715 8459 -3699
rect 8511 -3557 8577 -3541
rect 8511 -3591 8527 -3557
rect 8561 -3591 8577 -3557
rect 8511 -3665 8577 -3591
rect 8511 -3699 8527 -3665
rect 8561 -3699 8577 -3665
rect 8511 -3715 8577 -3699
rect 8629 -3557 8695 -3541
rect 8629 -3591 8645 -3557
rect 8679 -3591 8695 -3557
rect 8629 -3665 8695 -3591
rect 8629 -3699 8645 -3665
rect 8679 -3699 8695 -3665
rect 8629 -3715 8695 -3699
rect 8747 -3557 8813 -3541
rect 8747 -3591 8763 -3557
rect 8797 -3591 8813 -3557
rect 8747 -3665 8813 -3591
rect 8747 -3699 8763 -3665
rect 8797 -3699 8813 -3665
rect 8747 -3715 8813 -3699
rect 8865 -3557 8931 -3541
rect 8865 -3591 8881 -3557
rect 8915 -3591 8931 -3557
rect 8865 -3665 8931 -3591
rect 8865 -3699 8881 -3665
rect 8915 -3699 8931 -3665
rect 8865 -3715 8931 -3699
rect 8983 -3557 9049 -3541
rect 8983 -3591 8999 -3557
rect 9033 -3591 9049 -3557
rect 8983 -3665 9049 -3591
rect 8983 -3699 8999 -3665
rect 9033 -3699 9049 -3665
rect 8983 -3715 9049 -3699
rect 9101 -3557 9167 -3541
rect 9101 -3591 9117 -3557
rect 9151 -3591 9167 -3557
rect 9101 -3665 9167 -3591
rect 9101 -3699 9117 -3665
rect 9151 -3699 9167 -3665
rect 9101 -3715 9167 -3699
rect 9219 -3557 9285 -3541
rect 9219 -3591 9235 -3557
rect 9269 -3591 9285 -3557
rect 9219 -3665 9285 -3591
rect 9219 -3699 9235 -3665
rect 9269 -3699 9285 -3665
rect 9219 -3715 9285 -3699
rect 9337 -3557 9403 -3541
rect 9337 -3591 9353 -3557
rect 9387 -3591 9403 -3557
rect 9337 -3665 9403 -3591
rect 9337 -3699 9353 -3665
rect 9387 -3699 9403 -3665
rect 9337 -3715 9403 -3699
rect 9455 -3557 9521 -3541
rect 9455 -3591 9471 -3557
rect 9505 -3591 9521 -3557
rect 9455 -3665 9521 -3591
rect 9455 -3699 9471 -3665
rect 9505 -3699 9521 -3665
rect 9455 -3715 9521 -3699
rect 9573 -3557 9639 -3541
rect 9573 -3591 9589 -3557
rect 9623 -3591 9639 -3557
rect 9573 -3665 9639 -3591
rect 9573 -3699 9589 -3665
rect 9623 -3699 9639 -3665
rect 9573 -3715 9639 -3699
rect 9691 -3557 9757 -3541
rect 9691 -3591 9707 -3557
rect 9741 -3591 9757 -3557
rect 9691 -3665 9757 -3591
rect 9691 -3699 9707 -3665
rect 9741 -3699 9757 -3665
rect 9691 -3715 9757 -3699
rect 9809 -3557 9875 -3541
rect 9809 -3591 9825 -3557
rect 9859 -3591 9875 -3557
rect 9809 -3665 9875 -3591
rect 9809 -3699 9825 -3665
rect 9859 -3699 9875 -3665
rect 9809 -3715 9875 -3699
rect 9927 -3557 9993 -3541
rect 9927 -3591 9943 -3557
rect 9977 -3591 9993 -3557
rect 9927 -3665 9993 -3591
rect 9927 -3699 9943 -3665
rect 9977 -3699 9993 -3665
rect 9927 -3715 9993 -3699
rect 10045 -3557 10111 -3541
rect 10045 -3591 10061 -3557
rect 10095 -3591 10111 -3557
rect 10045 -3665 10111 -3591
rect 10045 -3699 10061 -3665
rect 10095 -3699 10111 -3665
rect 10045 -3715 10111 -3699
rect 10163 -3557 10229 -3541
rect 10163 -3591 10179 -3557
rect 10213 -3591 10229 -3557
rect 10163 -3665 10229 -3591
rect 10163 -3699 10179 -3665
rect 10213 -3699 10229 -3665
rect 10163 -3715 10229 -3699
rect 10281 -3557 10347 -3541
rect 10281 -3591 10297 -3557
rect 10331 -3591 10347 -3557
rect 10281 -3665 10347 -3591
rect 10281 -3699 10297 -3665
rect 10331 -3699 10347 -3665
rect 10281 -3715 10347 -3699
rect 10399 -3557 10465 -3541
rect 10399 -3591 10415 -3557
rect 10449 -3591 10465 -3557
rect 10399 -3665 10465 -3591
rect 10399 -3699 10415 -3665
rect 10449 -3699 10465 -3665
rect 10399 -3715 10465 -3699
rect 10517 -3557 10583 -3541
rect 10517 -3591 10533 -3557
rect 10567 -3591 10583 -3557
rect 10517 -3665 10583 -3591
rect 10517 -3699 10533 -3665
rect 10567 -3699 10583 -3665
rect 10517 -3715 10583 -3699
rect 10635 -3557 10701 -3541
rect 10635 -3591 10651 -3557
rect 10685 -3591 10701 -3557
rect 10635 -3665 10701 -3591
rect 10635 -3699 10651 -3665
rect 10685 -3699 10701 -3665
rect 10635 -3715 10701 -3699
rect 4856 -3746 4916 -3715
rect 4974 -3746 5034 -3715
rect 5092 -3746 5152 -3715
rect 5210 -3746 5270 -3715
rect 5328 -3746 5388 -3715
rect 5446 -3746 5506 -3715
rect 5564 -3746 5624 -3715
rect 5682 -3746 5742 -3715
rect 5800 -3746 5860 -3715
rect 5918 -3746 5978 -3715
rect 6036 -3746 6096 -3715
rect 6154 -3746 6214 -3715
rect 6272 -3746 6332 -3715
rect 6390 -3746 6450 -3715
rect 6508 -3746 6568 -3715
rect 6626 -3746 6686 -3715
rect 6744 -3746 6804 -3715
rect 6862 -3746 6922 -3715
rect 6980 -3746 7040 -3715
rect 7098 -3746 7158 -3715
rect 7216 -3746 7276 -3715
rect 7334 -3746 7394 -3715
rect 7452 -3746 7512 -3715
rect 7570 -3746 7630 -3715
rect 7688 -3746 7748 -3715
rect 7806 -3746 7866 -3715
rect 7924 -3746 7984 -3715
rect 8042 -3746 8102 -3715
rect 8160 -3746 8220 -3715
rect 8278 -3746 8338 -3715
rect 8396 -3746 8456 -3715
rect 8514 -3746 8574 -3715
rect 8632 -3746 8692 -3715
rect 8750 -3746 8810 -3715
rect 8868 -3746 8928 -3715
rect 8986 -3746 9046 -3715
rect 9104 -3746 9164 -3715
rect 9222 -3746 9282 -3715
rect 9340 -3746 9400 -3715
rect 9458 -3746 9518 -3715
rect 9576 -3746 9636 -3715
rect 9694 -3746 9754 -3715
rect 9812 -3746 9872 -3715
rect 9930 -3746 9990 -3715
rect 10048 -3746 10108 -3715
rect 10166 -3746 10226 -3715
rect 10284 -3746 10344 -3715
rect 10402 -3746 10462 -3715
rect 10520 -3746 10580 -3715
rect 10638 -3746 10698 -3715
rect 4856 -4377 4916 -4346
rect 4974 -4377 5034 -4346
rect 5092 -4377 5152 -4346
rect 5210 -4377 5270 -4346
rect 5328 -4377 5388 -4346
rect 5446 -4377 5506 -4346
rect 5564 -4377 5624 -4346
rect 5682 -4377 5742 -4346
rect 5800 -4377 5860 -4346
rect 5918 -4377 5978 -4346
rect 6036 -4377 6096 -4346
rect 6154 -4377 6214 -4346
rect 6272 -4377 6332 -4346
rect 6390 -4377 6450 -4346
rect 6508 -4377 6568 -4346
rect 6626 -4377 6686 -4346
rect 6744 -4377 6804 -4346
rect 6862 -4377 6922 -4346
rect 6980 -4377 7040 -4346
rect 7098 -4377 7158 -4346
rect 7216 -4377 7276 -4346
rect 7334 -4377 7394 -4346
rect 7452 -4377 7512 -4346
rect 7570 -4377 7630 -4346
rect 7688 -4377 7748 -4346
rect 7806 -4377 7866 -4346
rect 7924 -4377 7984 -4346
rect 8042 -4377 8102 -4346
rect 8160 -4377 8220 -4346
rect 8278 -4377 8338 -4346
rect 8396 -4377 8456 -4346
rect 8514 -4377 8574 -4346
rect 8632 -4377 8692 -4346
rect 8750 -4377 8810 -4346
rect 8868 -4377 8928 -4346
rect 8986 -4377 9046 -4346
rect 9104 -4377 9164 -4346
rect 9222 -4377 9282 -4346
rect 9340 -4377 9400 -4346
rect 9458 -4377 9518 -4346
rect 9576 -4377 9636 -4346
rect 9694 -4377 9754 -4346
rect 9812 -4377 9872 -4346
rect 9930 -4377 9990 -4346
rect 10048 -4377 10108 -4346
rect 10166 -4377 10226 -4346
rect 10284 -4377 10344 -4346
rect 10402 -4377 10462 -4346
rect 10520 -4377 10580 -4346
rect 10638 -4377 10698 -4346
rect 4853 -4443 4919 -4377
rect 4971 -4443 5037 -4377
rect 5089 -4443 5155 -4377
rect 5207 -4443 5273 -4377
rect 5325 -4443 5391 -4377
rect 5443 -4443 5509 -4377
rect 5561 -4443 5627 -4377
rect 5679 -4443 5745 -4377
rect 5797 -4443 5863 -4377
rect 5915 -4443 5981 -4377
rect 6033 -4443 6099 -4377
rect 6151 -4443 6217 -4377
rect 6269 -4443 6335 -4377
rect 6387 -4443 6453 -4377
rect 6505 -4443 6571 -4377
rect 6623 -4443 6689 -4377
rect 6741 -4443 6807 -4377
rect 6859 -4443 6925 -4377
rect 6977 -4443 7043 -4377
rect 7095 -4443 7161 -4377
rect 7213 -4443 7279 -4377
rect 7331 -4443 7397 -4377
rect 7449 -4443 7515 -4377
rect 7567 -4443 7633 -4377
rect 7685 -4443 7751 -4377
rect 7803 -4443 7869 -4377
rect 7921 -4443 7987 -4377
rect 8039 -4443 8105 -4377
rect 8157 -4443 8223 -4377
rect 8275 -4443 8341 -4377
rect 8393 -4443 8459 -4377
rect 8511 -4443 8577 -4377
rect 8629 -4443 8695 -4377
rect 8747 -4443 8813 -4377
rect 8865 -4443 8931 -4377
rect 8983 -4443 9049 -4377
rect 9101 -4443 9167 -4377
rect 9219 -4443 9285 -4377
rect 9337 -4443 9403 -4377
rect 9455 -4443 9521 -4377
rect 9573 -4443 9639 -4377
rect 9691 -4443 9757 -4377
rect 9809 -4443 9875 -4377
rect 9927 -4443 9993 -4377
rect 10045 -4443 10111 -4377
rect 10163 -4443 10229 -4377
rect 10281 -4443 10347 -4377
rect 10399 -4443 10465 -4377
rect 10517 -4443 10583 -4377
rect 10635 -4443 10701 -4377
rect 4853 -5607 4919 -5591
rect 4853 -5641 4869 -5607
rect 4903 -5641 4919 -5607
rect 4853 -5715 4919 -5641
rect 4853 -5749 4869 -5715
rect 4903 -5749 4919 -5715
rect 4853 -5765 4919 -5749
rect 4971 -5607 5037 -5591
rect 4971 -5641 4987 -5607
rect 5021 -5641 5037 -5607
rect 4971 -5715 5037 -5641
rect 4971 -5749 4987 -5715
rect 5021 -5749 5037 -5715
rect 4971 -5765 5037 -5749
rect 5089 -5607 5155 -5591
rect 5089 -5641 5105 -5607
rect 5139 -5641 5155 -5607
rect 5089 -5715 5155 -5641
rect 5089 -5749 5105 -5715
rect 5139 -5749 5155 -5715
rect 5089 -5765 5155 -5749
rect 5207 -5607 5273 -5591
rect 5207 -5641 5223 -5607
rect 5257 -5641 5273 -5607
rect 5207 -5715 5273 -5641
rect 5207 -5749 5223 -5715
rect 5257 -5749 5273 -5715
rect 5207 -5765 5273 -5749
rect 5325 -5607 5391 -5591
rect 5325 -5641 5341 -5607
rect 5375 -5641 5391 -5607
rect 5325 -5715 5391 -5641
rect 5325 -5749 5341 -5715
rect 5375 -5749 5391 -5715
rect 5325 -5765 5391 -5749
rect 5443 -5607 5509 -5591
rect 5443 -5641 5459 -5607
rect 5493 -5641 5509 -5607
rect 5443 -5715 5509 -5641
rect 5443 -5749 5459 -5715
rect 5493 -5749 5509 -5715
rect 5443 -5765 5509 -5749
rect 5561 -5607 5627 -5591
rect 5561 -5641 5577 -5607
rect 5611 -5641 5627 -5607
rect 5561 -5715 5627 -5641
rect 5561 -5749 5577 -5715
rect 5611 -5749 5627 -5715
rect 5561 -5765 5627 -5749
rect 5679 -5607 5745 -5591
rect 5679 -5641 5695 -5607
rect 5729 -5641 5745 -5607
rect 5679 -5715 5745 -5641
rect 5679 -5749 5695 -5715
rect 5729 -5749 5745 -5715
rect 5679 -5765 5745 -5749
rect 5797 -5607 5863 -5591
rect 5797 -5641 5813 -5607
rect 5847 -5641 5863 -5607
rect 5797 -5715 5863 -5641
rect 5797 -5749 5813 -5715
rect 5847 -5749 5863 -5715
rect 5797 -5765 5863 -5749
rect 5915 -5607 5981 -5591
rect 5915 -5641 5931 -5607
rect 5965 -5641 5981 -5607
rect 5915 -5715 5981 -5641
rect 5915 -5749 5931 -5715
rect 5965 -5749 5981 -5715
rect 5915 -5765 5981 -5749
rect 6033 -5607 6099 -5591
rect 6033 -5641 6049 -5607
rect 6083 -5641 6099 -5607
rect 6033 -5715 6099 -5641
rect 6033 -5749 6049 -5715
rect 6083 -5749 6099 -5715
rect 6033 -5765 6099 -5749
rect 6151 -5607 6217 -5591
rect 6151 -5641 6167 -5607
rect 6201 -5641 6217 -5607
rect 6151 -5715 6217 -5641
rect 6151 -5749 6167 -5715
rect 6201 -5749 6217 -5715
rect 6151 -5765 6217 -5749
rect 6269 -5607 6335 -5591
rect 6269 -5641 6285 -5607
rect 6319 -5641 6335 -5607
rect 6269 -5715 6335 -5641
rect 6269 -5749 6285 -5715
rect 6319 -5749 6335 -5715
rect 6269 -5765 6335 -5749
rect 6387 -5607 6453 -5591
rect 6387 -5641 6403 -5607
rect 6437 -5641 6453 -5607
rect 6387 -5715 6453 -5641
rect 6387 -5749 6403 -5715
rect 6437 -5749 6453 -5715
rect 6387 -5765 6453 -5749
rect 6505 -5607 6571 -5591
rect 6505 -5641 6521 -5607
rect 6555 -5641 6571 -5607
rect 6505 -5715 6571 -5641
rect 6505 -5749 6521 -5715
rect 6555 -5749 6571 -5715
rect 6505 -5765 6571 -5749
rect 6623 -5607 6689 -5591
rect 6623 -5641 6639 -5607
rect 6673 -5641 6689 -5607
rect 6623 -5715 6689 -5641
rect 6623 -5749 6639 -5715
rect 6673 -5749 6689 -5715
rect 6623 -5765 6689 -5749
rect 6741 -5607 6807 -5591
rect 6741 -5641 6757 -5607
rect 6791 -5641 6807 -5607
rect 6741 -5715 6807 -5641
rect 6741 -5749 6757 -5715
rect 6791 -5749 6807 -5715
rect 6741 -5765 6807 -5749
rect 6859 -5607 6925 -5591
rect 6859 -5641 6875 -5607
rect 6909 -5641 6925 -5607
rect 6859 -5715 6925 -5641
rect 6859 -5749 6875 -5715
rect 6909 -5749 6925 -5715
rect 6859 -5765 6925 -5749
rect 6977 -5607 7043 -5591
rect 6977 -5641 6993 -5607
rect 7027 -5641 7043 -5607
rect 6977 -5715 7043 -5641
rect 6977 -5749 6993 -5715
rect 7027 -5749 7043 -5715
rect 6977 -5765 7043 -5749
rect 7095 -5607 7161 -5591
rect 7095 -5641 7111 -5607
rect 7145 -5641 7161 -5607
rect 7095 -5715 7161 -5641
rect 7095 -5749 7111 -5715
rect 7145 -5749 7161 -5715
rect 7095 -5765 7161 -5749
rect 7213 -5607 7279 -5591
rect 7213 -5641 7229 -5607
rect 7263 -5641 7279 -5607
rect 7213 -5715 7279 -5641
rect 7213 -5749 7229 -5715
rect 7263 -5749 7279 -5715
rect 7213 -5765 7279 -5749
rect 7331 -5607 7397 -5591
rect 7331 -5641 7347 -5607
rect 7381 -5641 7397 -5607
rect 7331 -5715 7397 -5641
rect 7331 -5749 7347 -5715
rect 7381 -5749 7397 -5715
rect 7331 -5765 7397 -5749
rect 7449 -5607 7515 -5591
rect 7449 -5641 7465 -5607
rect 7499 -5641 7515 -5607
rect 7449 -5715 7515 -5641
rect 7449 -5749 7465 -5715
rect 7499 -5749 7515 -5715
rect 7449 -5765 7515 -5749
rect 7567 -5607 7633 -5591
rect 7567 -5641 7583 -5607
rect 7617 -5641 7633 -5607
rect 7567 -5715 7633 -5641
rect 7567 -5749 7583 -5715
rect 7617 -5749 7633 -5715
rect 7567 -5765 7633 -5749
rect 7685 -5607 7751 -5591
rect 7685 -5641 7701 -5607
rect 7735 -5641 7751 -5607
rect 7685 -5715 7751 -5641
rect 7685 -5749 7701 -5715
rect 7735 -5749 7751 -5715
rect 7685 -5765 7751 -5749
rect 7803 -5607 7869 -5591
rect 7803 -5641 7819 -5607
rect 7853 -5641 7869 -5607
rect 7803 -5715 7869 -5641
rect 7803 -5749 7819 -5715
rect 7853 -5749 7869 -5715
rect 7803 -5765 7869 -5749
rect 7921 -5607 7987 -5591
rect 7921 -5641 7937 -5607
rect 7971 -5641 7987 -5607
rect 7921 -5715 7987 -5641
rect 7921 -5749 7937 -5715
rect 7971 -5749 7987 -5715
rect 7921 -5765 7987 -5749
rect 8039 -5607 8105 -5591
rect 8039 -5641 8055 -5607
rect 8089 -5641 8105 -5607
rect 8039 -5715 8105 -5641
rect 8039 -5749 8055 -5715
rect 8089 -5749 8105 -5715
rect 8039 -5765 8105 -5749
rect 8157 -5607 8223 -5591
rect 8157 -5641 8173 -5607
rect 8207 -5641 8223 -5607
rect 8157 -5715 8223 -5641
rect 8157 -5749 8173 -5715
rect 8207 -5749 8223 -5715
rect 8157 -5765 8223 -5749
rect 8275 -5607 8341 -5591
rect 8275 -5641 8291 -5607
rect 8325 -5641 8341 -5607
rect 8275 -5715 8341 -5641
rect 8275 -5749 8291 -5715
rect 8325 -5749 8341 -5715
rect 8275 -5765 8341 -5749
rect 8393 -5607 8459 -5591
rect 8393 -5641 8409 -5607
rect 8443 -5641 8459 -5607
rect 8393 -5715 8459 -5641
rect 8393 -5749 8409 -5715
rect 8443 -5749 8459 -5715
rect 8393 -5765 8459 -5749
rect 8511 -5607 8577 -5591
rect 8511 -5641 8527 -5607
rect 8561 -5641 8577 -5607
rect 8511 -5715 8577 -5641
rect 8511 -5749 8527 -5715
rect 8561 -5749 8577 -5715
rect 8511 -5765 8577 -5749
rect 8629 -5607 8695 -5591
rect 8629 -5641 8645 -5607
rect 8679 -5641 8695 -5607
rect 8629 -5715 8695 -5641
rect 8629 -5749 8645 -5715
rect 8679 -5749 8695 -5715
rect 8629 -5765 8695 -5749
rect 8747 -5607 8813 -5591
rect 8747 -5641 8763 -5607
rect 8797 -5641 8813 -5607
rect 8747 -5715 8813 -5641
rect 8747 -5749 8763 -5715
rect 8797 -5749 8813 -5715
rect 8747 -5765 8813 -5749
rect 8865 -5607 8931 -5591
rect 8865 -5641 8881 -5607
rect 8915 -5641 8931 -5607
rect 8865 -5715 8931 -5641
rect 8865 -5749 8881 -5715
rect 8915 -5749 8931 -5715
rect 8865 -5765 8931 -5749
rect 8983 -5607 9049 -5591
rect 8983 -5641 8999 -5607
rect 9033 -5641 9049 -5607
rect 8983 -5715 9049 -5641
rect 8983 -5749 8999 -5715
rect 9033 -5749 9049 -5715
rect 8983 -5765 9049 -5749
rect 9101 -5607 9167 -5591
rect 9101 -5641 9117 -5607
rect 9151 -5641 9167 -5607
rect 9101 -5715 9167 -5641
rect 9101 -5749 9117 -5715
rect 9151 -5749 9167 -5715
rect 9101 -5765 9167 -5749
rect 9219 -5607 9285 -5591
rect 9219 -5641 9235 -5607
rect 9269 -5641 9285 -5607
rect 9219 -5715 9285 -5641
rect 9219 -5749 9235 -5715
rect 9269 -5749 9285 -5715
rect 9219 -5765 9285 -5749
rect 9337 -5607 9403 -5591
rect 9337 -5641 9353 -5607
rect 9387 -5641 9403 -5607
rect 9337 -5715 9403 -5641
rect 9337 -5749 9353 -5715
rect 9387 -5749 9403 -5715
rect 9337 -5765 9403 -5749
rect 9455 -5607 9521 -5591
rect 9455 -5641 9471 -5607
rect 9505 -5641 9521 -5607
rect 9455 -5715 9521 -5641
rect 9455 -5749 9471 -5715
rect 9505 -5749 9521 -5715
rect 9455 -5765 9521 -5749
rect 9573 -5607 9639 -5591
rect 9573 -5641 9589 -5607
rect 9623 -5641 9639 -5607
rect 9573 -5715 9639 -5641
rect 9573 -5749 9589 -5715
rect 9623 -5749 9639 -5715
rect 9573 -5765 9639 -5749
rect 9691 -5607 9757 -5591
rect 9691 -5641 9707 -5607
rect 9741 -5641 9757 -5607
rect 9691 -5715 9757 -5641
rect 9691 -5749 9707 -5715
rect 9741 -5749 9757 -5715
rect 9691 -5765 9757 -5749
rect 9809 -5607 9875 -5591
rect 9809 -5641 9825 -5607
rect 9859 -5641 9875 -5607
rect 9809 -5715 9875 -5641
rect 9809 -5749 9825 -5715
rect 9859 -5749 9875 -5715
rect 9809 -5765 9875 -5749
rect 9927 -5607 9993 -5591
rect 9927 -5641 9943 -5607
rect 9977 -5641 9993 -5607
rect 9927 -5715 9993 -5641
rect 9927 -5749 9943 -5715
rect 9977 -5749 9993 -5715
rect 9927 -5765 9993 -5749
rect 10045 -5607 10111 -5591
rect 10045 -5641 10061 -5607
rect 10095 -5641 10111 -5607
rect 10045 -5715 10111 -5641
rect 10045 -5749 10061 -5715
rect 10095 -5749 10111 -5715
rect 10045 -5765 10111 -5749
rect 10163 -5607 10229 -5591
rect 10163 -5641 10179 -5607
rect 10213 -5641 10229 -5607
rect 10163 -5715 10229 -5641
rect 10163 -5749 10179 -5715
rect 10213 -5749 10229 -5715
rect 10163 -5765 10229 -5749
rect 10281 -5607 10347 -5591
rect 10281 -5641 10297 -5607
rect 10331 -5641 10347 -5607
rect 10281 -5715 10347 -5641
rect 10281 -5749 10297 -5715
rect 10331 -5749 10347 -5715
rect 10281 -5765 10347 -5749
rect 10399 -5607 10465 -5591
rect 10399 -5641 10415 -5607
rect 10449 -5641 10465 -5607
rect 10399 -5715 10465 -5641
rect 10399 -5749 10415 -5715
rect 10449 -5749 10465 -5715
rect 10399 -5765 10465 -5749
rect 10517 -5607 10583 -5591
rect 10517 -5641 10533 -5607
rect 10567 -5641 10583 -5607
rect 10517 -5715 10583 -5641
rect 10517 -5749 10533 -5715
rect 10567 -5749 10583 -5715
rect 10517 -5765 10583 -5749
rect 10635 -5607 10701 -5591
rect 10635 -5641 10651 -5607
rect 10685 -5641 10701 -5607
rect 10635 -5715 10701 -5641
rect 10635 -5749 10651 -5715
rect 10685 -5749 10701 -5715
rect 10635 -5765 10701 -5749
rect 5919 -7841 5985 -7825
rect 5919 -7875 5935 -7841
rect 5969 -7875 5985 -7841
rect 5919 -7949 5985 -7875
rect 5919 -7983 5935 -7949
rect 5969 -7983 5985 -7949
rect 5919 -7999 5985 -7983
rect 6037 -7841 6103 -7825
rect 6037 -7875 6053 -7841
rect 6087 -7875 6103 -7841
rect 6037 -7949 6103 -7875
rect 6037 -7983 6053 -7949
rect 6087 -7983 6103 -7949
rect 6037 -7999 6103 -7983
rect 6155 -7841 6221 -7825
rect 6155 -7875 6171 -7841
rect 6205 -7875 6221 -7841
rect 6155 -7949 6221 -7875
rect 6155 -7983 6171 -7949
rect 6205 -7983 6221 -7949
rect 6155 -7999 6221 -7983
rect 6273 -7841 6339 -7825
rect 6273 -7875 6289 -7841
rect 6323 -7875 6339 -7841
rect 6273 -7949 6339 -7875
rect 6273 -7983 6289 -7949
rect 6323 -7983 6339 -7949
rect 6273 -7999 6339 -7983
rect 6391 -7841 6457 -7825
rect 6391 -7875 6407 -7841
rect 6441 -7875 6457 -7841
rect 6391 -7949 6457 -7875
rect 6391 -7983 6407 -7949
rect 6441 -7983 6457 -7949
rect 6391 -7999 6457 -7983
rect 6509 -7841 6575 -7825
rect 6509 -7875 6525 -7841
rect 6559 -7875 6575 -7841
rect 6509 -7949 6575 -7875
rect 6509 -7983 6525 -7949
rect 6559 -7983 6575 -7949
rect 6509 -7999 6575 -7983
rect 6627 -7841 6693 -7825
rect 6627 -7875 6643 -7841
rect 6677 -7875 6693 -7841
rect 6627 -7949 6693 -7875
rect 6627 -7983 6643 -7949
rect 6677 -7983 6693 -7949
rect 6627 -7999 6693 -7983
rect 6745 -7841 6811 -7825
rect 6745 -7875 6761 -7841
rect 6795 -7875 6811 -7841
rect 6745 -7949 6811 -7875
rect 6745 -7983 6761 -7949
rect 6795 -7983 6811 -7949
rect 6745 -7999 6811 -7983
rect 6863 -7841 6929 -7825
rect 6863 -7875 6879 -7841
rect 6913 -7875 6929 -7841
rect 6863 -7949 6929 -7875
rect 6863 -7983 6879 -7949
rect 6913 -7983 6929 -7949
rect 6863 -7999 6929 -7983
rect 6981 -7841 7047 -7825
rect 6981 -7875 6997 -7841
rect 7031 -7875 7047 -7841
rect 6981 -7949 7047 -7875
rect 6981 -7983 6997 -7949
rect 7031 -7983 7047 -7949
rect 6981 -7999 7047 -7983
rect 7099 -7841 7165 -7825
rect 7099 -7875 7115 -7841
rect 7149 -7875 7165 -7841
rect 7099 -7949 7165 -7875
rect 7099 -7983 7115 -7949
rect 7149 -7983 7165 -7949
rect 7099 -7999 7165 -7983
rect 7217 -7841 7283 -7825
rect 7217 -7875 7233 -7841
rect 7267 -7875 7283 -7841
rect 7217 -7949 7283 -7875
rect 7217 -7983 7233 -7949
rect 7267 -7983 7283 -7949
rect 7217 -7999 7283 -7983
rect 7335 -7841 7401 -7825
rect 7335 -7875 7351 -7841
rect 7385 -7875 7401 -7841
rect 7335 -7949 7401 -7875
rect 7335 -7983 7351 -7949
rect 7385 -7983 7401 -7949
rect 7335 -7999 7401 -7983
rect 7453 -7841 7519 -7825
rect 7453 -7875 7469 -7841
rect 7503 -7875 7519 -7841
rect 7453 -7949 7519 -7875
rect 7453 -7983 7469 -7949
rect 7503 -7983 7519 -7949
rect 7453 -7999 7519 -7983
rect 7571 -7841 7637 -7825
rect 7571 -7875 7587 -7841
rect 7621 -7875 7637 -7841
rect 7571 -7949 7637 -7875
rect 7571 -7983 7587 -7949
rect 7621 -7983 7637 -7949
rect 7571 -7999 7637 -7983
rect 7917 -7841 7983 -7825
rect 7917 -7875 7933 -7841
rect 7967 -7875 7983 -7841
rect 7917 -7949 7983 -7875
rect 7917 -7983 7933 -7949
rect 7967 -7983 7983 -7949
rect 7917 -7999 7983 -7983
rect 8035 -7841 8101 -7825
rect 8035 -7875 8051 -7841
rect 8085 -7875 8101 -7841
rect 8035 -7949 8101 -7875
rect 8035 -7983 8051 -7949
rect 8085 -7983 8101 -7949
rect 8035 -7999 8101 -7983
rect 8153 -7841 8219 -7825
rect 8153 -7875 8169 -7841
rect 8203 -7875 8219 -7841
rect 8153 -7949 8219 -7875
rect 8153 -7983 8169 -7949
rect 8203 -7983 8219 -7949
rect 8153 -7999 8219 -7983
rect 8271 -7841 8337 -7825
rect 8271 -7875 8287 -7841
rect 8321 -7875 8337 -7841
rect 8271 -7949 8337 -7875
rect 8271 -7983 8287 -7949
rect 8321 -7983 8337 -7949
rect 8271 -7999 8337 -7983
rect 8389 -7841 8455 -7825
rect 8389 -7875 8405 -7841
rect 8439 -7875 8455 -7841
rect 8389 -7949 8455 -7875
rect 8389 -7983 8405 -7949
rect 8439 -7983 8455 -7949
rect 8389 -7999 8455 -7983
rect 8507 -7841 8573 -7825
rect 8507 -7875 8523 -7841
rect 8557 -7875 8573 -7841
rect 8507 -7949 8573 -7875
rect 8507 -7983 8523 -7949
rect 8557 -7983 8573 -7949
rect 8507 -7999 8573 -7983
rect 8625 -7841 8691 -7825
rect 8625 -7875 8641 -7841
rect 8675 -7875 8691 -7841
rect 8625 -7949 8691 -7875
rect 8625 -7983 8641 -7949
rect 8675 -7983 8691 -7949
rect 8625 -7999 8691 -7983
rect 8743 -7841 8809 -7825
rect 8743 -7875 8759 -7841
rect 8793 -7875 8809 -7841
rect 8743 -7949 8809 -7875
rect 8743 -7983 8759 -7949
rect 8793 -7983 8809 -7949
rect 8743 -7999 8809 -7983
rect 8861 -7841 8927 -7825
rect 8861 -7875 8877 -7841
rect 8911 -7875 8927 -7841
rect 8861 -7949 8927 -7875
rect 8861 -7983 8877 -7949
rect 8911 -7983 8927 -7949
rect 8861 -7999 8927 -7983
rect 8979 -7841 9045 -7825
rect 8979 -7875 8995 -7841
rect 9029 -7875 9045 -7841
rect 8979 -7949 9045 -7875
rect 8979 -7983 8995 -7949
rect 9029 -7983 9045 -7949
rect 8979 -7999 9045 -7983
rect 9097 -7841 9163 -7825
rect 9097 -7875 9113 -7841
rect 9147 -7875 9163 -7841
rect 9097 -7949 9163 -7875
rect 9097 -7983 9113 -7949
rect 9147 -7983 9163 -7949
rect 9097 -7999 9163 -7983
rect 9215 -7841 9281 -7825
rect 9215 -7875 9231 -7841
rect 9265 -7875 9281 -7841
rect 9215 -7949 9281 -7875
rect 9215 -7983 9231 -7949
rect 9265 -7983 9281 -7949
rect 9215 -7999 9281 -7983
rect 9333 -7841 9399 -7825
rect 9333 -7875 9349 -7841
rect 9383 -7875 9399 -7841
rect 9333 -7949 9399 -7875
rect 9333 -7983 9349 -7949
rect 9383 -7983 9399 -7949
rect 9333 -7999 9399 -7983
rect 9451 -7841 9517 -7825
rect 9451 -7875 9467 -7841
rect 9501 -7875 9517 -7841
rect 9451 -7949 9517 -7875
rect 9451 -7983 9467 -7949
rect 9501 -7983 9517 -7949
rect 9451 -7999 9517 -7983
rect 9569 -7841 9635 -7825
rect 9569 -7875 9585 -7841
rect 9619 -7875 9635 -7841
rect 9569 -7949 9635 -7875
rect 9569 -7983 9585 -7949
rect 9619 -7983 9635 -7949
rect 9569 -7999 9635 -7983
rect 12580 -8289 12670 -8135
rect 12728 -8299 12818 -8125
rect 12876 -8299 12966 -8125
rect 13024 -8299 13114 -8125
rect 13172 -8141 13262 -8125
rect 13172 -8175 13188 -8141
rect 13246 -8175 13262 -8141
rect 13172 -8249 13262 -8175
rect 13172 -8283 13188 -8249
rect 13246 -8283 13262 -8249
rect 13172 -8299 13262 -8283
rect 13320 -8141 13410 -8125
rect 13320 -8175 13336 -8141
rect 13394 -8175 13410 -8141
rect 13320 -8249 13410 -8175
rect 13320 -8283 13336 -8249
rect 13394 -8283 13410 -8249
rect 13320 -8299 13410 -8283
rect 13468 -8141 13558 -8125
rect 13468 -8175 13484 -8141
rect 13542 -8175 13558 -8141
rect 13468 -8249 13558 -8175
rect 13468 -8283 13484 -8249
rect 13542 -8283 13558 -8249
rect 13468 -8299 13558 -8283
rect 13616 -8141 13706 -8125
rect 13616 -8175 13632 -8141
rect 13690 -8175 13706 -8141
rect 13616 -8249 13706 -8175
rect 13616 -8283 13632 -8249
rect 13690 -8283 13706 -8249
rect 13616 -8299 13706 -8283
rect 13764 -8141 13854 -8125
rect 13764 -8175 13780 -8141
rect 13838 -8175 13854 -8141
rect 13764 -8249 13854 -8175
rect 13764 -8283 13780 -8249
rect 13838 -8283 13854 -8249
rect 13764 -8299 13854 -8283
rect 13912 -8141 14002 -8125
rect 13912 -8175 13928 -8141
rect 13986 -8175 14002 -8141
rect 13912 -8249 14002 -8175
rect 13912 -8283 13928 -8249
rect 13986 -8283 14002 -8249
rect 13912 -8299 14002 -8283
rect 14060 -8299 14150 -8125
rect 14208 -8299 14298 -8125
rect 14356 -8299 14446 -8125
rect 14504 -8299 14594 -8125
rect 14652 -8141 14742 -8125
rect 14652 -8175 14668 -8141
rect 14726 -8175 14742 -8141
rect 14652 -8249 14742 -8175
rect 14652 -8283 14668 -8249
rect 14726 -8283 14742 -8249
rect 14652 -8299 14742 -8283
rect 14800 -8141 14890 -8125
rect 14800 -8175 14816 -8141
rect 14874 -8175 14890 -8141
rect 14800 -8249 14890 -8175
rect 14800 -8283 14816 -8249
rect 14874 -8283 14890 -8249
rect 14800 -8299 14890 -8283
rect 14948 -8141 15038 -8125
rect 14948 -8175 14964 -8141
rect 15022 -8175 15038 -8141
rect 14948 -8249 15038 -8175
rect 14948 -8283 14964 -8249
rect 15022 -8283 15038 -8249
rect 14948 -8299 15038 -8283
rect 15096 -8141 15186 -8125
rect 15096 -8175 15112 -8141
rect 15170 -8175 15186 -8141
rect 15096 -8249 15186 -8175
rect 15096 -8283 15112 -8249
rect 15170 -8283 15186 -8249
rect 15096 -8299 15186 -8283
rect 15244 -8141 15334 -8125
rect 15244 -8175 15260 -8141
rect 15318 -8175 15334 -8141
rect 15244 -8249 15334 -8175
rect 15244 -8283 15260 -8249
rect 15318 -8283 15334 -8249
rect 15244 -8299 15334 -8283
rect 15392 -8141 15482 -8125
rect 15392 -8175 15408 -8141
rect 15466 -8175 15482 -8141
rect 15392 -8249 15482 -8175
rect 15392 -8283 15408 -8249
rect 15466 -8283 15482 -8249
rect 15392 -8299 15482 -8283
rect 15540 -8141 15630 -8125
rect 15540 -8175 15556 -8141
rect 15614 -8175 15630 -8141
rect 15540 -8249 15630 -8175
rect 15540 -8283 15556 -8249
rect 15614 -8283 15630 -8249
rect 15540 -8299 15630 -8283
rect 15688 -8141 15778 -8125
rect 15688 -8175 15704 -8141
rect 15762 -8175 15778 -8141
rect 15688 -8249 15778 -8175
rect 15688 -8283 15704 -8249
rect 15762 -8283 15778 -8249
rect 15688 -8299 15778 -8283
rect 15836 -8141 15926 -8125
rect 15836 -8175 15852 -8141
rect 15910 -8175 15926 -8141
rect 15836 -8249 15926 -8175
rect 15836 -8283 15852 -8249
rect 15910 -8283 15926 -8249
rect 15836 -8299 15926 -8283
rect 15984 -8141 16074 -8125
rect 15984 -8175 16000 -8141
rect 16058 -8175 16074 -8141
rect 15984 -8249 16074 -8175
rect 15984 -8283 16000 -8249
rect 16058 -8283 16074 -8249
rect 15984 -8299 16074 -8283
rect 16132 -8141 16222 -8125
rect 16132 -8175 16148 -8141
rect 16206 -8175 16222 -8141
rect 16132 -8249 16222 -8175
rect 16132 -8283 16148 -8249
rect 16206 -8283 16222 -8249
rect 16132 -8299 16222 -8283
rect 16280 -8141 16370 -8125
rect 16280 -8175 16296 -8141
rect 16354 -8175 16370 -8141
rect 16280 -8249 16370 -8175
rect 16280 -8283 16296 -8249
rect 16354 -8283 16370 -8249
rect 16280 -8299 16370 -8283
rect 16428 -8141 16518 -8125
rect 16428 -8175 16444 -8141
rect 16502 -8175 16518 -8141
rect 16428 -8249 16518 -8175
rect 16428 -8283 16444 -8249
rect 16502 -8283 16518 -8249
rect 16428 -8299 16518 -8283
rect 16576 -8141 16666 -8125
rect 16576 -8175 16592 -8141
rect 16650 -8175 16666 -8141
rect 16576 -8249 16666 -8175
rect 16576 -8283 16592 -8249
rect 16650 -8283 16666 -8249
rect 16576 -8299 16666 -8283
rect 16724 -8141 16814 -8125
rect 16724 -8175 16740 -8141
rect 16798 -8175 16814 -8141
rect 16724 -8249 16814 -8175
rect 16724 -8283 16740 -8249
rect 16798 -8283 16814 -8249
rect 16724 -8299 16814 -8283
rect 16872 -8141 16962 -8125
rect 16872 -8175 16888 -8141
rect 16946 -8175 16962 -8141
rect 16872 -8249 16962 -8175
rect 16872 -8283 16888 -8249
rect 16946 -8283 16962 -8249
rect 16872 -8299 16962 -8283
rect 17020 -8141 17110 -8125
rect 17020 -8175 17036 -8141
rect 17094 -8175 17110 -8141
rect 17020 -8249 17110 -8175
rect 17020 -8283 17036 -8249
rect 17094 -8283 17110 -8249
rect 17020 -8299 17110 -8283
rect 17168 -8141 17258 -8125
rect 17168 -8175 17184 -8141
rect 17242 -8175 17258 -8141
rect 17168 -8249 17258 -8175
rect 17168 -8283 17184 -8249
rect 17242 -8283 17258 -8249
rect 17168 -8299 17258 -8283
rect 17316 -8141 17406 -8125
rect 17316 -8175 17332 -8141
rect 17390 -8175 17406 -8141
rect 17316 -8249 17406 -8175
rect 17316 -8283 17332 -8249
rect 17390 -8283 17406 -8249
rect 17316 -8299 17406 -8283
rect 17464 -8141 17554 -8125
rect 17464 -8175 17480 -8141
rect 17538 -8175 17554 -8141
rect 17464 -8249 17554 -8175
rect 17464 -8283 17480 -8249
rect 17538 -8283 17554 -8249
rect 17464 -8299 17554 -8283
rect 17612 -8141 17702 -8125
rect 17612 -8175 17628 -8141
rect 17686 -8175 17702 -8141
rect 17612 -8249 17702 -8175
rect 17612 -8283 17628 -8249
rect 17686 -8283 17702 -8249
rect 17612 -8299 17702 -8283
rect 17760 -8141 17850 -8125
rect 17760 -8175 17776 -8141
rect 17834 -8175 17850 -8141
rect 17760 -8249 17850 -8175
rect 17760 -8283 17776 -8249
rect 17834 -8283 17850 -8249
rect 17760 -8299 17850 -8283
rect 17908 -8141 17998 -8125
rect 17908 -8175 17924 -8141
rect 17982 -8175 17998 -8141
rect 17908 -8249 17998 -8175
rect 17908 -8283 17924 -8249
rect 17982 -8283 17998 -8249
rect 17908 -8299 17998 -8283
rect 18056 -8141 18146 -8125
rect 18056 -8175 18072 -8141
rect 18130 -8175 18146 -8141
rect 18056 -8249 18146 -8175
rect 18056 -8283 18072 -8249
rect 18130 -8283 18146 -8249
rect 18056 -8299 18146 -8283
rect 18204 -8141 18294 -8125
rect 18204 -8175 18220 -8141
rect 18278 -8175 18294 -8141
rect 18204 -8249 18294 -8175
rect 18204 -8283 18220 -8249
rect 18278 -8283 18294 -8249
rect 18204 -8299 18294 -8283
rect 18352 -8141 18442 -8125
rect 18352 -8175 18368 -8141
rect 18426 -8175 18442 -8141
rect 18352 -8249 18442 -8175
rect 18352 -8283 18368 -8249
rect 18426 -8283 18442 -8249
rect 18352 -8299 18442 -8283
rect 18500 -8141 18590 -8125
rect 18500 -8175 18516 -8141
rect 18574 -8175 18590 -8141
rect 18500 -8249 18590 -8175
rect 18500 -8283 18516 -8249
rect 18574 -8283 18590 -8249
rect 18500 -8299 18590 -8283
rect 18648 -8141 18738 -8125
rect 18648 -8175 18664 -8141
rect 18722 -8175 18738 -8141
rect 18648 -8249 18738 -8175
rect 18648 -8283 18664 -8249
rect 18722 -8283 18738 -8249
rect 18648 -8299 18738 -8283
rect 18796 -8141 18886 -8125
rect 18796 -8175 18812 -8141
rect 18870 -8175 18886 -8141
rect 18796 -8249 18886 -8175
rect 18796 -8283 18812 -8249
rect 18870 -8283 18886 -8249
rect 18796 -8299 18886 -8283
rect 18944 -8141 19034 -8125
rect 18944 -8175 18960 -8141
rect 19018 -8175 19034 -8141
rect 18944 -8249 19034 -8175
rect 18944 -8283 18960 -8249
rect 19018 -8283 19034 -8249
rect 18944 -8299 19034 -8283
rect 19092 -8141 19182 -8125
rect 19092 -8175 19108 -8141
rect 19166 -8175 19182 -8141
rect 19092 -8249 19182 -8175
rect 19092 -8283 19108 -8249
rect 19166 -8283 19182 -8249
rect 19092 -8299 19182 -8283
rect 19240 -8299 19330 -8125
rect 19388 -8299 19478 -8125
rect 19536 -8299 19626 -8125
rect 19684 -8299 19774 -8125
rect 19832 -8141 19922 -8125
rect 19832 -8175 19848 -8141
rect 19906 -8175 19922 -8141
rect 19832 -8249 19922 -8175
rect 19832 -8283 19848 -8249
rect 19906 -8283 19922 -8249
rect 19832 -8299 19922 -8283
rect 19980 -8141 20070 -8125
rect 19980 -8175 19996 -8141
rect 20054 -8175 20070 -8141
rect 19980 -8249 20070 -8175
rect 19980 -8283 19996 -8249
rect 20054 -8283 20070 -8249
rect 19980 -8299 20070 -8283
rect 20128 -8141 20218 -8125
rect 20128 -8175 20144 -8141
rect 20202 -8175 20218 -8141
rect 20128 -8249 20218 -8175
rect 20128 -8283 20144 -8249
rect 20202 -8283 20218 -8249
rect 20128 -8299 20218 -8283
rect 20276 -8141 20366 -8125
rect 20276 -8175 20292 -8141
rect 20350 -8175 20366 -8141
rect 20276 -8249 20366 -8175
rect 20276 -8283 20292 -8249
rect 20350 -8283 20366 -8249
rect 20276 -8299 20366 -8283
rect 20424 -8141 20514 -8125
rect 20424 -8175 20440 -8141
rect 20498 -8175 20514 -8141
rect 20424 -8249 20514 -8175
rect 20424 -8283 20440 -8249
rect 20498 -8283 20514 -8249
rect 20424 -8299 20514 -8283
rect 20572 -8141 20662 -8125
rect 20572 -8175 20588 -8141
rect 20646 -8175 20662 -8141
rect 20572 -8249 20662 -8175
rect 20572 -8283 20588 -8249
rect 20646 -8283 20662 -8249
rect 20572 -8299 20662 -8283
rect 20720 -8141 20810 -8125
rect 20720 -8175 20736 -8141
rect 20794 -8175 20810 -8141
rect 20720 -8249 20810 -8175
rect 20720 -8283 20736 -8249
rect 20794 -8283 20810 -8249
rect 20720 -8299 20810 -8283
rect 20868 -8141 20958 -8125
rect 20868 -8175 20884 -8141
rect 20942 -8175 20958 -8141
rect 20868 -8249 20958 -8175
rect 20868 -8283 20884 -8249
rect 20942 -8283 20958 -8249
rect 20868 -8299 20958 -8283
rect 21016 -8141 21106 -8125
rect 21016 -8175 21032 -8141
rect 21090 -8175 21106 -8141
rect 21016 -8249 21106 -8175
rect 21016 -8283 21032 -8249
rect 21090 -8283 21106 -8249
rect 21016 -8299 21106 -8283
rect 21164 -8141 21254 -8125
rect 21164 -8175 21180 -8141
rect 21238 -8175 21254 -8141
rect 21164 -8249 21254 -8175
rect 21164 -8283 21180 -8249
rect 21238 -8283 21254 -8249
rect 21164 -8299 21254 -8283
rect 21312 -8141 21402 -8125
rect 21312 -8175 21328 -8141
rect 21386 -8175 21402 -8141
rect 21312 -8249 21402 -8175
rect 21312 -8283 21328 -8249
rect 21386 -8283 21402 -8249
rect 21312 -8299 21402 -8283
rect 21460 -8141 21550 -8125
rect 21460 -8175 21476 -8141
rect 21534 -8175 21550 -8141
rect 21460 -8249 21550 -8175
rect 21460 -8283 21476 -8249
rect 21534 -8283 21550 -8249
rect 21460 -8299 21550 -8283
rect 21608 -8141 21698 -8125
rect 21608 -8175 21624 -8141
rect 21682 -8175 21698 -8141
rect 21608 -8249 21698 -8175
rect 21608 -8283 21624 -8249
rect 21682 -8283 21698 -8249
rect 21608 -8299 21698 -8283
rect 21756 -8141 21846 -8125
rect 21756 -8175 21772 -8141
rect 21830 -8175 21846 -8141
rect 21756 -8249 21846 -8175
rect 21756 -8283 21772 -8249
rect 21830 -8283 21846 -8249
rect 21756 -8299 21846 -8283
rect 21904 -8141 21994 -8125
rect 21904 -8175 21920 -8141
rect 21978 -8175 21994 -8141
rect 21904 -8249 21994 -8175
rect 21904 -8283 21920 -8249
rect 21978 -8283 21994 -8249
rect 21904 -8299 21994 -8283
rect 22052 -8141 22142 -8125
rect 22052 -8175 22068 -8141
rect 22126 -8175 22142 -8141
rect 22052 -8249 22142 -8175
rect 22052 -8283 22068 -8249
rect 22126 -8283 22142 -8249
rect 22052 -8299 22142 -8283
rect 22200 -8141 22290 -8125
rect 22200 -8175 22216 -8141
rect 22274 -8175 22290 -8141
rect 22200 -8249 22290 -8175
rect 22200 -8283 22216 -8249
rect 22274 -8283 22290 -8249
rect 22200 -8299 22290 -8283
rect 22348 -8141 22438 -8125
rect 22348 -8175 22364 -8141
rect 22422 -8175 22438 -8141
rect 22348 -8249 22438 -8175
rect 22348 -8283 22364 -8249
rect 22422 -8283 22438 -8249
rect 22348 -8299 22438 -8283
rect 22496 -8141 22586 -8125
rect 22496 -8175 22512 -8141
rect 22570 -8175 22586 -8141
rect 22496 -8249 22586 -8175
rect 22496 -8283 22512 -8249
rect 22570 -8283 22586 -8249
rect 22496 -8299 22586 -8283
rect 22644 -8141 22734 -8125
rect 22644 -8175 22660 -8141
rect 22718 -8175 22734 -8141
rect 22644 -8249 22734 -8175
rect 22644 -8283 22660 -8249
rect 22718 -8283 22734 -8249
rect 22644 -8299 22734 -8283
rect 22792 -8141 22882 -8125
rect 22792 -8175 22808 -8141
rect 22866 -8175 22882 -8141
rect 22792 -8249 22882 -8175
rect 22792 -8283 22808 -8249
rect 22866 -8283 22882 -8249
rect 22792 -8299 22882 -8283
rect 22940 -8141 23030 -8125
rect 22940 -8175 22956 -8141
rect 23014 -8175 23030 -8141
rect 22940 -8249 23030 -8175
rect 22940 -8283 22956 -8249
rect 23014 -8283 23030 -8249
rect 22940 -8299 23030 -8283
rect 23088 -8141 23178 -8125
rect 23088 -8175 23104 -8141
rect 23162 -8175 23178 -8141
rect 23088 -8249 23178 -8175
rect 23088 -8283 23104 -8249
rect 23162 -8283 23178 -8249
rect 23088 -8299 23178 -8283
rect 23236 -8141 23326 -8125
rect 23236 -8175 23252 -8141
rect 23310 -8175 23326 -8141
rect 23236 -8249 23326 -8175
rect 23236 -8283 23252 -8249
rect 23310 -8283 23326 -8249
rect 23236 -8299 23326 -8283
rect 23384 -8141 23474 -8125
rect 23384 -8175 23400 -8141
rect 23458 -8175 23474 -8141
rect 23384 -8249 23474 -8175
rect 23384 -8283 23400 -8249
rect 23458 -8283 23474 -8249
rect 23384 -8299 23474 -8283
rect 23532 -8141 23622 -8125
rect 23532 -8175 23548 -8141
rect 23606 -8175 23622 -8141
rect 23532 -8249 23622 -8175
rect 23532 -8283 23548 -8249
rect 23606 -8283 23622 -8249
rect 23532 -8299 23622 -8283
<< polycont >>
rect 7811 2006 7845 2040
rect 7929 2006 7963 2040
rect 8047 2006 8081 2040
rect 8165 2006 8199 2040
rect 8283 2006 8317 2040
rect 8401 2006 8435 2040
rect 8519 2006 8553 2040
rect 8865 2006 8899 2040
rect 8983 2006 9017 2040
rect 9101 2006 9135 2040
rect 9219 2006 9253 2040
rect 9337 2006 9371 2040
rect 9455 2006 9489 2040
rect 9573 2006 9607 2040
rect 9691 2006 9725 2040
rect 9809 2006 9843 2040
rect 9927 2006 9961 2040
rect 10045 2006 10079 2040
rect 10163 2006 10197 2040
rect 10281 2006 10315 2040
rect 10399 2006 10433 2040
rect 10517 2006 10551 2040
rect 12677 2005 12711 2039
rect 12795 2005 12829 2039
rect 12913 2005 12947 2039
rect 13031 2005 13065 2039
rect 13149 2005 13183 2039
rect 13267 2005 13301 2039
rect 13385 2005 13419 2039
rect 13503 2005 13537 2039
rect 13621 2005 13655 2039
rect 13739 2005 13773 2039
rect 13857 2005 13891 2039
rect 13975 2005 14009 2039
rect 14093 2005 14127 2039
rect 14211 2005 14245 2039
rect 14329 2005 14363 2039
rect 14447 2005 14481 2039
rect 14565 2005 14599 2039
rect 14683 2005 14717 2039
rect 14801 2005 14835 2039
rect 14919 2005 14953 2039
rect 15037 2005 15071 2039
rect 15155 2005 15189 2039
rect 15273 2005 15307 2039
rect 15391 2005 15425 2039
rect 16800 2005 16834 2039
rect 16918 2005 16952 2039
rect 17036 2005 17070 2039
rect 17154 2005 17188 2039
rect 17272 2005 17306 2039
rect 17390 2005 17424 2039
rect 17508 2005 17542 2039
rect 17626 2005 17660 2039
rect 17744 2005 17778 2039
rect 17862 2005 17896 2039
rect 17980 2005 18014 2039
rect 18098 2005 18132 2039
rect 18216 2005 18250 2039
rect 18334 2005 18368 2039
rect 18452 2005 18486 2039
rect 18570 2005 18604 2039
rect 18688 2005 18722 2039
rect 18806 2005 18840 2039
rect 18924 2005 18958 2039
rect 19042 2005 19076 2039
rect 19160 2005 19194 2039
rect 19278 2005 19312 2039
rect 19396 2005 19430 2039
rect 19514 2005 19548 2039
rect 20923 2005 20957 2039
rect 21041 2005 21075 2039
rect 21159 2005 21193 2039
rect 21277 2005 21311 2039
rect 21395 2005 21429 2039
rect 21513 2005 21547 2039
rect 21631 2005 21665 2039
rect 21749 2005 21783 2039
rect 21867 2005 21901 2039
rect 21985 2005 22019 2039
rect 22103 2005 22137 2039
rect 22221 2005 22255 2039
rect 22339 2005 22373 2039
rect 22457 2005 22491 2039
rect 22575 2005 22609 2039
rect 22693 2005 22727 2039
rect 22811 2005 22845 2039
rect 22929 2005 22963 2039
rect 23047 2005 23081 2039
rect 23165 2005 23199 2039
rect 23283 2005 23317 2039
rect 23401 2005 23435 2039
rect 23519 2005 23553 2039
rect 23637 2005 23671 2039
rect 12677 1897 12711 1931
rect 12795 1897 12829 1931
rect 12913 1897 12947 1931
rect 13031 1897 13065 1931
rect 13149 1897 13183 1931
rect 13267 1897 13301 1931
rect 13385 1897 13419 1931
rect 13503 1897 13537 1931
rect 13621 1897 13655 1931
rect 13739 1897 13773 1931
rect 13857 1897 13891 1931
rect 13975 1897 14009 1931
rect 14093 1897 14127 1931
rect 14211 1897 14245 1931
rect 14329 1897 14363 1931
rect 14447 1897 14481 1931
rect 14565 1897 14599 1931
rect 14683 1897 14717 1931
rect 14801 1897 14835 1931
rect 14919 1897 14953 1931
rect 15037 1897 15071 1931
rect 15155 1897 15189 1931
rect 15273 1897 15307 1931
rect 15391 1897 15425 1931
rect 16800 1897 16834 1931
rect 16918 1897 16952 1931
rect 17036 1897 17070 1931
rect 17154 1897 17188 1931
rect 17272 1897 17306 1931
rect 17390 1897 17424 1931
rect 17508 1897 17542 1931
rect 17626 1897 17660 1931
rect 17744 1897 17778 1931
rect 17862 1897 17896 1931
rect 17980 1897 18014 1931
rect 18098 1897 18132 1931
rect 18216 1897 18250 1931
rect 18334 1897 18368 1931
rect 18452 1897 18486 1931
rect 18570 1897 18604 1931
rect 18688 1897 18722 1931
rect 18806 1897 18840 1931
rect 18924 1897 18958 1931
rect 19042 1897 19076 1931
rect 19160 1897 19194 1931
rect 19278 1897 19312 1931
rect 19396 1897 19430 1931
rect 19514 1897 19548 1931
rect 20923 1897 20957 1931
rect 21041 1897 21075 1931
rect 21159 1897 21193 1931
rect 21277 1897 21311 1931
rect 21395 1897 21429 1931
rect 21513 1897 21547 1931
rect 21631 1897 21665 1931
rect 21749 1897 21783 1931
rect 21867 1897 21901 1931
rect 21985 1897 22019 1931
rect 22103 1897 22137 1931
rect 22221 1897 22255 1931
rect 22339 1897 22373 1931
rect 22457 1897 22491 1931
rect 22575 1897 22609 1931
rect 22693 1897 22727 1931
rect 22811 1897 22845 1931
rect 22929 1897 22963 1931
rect 23047 1897 23081 1931
rect 23165 1897 23199 1931
rect 23283 1897 23317 1931
rect 23401 1897 23435 1931
rect 23519 1897 23553 1931
rect 23637 1897 23671 1931
rect 4869 509 4903 543
rect 4869 401 4903 435
rect 4987 509 5021 543
rect 4987 401 5021 435
rect 5105 509 5139 543
rect 5105 401 5139 435
rect 5223 509 5257 543
rect 5223 401 5257 435
rect 5341 509 5375 543
rect 5341 401 5375 435
rect 5459 509 5493 543
rect 5459 401 5493 435
rect 5577 509 5611 543
rect 5577 401 5611 435
rect 5695 509 5729 543
rect 5695 401 5729 435
rect 5813 509 5847 543
rect 5813 401 5847 435
rect 5931 509 5965 543
rect 5931 401 5965 435
rect 6049 509 6083 543
rect 6049 401 6083 435
rect 6167 509 6201 543
rect 6167 401 6201 435
rect 6285 509 6319 543
rect 6285 401 6319 435
rect 6403 509 6437 543
rect 6403 401 6437 435
rect 6521 509 6555 543
rect 6521 401 6555 435
rect 6639 509 6673 543
rect 6639 401 6673 435
rect 6757 509 6791 543
rect 6757 401 6791 435
rect 6875 509 6909 543
rect 6875 401 6909 435
rect 6993 509 7027 543
rect 6993 401 7027 435
rect 7111 509 7145 543
rect 7111 401 7145 435
rect 7229 509 7263 543
rect 7229 401 7263 435
rect 7347 509 7381 543
rect 7347 401 7381 435
rect 7465 509 7499 543
rect 7465 401 7499 435
rect 7583 509 7617 543
rect 7583 401 7617 435
rect 7701 509 7735 543
rect 7701 401 7735 435
rect 7819 509 7853 543
rect 7819 401 7853 435
rect 7937 509 7971 543
rect 7937 401 7971 435
rect 8055 509 8089 543
rect 8055 401 8089 435
rect 8173 509 8207 543
rect 8173 401 8207 435
rect 8291 509 8325 543
rect 8291 401 8325 435
rect 8409 509 8443 543
rect 8409 401 8443 435
rect 8527 509 8561 543
rect 8527 401 8561 435
rect 8645 509 8679 543
rect 8645 401 8679 435
rect 8763 509 8797 543
rect 8763 401 8797 435
rect 8881 509 8915 543
rect 8881 401 8915 435
rect 8999 509 9033 543
rect 8999 401 9033 435
rect 9117 509 9151 543
rect 9117 401 9151 435
rect 9235 509 9269 543
rect 9235 401 9269 435
rect 9353 509 9387 543
rect 9353 401 9387 435
rect 9471 509 9505 543
rect 9471 401 9505 435
rect 9589 509 9623 543
rect 9589 401 9623 435
rect 9707 509 9741 543
rect 9707 401 9741 435
rect 9825 509 9859 543
rect 9825 401 9859 435
rect 9943 509 9977 543
rect 9943 401 9977 435
rect 10061 509 10095 543
rect 10061 401 10095 435
rect 10179 509 10213 543
rect 10179 401 10213 435
rect 10297 509 10331 543
rect 10297 401 10331 435
rect 10415 509 10449 543
rect 10415 401 10449 435
rect 10533 509 10567 543
rect 10533 401 10567 435
rect 10651 509 10685 543
rect 10651 401 10685 435
rect 4869 -1541 4903 -1507
rect 4869 -1649 4903 -1615
rect 4987 -1541 5021 -1507
rect 4987 -1649 5021 -1615
rect 5105 -1541 5139 -1507
rect 5105 -1649 5139 -1615
rect 5223 -1541 5257 -1507
rect 5223 -1649 5257 -1615
rect 5341 -1541 5375 -1507
rect 5341 -1649 5375 -1615
rect 5459 -1541 5493 -1507
rect 5459 -1649 5493 -1615
rect 5577 -1541 5611 -1507
rect 5577 -1649 5611 -1615
rect 5695 -1541 5729 -1507
rect 5695 -1649 5729 -1615
rect 5813 -1541 5847 -1507
rect 5813 -1649 5847 -1615
rect 5931 -1541 5965 -1507
rect 5931 -1649 5965 -1615
rect 6049 -1541 6083 -1507
rect 6049 -1649 6083 -1615
rect 6167 -1541 6201 -1507
rect 6167 -1649 6201 -1615
rect 6285 -1541 6319 -1507
rect 6285 -1649 6319 -1615
rect 6403 -1541 6437 -1507
rect 6403 -1649 6437 -1615
rect 6521 -1541 6555 -1507
rect 6521 -1649 6555 -1615
rect 6639 -1541 6673 -1507
rect 6639 -1649 6673 -1615
rect 6757 -1541 6791 -1507
rect 6757 -1649 6791 -1615
rect 6875 -1541 6909 -1507
rect 6875 -1649 6909 -1615
rect 6993 -1541 7027 -1507
rect 6993 -1649 7027 -1615
rect 7111 -1541 7145 -1507
rect 7111 -1649 7145 -1615
rect 7229 -1541 7263 -1507
rect 7229 -1649 7263 -1615
rect 7347 -1541 7381 -1507
rect 7347 -1649 7381 -1615
rect 7465 -1541 7499 -1507
rect 7465 -1649 7499 -1615
rect 7583 -1541 7617 -1507
rect 7583 -1649 7617 -1615
rect 7701 -1541 7735 -1507
rect 7701 -1649 7735 -1615
rect 7819 -1541 7853 -1507
rect 7819 -1649 7853 -1615
rect 7937 -1541 7971 -1507
rect 7937 -1649 7971 -1615
rect 8055 -1541 8089 -1507
rect 8055 -1649 8089 -1615
rect 8173 -1541 8207 -1507
rect 8173 -1649 8207 -1615
rect 8291 -1541 8325 -1507
rect 8291 -1649 8325 -1615
rect 8409 -1541 8443 -1507
rect 8409 -1649 8443 -1615
rect 8527 -1541 8561 -1507
rect 8527 -1649 8561 -1615
rect 8645 -1541 8679 -1507
rect 8645 -1649 8679 -1615
rect 8763 -1541 8797 -1507
rect 8763 -1649 8797 -1615
rect 8881 -1541 8915 -1507
rect 8881 -1649 8915 -1615
rect 8999 -1541 9033 -1507
rect 8999 -1649 9033 -1615
rect 9117 -1541 9151 -1507
rect 9117 -1649 9151 -1615
rect 9235 -1541 9269 -1507
rect 9235 -1649 9269 -1615
rect 9353 -1541 9387 -1507
rect 9353 -1649 9387 -1615
rect 9471 -1541 9505 -1507
rect 9471 -1649 9505 -1615
rect 9589 -1541 9623 -1507
rect 9589 -1649 9623 -1615
rect 9707 -1541 9741 -1507
rect 9707 -1649 9741 -1615
rect 9825 -1541 9859 -1507
rect 9825 -1649 9859 -1615
rect 9943 -1541 9977 -1507
rect 9943 -1649 9977 -1615
rect 10061 -1541 10095 -1507
rect 10061 -1649 10095 -1615
rect 10179 -1541 10213 -1507
rect 10179 -1649 10213 -1615
rect 10297 -1541 10331 -1507
rect 10297 -1649 10331 -1615
rect 10415 -1541 10449 -1507
rect 10415 -1649 10449 -1615
rect 10533 -1541 10567 -1507
rect 10533 -1649 10567 -1615
rect 10651 -1541 10685 -1507
rect 10651 -1649 10685 -1615
rect 4869 -3591 4903 -3557
rect 4869 -3699 4903 -3665
rect 4987 -3591 5021 -3557
rect 4987 -3699 5021 -3665
rect 5105 -3591 5139 -3557
rect 5105 -3699 5139 -3665
rect 5223 -3591 5257 -3557
rect 5223 -3699 5257 -3665
rect 5341 -3591 5375 -3557
rect 5341 -3699 5375 -3665
rect 5459 -3591 5493 -3557
rect 5459 -3699 5493 -3665
rect 5577 -3591 5611 -3557
rect 5577 -3699 5611 -3665
rect 5695 -3591 5729 -3557
rect 5695 -3699 5729 -3665
rect 5813 -3591 5847 -3557
rect 5813 -3699 5847 -3665
rect 5931 -3591 5965 -3557
rect 5931 -3699 5965 -3665
rect 6049 -3591 6083 -3557
rect 6049 -3699 6083 -3665
rect 6167 -3591 6201 -3557
rect 6167 -3699 6201 -3665
rect 6285 -3591 6319 -3557
rect 6285 -3699 6319 -3665
rect 6403 -3591 6437 -3557
rect 6403 -3699 6437 -3665
rect 6521 -3591 6555 -3557
rect 6521 -3699 6555 -3665
rect 6639 -3591 6673 -3557
rect 6639 -3699 6673 -3665
rect 6757 -3591 6791 -3557
rect 6757 -3699 6791 -3665
rect 6875 -3591 6909 -3557
rect 6875 -3699 6909 -3665
rect 6993 -3591 7027 -3557
rect 6993 -3699 7027 -3665
rect 7111 -3591 7145 -3557
rect 7111 -3699 7145 -3665
rect 7229 -3591 7263 -3557
rect 7229 -3699 7263 -3665
rect 7347 -3591 7381 -3557
rect 7347 -3699 7381 -3665
rect 7465 -3591 7499 -3557
rect 7465 -3699 7499 -3665
rect 7583 -3591 7617 -3557
rect 7583 -3699 7617 -3665
rect 7701 -3591 7735 -3557
rect 7701 -3699 7735 -3665
rect 7819 -3591 7853 -3557
rect 7819 -3699 7853 -3665
rect 7937 -3591 7971 -3557
rect 7937 -3699 7971 -3665
rect 8055 -3591 8089 -3557
rect 8055 -3699 8089 -3665
rect 8173 -3591 8207 -3557
rect 8173 -3699 8207 -3665
rect 8291 -3591 8325 -3557
rect 8291 -3699 8325 -3665
rect 8409 -3591 8443 -3557
rect 8409 -3699 8443 -3665
rect 8527 -3591 8561 -3557
rect 8527 -3699 8561 -3665
rect 8645 -3591 8679 -3557
rect 8645 -3699 8679 -3665
rect 8763 -3591 8797 -3557
rect 8763 -3699 8797 -3665
rect 8881 -3591 8915 -3557
rect 8881 -3699 8915 -3665
rect 8999 -3591 9033 -3557
rect 8999 -3699 9033 -3665
rect 9117 -3591 9151 -3557
rect 9117 -3699 9151 -3665
rect 9235 -3591 9269 -3557
rect 9235 -3699 9269 -3665
rect 9353 -3591 9387 -3557
rect 9353 -3699 9387 -3665
rect 9471 -3591 9505 -3557
rect 9471 -3699 9505 -3665
rect 9589 -3591 9623 -3557
rect 9589 -3699 9623 -3665
rect 9707 -3591 9741 -3557
rect 9707 -3699 9741 -3665
rect 9825 -3591 9859 -3557
rect 9825 -3699 9859 -3665
rect 9943 -3591 9977 -3557
rect 9943 -3699 9977 -3665
rect 10061 -3591 10095 -3557
rect 10061 -3699 10095 -3665
rect 10179 -3591 10213 -3557
rect 10179 -3699 10213 -3665
rect 10297 -3591 10331 -3557
rect 10297 -3699 10331 -3665
rect 10415 -3591 10449 -3557
rect 10415 -3699 10449 -3665
rect 10533 -3591 10567 -3557
rect 10533 -3699 10567 -3665
rect 10651 -3591 10685 -3557
rect 10651 -3699 10685 -3665
rect 4869 -5641 4903 -5607
rect 4869 -5749 4903 -5715
rect 4987 -5641 5021 -5607
rect 4987 -5749 5021 -5715
rect 5105 -5641 5139 -5607
rect 5105 -5749 5139 -5715
rect 5223 -5641 5257 -5607
rect 5223 -5749 5257 -5715
rect 5341 -5641 5375 -5607
rect 5341 -5749 5375 -5715
rect 5459 -5641 5493 -5607
rect 5459 -5749 5493 -5715
rect 5577 -5641 5611 -5607
rect 5577 -5749 5611 -5715
rect 5695 -5641 5729 -5607
rect 5695 -5749 5729 -5715
rect 5813 -5641 5847 -5607
rect 5813 -5749 5847 -5715
rect 5931 -5641 5965 -5607
rect 5931 -5749 5965 -5715
rect 6049 -5641 6083 -5607
rect 6049 -5749 6083 -5715
rect 6167 -5641 6201 -5607
rect 6167 -5749 6201 -5715
rect 6285 -5641 6319 -5607
rect 6285 -5749 6319 -5715
rect 6403 -5641 6437 -5607
rect 6403 -5749 6437 -5715
rect 6521 -5641 6555 -5607
rect 6521 -5749 6555 -5715
rect 6639 -5641 6673 -5607
rect 6639 -5749 6673 -5715
rect 6757 -5641 6791 -5607
rect 6757 -5749 6791 -5715
rect 6875 -5641 6909 -5607
rect 6875 -5749 6909 -5715
rect 6993 -5641 7027 -5607
rect 6993 -5749 7027 -5715
rect 7111 -5641 7145 -5607
rect 7111 -5749 7145 -5715
rect 7229 -5641 7263 -5607
rect 7229 -5749 7263 -5715
rect 7347 -5641 7381 -5607
rect 7347 -5749 7381 -5715
rect 7465 -5641 7499 -5607
rect 7465 -5749 7499 -5715
rect 7583 -5641 7617 -5607
rect 7583 -5749 7617 -5715
rect 7701 -5641 7735 -5607
rect 7701 -5749 7735 -5715
rect 7819 -5641 7853 -5607
rect 7819 -5749 7853 -5715
rect 7937 -5641 7971 -5607
rect 7937 -5749 7971 -5715
rect 8055 -5641 8089 -5607
rect 8055 -5749 8089 -5715
rect 8173 -5641 8207 -5607
rect 8173 -5749 8207 -5715
rect 8291 -5641 8325 -5607
rect 8291 -5749 8325 -5715
rect 8409 -5641 8443 -5607
rect 8409 -5749 8443 -5715
rect 8527 -5641 8561 -5607
rect 8527 -5749 8561 -5715
rect 8645 -5641 8679 -5607
rect 8645 -5749 8679 -5715
rect 8763 -5641 8797 -5607
rect 8763 -5749 8797 -5715
rect 8881 -5641 8915 -5607
rect 8881 -5749 8915 -5715
rect 8999 -5641 9033 -5607
rect 8999 -5749 9033 -5715
rect 9117 -5641 9151 -5607
rect 9117 -5749 9151 -5715
rect 9235 -5641 9269 -5607
rect 9235 -5749 9269 -5715
rect 9353 -5641 9387 -5607
rect 9353 -5749 9387 -5715
rect 9471 -5641 9505 -5607
rect 9471 -5749 9505 -5715
rect 9589 -5641 9623 -5607
rect 9589 -5749 9623 -5715
rect 9707 -5641 9741 -5607
rect 9707 -5749 9741 -5715
rect 9825 -5641 9859 -5607
rect 9825 -5749 9859 -5715
rect 9943 -5641 9977 -5607
rect 9943 -5749 9977 -5715
rect 10061 -5641 10095 -5607
rect 10061 -5749 10095 -5715
rect 10179 -5641 10213 -5607
rect 10179 -5749 10213 -5715
rect 10297 -5641 10331 -5607
rect 10297 -5749 10331 -5715
rect 10415 -5641 10449 -5607
rect 10415 -5749 10449 -5715
rect 10533 -5641 10567 -5607
rect 10533 -5749 10567 -5715
rect 10651 -5641 10685 -5607
rect 10651 -5749 10685 -5715
rect 5935 -7875 5969 -7841
rect 5935 -7983 5969 -7949
rect 6053 -7875 6087 -7841
rect 6053 -7983 6087 -7949
rect 6171 -7875 6205 -7841
rect 6171 -7983 6205 -7949
rect 6289 -7875 6323 -7841
rect 6289 -7983 6323 -7949
rect 6407 -7875 6441 -7841
rect 6407 -7983 6441 -7949
rect 6525 -7875 6559 -7841
rect 6525 -7983 6559 -7949
rect 6643 -7875 6677 -7841
rect 6643 -7983 6677 -7949
rect 6761 -7875 6795 -7841
rect 6761 -7983 6795 -7949
rect 6879 -7875 6913 -7841
rect 6879 -7983 6913 -7949
rect 6997 -7875 7031 -7841
rect 6997 -7983 7031 -7949
rect 7115 -7875 7149 -7841
rect 7115 -7983 7149 -7949
rect 7233 -7875 7267 -7841
rect 7233 -7983 7267 -7949
rect 7351 -7875 7385 -7841
rect 7351 -7983 7385 -7949
rect 7469 -7875 7503 -7841
rect 7469 -7983 7503 -7949
rect 7587 -7875 7621 -7841
rect 7587 -7983 7621 -7949
rect 13188 -8175 13246 -8141
rect 13188 -8283 13246 -8249
rect 13336 -8175 13394 -8141
rect 13336 -8283 13394 -8249
rect 13484 -8175 13542 -8141
rect 13484 -8283 13542 -8249
rect 13632 -8175 13690 -8141
rect 13632 -8283 13690 -8249
rect 13780 -8175 13838 -8141
rect 13780 -8283 13838 -8249
rect 13928 -8175 13986 -8141
rect 13928 -8283 13986 -8249
rect 15556 -8175 15614 -8141
rect 15556 -8283 15614 -8249
rect 15704 -8175 15762 -8141
rect 15704 -8283 15762 -8249
rect 15852 -8175 15910 -8141
rect 15852 -8283 15910 -8249
rect 16000 -8175 16058 -8141
rect 16000 -8283 16058 -8249
rect 16148 -8175 16206 -8141
rect 16148 -8283 16206 -8249
rect 16296 -8175 16354 -8141
rect 16296 -8283 16354 -8249
rect 16444 -8175 16502 -8141
rect 16444 -8283 16502 -8249
rect 16592 -8175 16650 -8141
rect 16592 -8283 16650 -8249
rect 16740 -8175 16798 -8141
rect 16740 -8283 16798 -8249
rect 16888 -8175 16946 -8141
rect 16888 -8283 16946 -8249
rect 17036 -8175 17094 -8141
rect 17036 -8283 17094 -8249
rect 17184 -8175 17242 -8141
rect 17184 -8283 17242 -8249
rect 17332 -8175 17390 -8141
rect 17332 -8283 17390 -8249
rect 17480 -8175 17538 -8141
rect 17480 -8283 17538 -8249
rect 17628 -8175 17686 -8141
rect 17628 -8283 17686 -8249
rect 17776 -8175 17834 -8141
rect 17776 -8283 17834 -8249
rect 17924 -8175 17982 -8141
rect 17924 -8283 17982 -8249
rect 18072 -8175 18130 -8141
rect 18072 -8283 18130 -8249
rect 18220 -8175 18278 -8141
rect 18220 -8283 18278 -8249
rect 18368 -8175 18426 -8141
rect 18368 -8283 18426 -8249
<< locali >>
rect 4730 3118 4768 3152
rect 12420 3117 12458 3151
rect 18468 3117 18597 3151
rect 4760 3030 4768 3064
rect 10778 3030 10808 3064
rect 12450 3029 12458 3063
rect 18468 3029 18597 3063
rect 24607 3029 24637 3063
rect 4760 2942 4768 2976
rect 10778 2942 10808 2976
rect 12450 2941 12458 2975
rect 18468 2941 18597 2975
rect 24607 2941 24637 2975
rect 15693 2653 15731 2687
rect 15765 2653 15803 2687
rect 15837 2653 15875 2687
rect 15909 2653 15947 2687
rect 15981 2653 16019 2687
rect 16053 2653 16091 2687
rect 16125 2653 16163 2687
rect 16197 2653 16235 2687
rect 16269 2653 16307 2687
rect 16341 2653 16379 2687
rect 15693 2579 15731 2613
rect 15765 2579 15803 2613
rect 15837 2579 15875 2613
rect 15909 2579 15947 2613
rect 15981 2579 16019 2613
rect 16053 2579 16091 2613
rect 16125 2579 16163 2613
rect 16197 2579 16235 2613
rect 16269 2579 16307 2613
rect 16341 2579 16379 2613
rect 15693 2505 15731 2539
rect 15765 2505 15803 2539
rect 15837 2505 15875 2539
rect 15909 2505 15947 2539
rect 15981 2505 16019 2539
rect 16053 2505 16091 2539
rect 16125 2505 16163 2539
rect 16197 2505 16235 2539
rect 16269 2505 16307 2539
rect 16341 2505 16379 2539
rect 15693 2431 15731 2465
rect 15765 2431 15803 2465
rect 15837 2431 15875 2465
rect 15909 2431 15947 2465
rect 15981 2431 16019 2465
rect 16053 2431 16091 2465
rect 16125 2431 16163 2465
rect 16197 2431 16235 2465
rect 16269 2431 16307 2465
rect 16341 2431 16379 2465
rect 15693 2357 15731 2391
rect 15765 2357 15803 2391
rect 15837 2357 15875 2391
rect 15909 2357 15947 2391
rect 15981 2357 16019 2391
rect 16053 2357 16091 2391
rect 16125 2357 16163 2391
rect 16197 2357 16235 2391
rect 16269 2357 16307 2391
rect 16341 2357 16379 2391
rect 15693 2283 15731 2317
rect 15765 2283 15803 2317
rect 15837 2283 15875 2317
rect 15909 2283 15947 2317
rect 15981 2283 16019 2317
rect 16053 2283 16091 2317
rect 16125 2283 16163 2317
rect 16197 2283 16235 2317
rect 16269 2283 16307 2317
rect 16341 2283 16379 2317
rect 15693 2209 15731 2243
rect 15765 2209 15803 2243
rect 15837 2209 15875 2243
rect 15909 2209 15947 2243
rect 15981 2209 16019 2243
rect 16053 2209 16091 2243
rect 16125 2209 16163 2243
rect 16197 2209 16235 2243
rect 16269 2209 16307 2243
rect 16341 2209 16379 2243
rect 15693 2135 15731 2169
rect 15765 2135 15803 2169
rect 15837 2135 15875 2169
rect 15909 2135 15947 2169
rect 15981 2135 16019 2169
rect 16053 2135 16091 2169
rect 16125 2135 16163 2169
rect 16197 2135 16235 2169
rect 16269 2135 16307 2169
rect 16341 2135 16379 2169
rect 19816 2653 19854 2687
rect 19888 2653 19926 2687
rect 19960 2653 19998 2687
rect 20032 2653 20070 2687
rect 20104 2653 20142 2687
rect 20176 2653 20214 2687
rect 20248 2653 20286 2687
rect 20320 2653 20358 2687
rect 20392 2653 20430 2687
rect 20464 2653 20502 2687
rect 19816 2579 19854 2613
rect 19888 2579 19926 2613
rect 19960 2579 19998 2613
rect 20032 2579 20070 2613
rect 20104 2579 20142 2613
rect 20176 2579 20214 2613
rect 20248 2579 20286 2613
rect 20320 2579 20358 2613
rect 20392 2579 20430 2613
rect 20464 2579 20502 2613
rect 19816 2505 19854 2539
rect 19888 2505 19926 2539
rect 19960 2505 19998 2539
rect 20032 2505 20070 2539
rect 20104 2505 20142 2539
rect 20176 2505 20214 2539
rect 20248 2505 20286 2539
rect 20320 2505 20358 2539
rect 20392 2505 20430 2539
rect 20464 2505 20502 2539
rect 19816 2431 19854 2465
rect 19888 2431 19926 2465
rect 19960 2431 19998 2465
rect 20032 2431 20070 2465
rect 20104 2431 20142 2465
rect 20176 2431 20214 2465
rect 20248 2431 20286 2465
rect 20320 2431 20358 2465
rect 20392 2431 20430 2465
rect 20464 2431 20502 2465
rect 19816 2357 19854 2391
rect 19888 2357 19926 2391
rect 19960 2357 19998 2391
rect 20032 2357 20070 2391
rect 20104 2357 20142 2391
rect 20176 2357 20214 2391
rect 20248 2357 20286 2391
rect 20320 2357 20358 2391
rect 20392 2357 20430 2391
rect 20464 2357 20502 2391
rect 19816 2283 19854 2317
rect 19888 2283 19926 2317
rect 19960 2283 19998 2317
rect 20032 2283 20070 2317
rect 20104 2283 20142 2317
rect 20176 2283 20214 2317
rect 20248 2283 20286 2317
rect 20320 2283 20358 2317
rect 20392 2283 20430 2317
rect 20464 2283 20502 2317
rect 19816 2209 19854 2243
rect 19888 2209 19926 2243
rect 19960 2209 19998 2243
rect 20032 2209 20070 2243
rect 20104 2209 20142 2243
rect 20176 2209 20214 2243
rect 20248 2209 20286 2243
rect 20320 2209 20358 2243
rect 20392 2209 20430 2243
rect 20464 2209 20502 2243
rect 19816 2135 19854 2169
rect 19888 2135 19926 2169
rect 19960 2135 19998 2169
rect 20032 2135 20070 2169
rect 20104 2135 20142 2169
rect 20176 2135 20214 2169
rect 20248 2135 20286 2169
rect 20320 2135 20358 2169
rect 20392 2135 20430 2169
rect 20464 2135 20502 2169
rect 23939 2653 23977 2687
rect 24011 2653 24049 2687
rect 24083 2653 24121 2687
rect 24155 2653 24193 2687
rect 24227 2653 24265 2687
rect 24299 2653 24337 2687
rect 24371 2653 24409 2687
rect 24443 2653 24481 2687
rect 24515 2653 24553 2687
rect 24587 2653 24625 2687
rect 23939 2579 23977 2613
rect 24011 2579 24049 2613
rect 24083 2579 24121 2613
rect 24155 2579 24193 2613
rect 24227 2579 24265 2613
rect 24299 2579 24337 2613
rect 24371 2579 24409 2613
rect 24443 2579 24481 2613
rect 24515 2579 24553 2613
rect 24587 2579 24625 2613
rect 23939 2505 23977 2539
rect 24011 2505 24049 2539
rect 24083 2505 24121 2539
rect 24155 2505 24193 2539
rect 24227 2505 24265 2539
rect 24299 2505 24337 2539
rect 24371 2505 24409 2539
rect 24443 2505 24481 2539
rect 24515 2505 24553 2539
rect 24587 2505 24625 2539
rect 23939 2431 23977 2465
rect 24011 2431 24049 2465
rect 24083 2431 24121 2465
rect 24155 2431 24193 2465
rect 24227 2431 24265 2465
rect 24299 2431 24337 2465
rect 24371 2431 24409 2465
rect 24443 2431 24481 2465
rect 24515 2431 24553 2465
rect 24587 2431 24625 2465
rect 23939 2357 23977 2391
rect 24011 2357 24049 2391
rect 24083 2357 24121 2391
rect 24155 2357 24193 2391
rect 24227 2357 24265 2391
rect 24299 2357 24337 2391
rect 24371 2357 24409 2391
rect 24443 2357 24481 2391
rect 24515 2357 24553 2391
rect 24587 2357 24625 2391
rect 23939 2283 23977 2317
rect 24011 2283 24049 2317
rect 24083 2283 24121 2317
rect 24155 2283 24193 2317
rect 24227 2283 24265 2317
rect 24299 2283 24337 2317
rect 24371 2283 24409 2317
rect 24443 2283 24481 2317
rect 24515 2283 24553 2317
rect 24587 2283 24625 2317
rect 23939 2209 23977 2243
rect 24011 2209 24049 2243
rect 24083 2209 24121 2243
rect 24155 2209 24193 2243
rect 24227 2209 24265 2243
rect 24299 2209 24337 2243
rect 24371 2209 24409 2243
rect 24443 2209 24481 2243
rect 24515 2209 24553 2243
rect 24587 2209 24625 2243
rect 23939 2135 23977 2169
rect 24011 2135 24049 2169
rect 24083 2135 24121 2169
rect 24155 2135 24193 2169
rect 24227 2135 24265 2169
rect 24299 2135 24337 2169
rect 24371 2135 24409 2169
rect 24443 2135 24481 2169
rect 24515 2135 24553 2169
rect 24587 2135 24625 2169
rect 15693 2061 15731 2095
rect 15765 2061 15803 2095
rect 15837 2061 15875 2095
rect 15909 2061 15947 2095
rect 15981 2061 16019 2095
rect 16053 2061 16091 2095
rect 16125 2061 16163 2095
rect 16197 2061 16235 2095
rect 16269 2061 16307 2095
rect 16341 2061 16379 2095
rect 19816 2061 19854 2095
rect 19888 2061 19926 2095
rect 19960 2061 19998 2095
rect 20032 2061 20070 2095
rect 20104 2061 20142 2095
rect 20176 2061 20214 2095
rect 20248 2061 20286 2095
rect 20320 2061 20358 2095
rect 20392 2061 20430 2095
rect 20464 2061 20502 2095
rect 23939 2061 23977 2095
rect 24011 2061 24049 2095
rect 24083 2061 24121 2095
rect 24155 2061 24193 2095
rect 24227 2061 24265 2095
rect 24299 2061 24337 2095
rect 24371 2061 24409 2095
rect 24443 2061 24481 2095
rect 24515 2061 24553 2095
rect 24587 2061 24625 2095
rect 7795 2006 7811 2040
rect 7845 2006 7861 2040
rect 7913 2006 7929 2040
rect 7963 2006 7979 2040
rect 8031 2006 8047 2040
rect 8081 2006 8097 2040
rect 8149 2006 8165 2040
rect 8199 2006 8215 2040
rect 8267 2006 8283 2040
rect 8317 2006 8333 2040
rect 8385 2006 8401 2040
rect 8435 2006 8451 2040
rect 8503 2006 8519 2040
rect 8553 2006 8569 2040
rect 8849 2006 8865 2040
rect 8899 2006 8915 2040
rect 8967 2006 8983 2040
rect 9017 2006 9033 2040
rect 9085 2006 9101 2040
rect 9135 2006 9151 2040
rect 9203 2006 9219 2040
rect 9253 2006 9269 2040
rect 9321 2006 9337 2040
rect 9371 2006 9387 2040
rect 9439 2006 9455 2040
rect 9489 2006 9505 2040
rect 9557 2006 9573 2040
rect 9607 2006 9623 2040
rect 9675 2006 9691 2040
rect 9725 2006 9741 2040
rect 9793 2006 9809 2040
rect 9843 2006 9859 2040
rect 9911 2006 9927 2040
rect 9961 2006 9977 2040
rect 10029 2006 10045 2040
rect 10079 2006 10095 2040
rect 10147 2006 10163 2040
rect 10197 2006 10213 2040
rect 10265 2006 10281 2040
rect 10315 2006 10331 2040
rect 10383 2006 10399 2040
rect 10433 2006 10449 2040
rect 10501 2006 10517 2040
rect 10551 2006 10567 2040
rect 12665 2005 12677 2039
rect 12711 2005 12723 2039
rect 12779 2005 12795 2039
rect 12829 2005 12845 2039
rect 12897 2005 12913 2039
rect 12947 2005 12963 2039
rect 13015 2005 13031 2039
rect 13065 2005 13081 2039
rect 13133 2005 13149 2039
rect 13183 2005 13199 2039
rect 13251 2005 13267 2039
rect 13301 2005 13317 2039
rect 13369 2005 13385 2039
rect 13419 2005 13435 2039
rect 13487 2005 13503 2039
rect 13537 2005 13553 2039
rect 13605 2005 13621 2039
rect 13655 2005 13671 2039
rect 13723 2005 13739 2039
rect 13773 2005 13789 2039
rect 13841 2005 13857 2039
rect 13891 2005 13907 2039
rect 13959 2005 13975 2039
rect 14009 2005 14025 2039
rect 14077 2005 14093 2039
rect 14127 2005 14143 2039
rect 14195 2005 14211 2039
rect 14245 2005 14261 2039
rect 14313 2005 14329 2039
rect 14363 2005 14379 2039
rect 14431 2005 14447 2039
rect 14481 2005 14497 2039
rect 14549 2005 14565 2039
rect 14599 2005 14615 2039
rect 14667 2005 14683 2039
rect 14717 2005 14733 2039
rect 14785 2005 14801 2039
rect 14835 2005 14851 2039
rect 14903 2005 14919 2039
rect 14953 2005 14969 2039
rect 15021 2005 15037 2039
rect 15071 2005 15087 2039
rect 15139 2005 15155 2039
rect 15189 2005 15205 2039
rect 15257 2005 15273 2039
rect 15307 2005 15323 2039
rect 15375 2005 15391 2039
rect 15425 2005 15441 2039
rect 15693 1987 15731 2021
rect 15765 1987 15803 2021
rect 15837 1987 15875 2021
rect 15909 1987 15947 2021
rect 15981 1987 16019 2021
rect 16053 1987 16091 2021
rect 16125 1987 16163 2021
rect 16197 1987 16235 2021
rect 16269 1987 16307 2021
rect 16341 1987 16379 2021
rect 16788 2005 16800 2039
rect 16834 2005 16846 2039
rect 16902 2005 16918 2039
rect 16952 2005 16968 2039
rect 17020 2005 17036 2039
rect 17070 2005 17086 2039
rect 17138 2005 17154 2039
rect 17188 2005 17204 2039
rect 17256 2005 17272 2039
rect 17306 2005 17322 2039
rect 17374 2005 17390 2039
rect 17424 2005 17440 2039
rect 17492 2005 17508 2039
rect 17542 2005 17558 2039
rect 17610 2005 17626 2039
rect 17660 2005 17676 2039
rect 17728 2005 17744 2039
rect 17778 2005 17794 2039
rect 17846 2005 17862 2039
rect 17896 2005 17912 2039
rect 17964 2005 17980 2039
rect 18014 2005 18030 2039
rect 18082 2005 18098 2039
rect 18132 2005 18148 2039
rect 18200 2005 18216 2039
rect 18250 2005 18266 2039
rect 18318 2005 18334 2039
rect 18368 2005 18384 2039
rect 18436 2005 18452 2039
rect 18486 2005 18502 2039
rect 18554 2005 18570 2039
rect 18604 2005 18620 2039
rect 18672 2005 18688 2039
rect 18722 2005 18738 2039
rect 18790 2005 18806 2039
rect 18840 2005 18856 2039
rect 18908 2005 18924 2039
rect 18958 2005 18974 2039
rect 19026 2005 19042 2039
rect 19076 2005 19092 2039
rect 19144 2005 19160 2039
rect 19194 2005 19210 2039
rect 19262 2005 19278 2039
rect 19312 2005 19328 2039
rect 19380 2005 19396 2039
rect 19430 2005 19446 2039
rect 19498 2005 19514 2039
rect 19548 2005 19564 2039
rect 19816 1987 19854 2021
rect 19888 1987 19926 2021
rect 19960 1987 19998 2021
rect 20032 1987 20070 2021
rect 20104 1987 20142 2021
rect 20176 1987 20214 2021
rect 20248 1987 20286 2021
rect 20320 1987 20358 2021
rect 20392 1987 20430 2021
rect 20464 1987 20502 2021
rect 20911 2005 20923 2039
rect 20957 2005 20969 2039
rect 21025 2005 21041 2039
rect 21075 2005 21091 2039
rect 21143 2005 21159 2039
rect 21193 2005 21209 2039
rect 21261 2005 21277 2039
rect 21311 2005 21327 2039
rect 21379 2005 21395 2039
rect 21429 2005 21445 2039
rect 21497 2005 21513 2039
rect 21547 2005 21563 2039
rect 21615 2005 21631 2039
rect 21665 2005 21681 2039
rect 21733 2005 21749 2039
rect 21783 2005 21799 2039
rect 21851 2005 21867 2039
rect 21901 2005 21917 2039
rect 21969 2005 21985 2039
rect 22019 2005 22035 2039
rect 22087 2005 22103 2039
rect 22137 2005 22153 2039
rect 22205 2005 22221 2039
rect 22255 2005 22271 2039
rect 22323 2005 22339 2039
rect 22373 2005 22389 2039
rect 22441 2005 22457 2039
rect 22491 2005 22507 2039
rect 22559 2005 22575 2039
rect 22609 2005 22625 2039
rect 22677 2005 22693 2039
rect 22727 2005 22743 2039
rect 22795 2005 22811 2039
rect 22845 2005 22861 2039
rect 22913 2005 22929 2039
rect 22963 2005 22979 2039
rect 23031 2005 23047 2039
rect 23081 2005 23097 2039
rect 23149 2005 23165 2039
rect 23199 2005 23215 2039
rect 23267 2005 23283 2039
rect 23317 2005 23333 2039
rect 23385 2005 23401 2039
rect 23435 2005 23451 2039
rect 23503 2005 23519 2039
rect 23553 2005 23569 2039
rect 23621 2005 23637 2039
rect 23671 2005 23687 2039
rect 23939 1987 23977 2021
rect 24011 1987 24049 2021
rect 24083 1987 24121 2021
rect 24155 1987 24193 2021
rect 24227 1987 24265 2021
rect 24299 1987 24337 2021
rect 24371 1987 24409 2021
rect 24443 1987 24481 2021
rect 24515 1987 24553 2021
rect 24587 1987 24625 2021
rect 12665 1897 12677 1931
rect 12711 1897 12723 1931
rect 12779 1897 12795 1931
rect 12829 1897 12845 1931
rect 12897 1897 12913 1931
rect 12947 1897 12963 1931
rect 13015 1897 13031 1931
rect 13065 1897 13081 1931
rect 13133 1897 13149 1931
rect 13183 1897 13199 1931
rect 13251 1897 13267 1931
rect 13301 1897 13317 1931
rect 13369 1897 13385 1931
rect 13419 1897 13435 1931
rect 13487 1897 13503 1931
rect 13537 1897 13553 1931
rect 13605 1897 13621 1931
rect 13655 1897 13671 1931
rect 13723 1897 13739 1931
rect 13773 1897 13789 1931
rect 13841 1897 13857 1931
rect 13891 1897 13907 1931
rect 13959 1897 13975 1931
rect 14009 1897 14025 1931
rect 14077 1897 14093 1931
rect 14127 1897 14143 1931
rect 14195 1897 14211 1931
rect 14245 1897 14261 1931
rect 14313 1897 14329 1931
rect 14363 1897 14379 1931
rect 14431 1897 14447 1931
rect 14481 1897 14497 1931
rect 14549 1897 14565 1931
rect 14599 1897 14615 1931
rect 14667 1897 14683 1931
rect 14717 1897 14733 1931
rect 14785 1897 14801 1931
rect 14835 1897 14851 1931
rect 14903 1897 14919 1931
rect 14953 1897 14969 1931
rect 15021 1897 15037 1931
rect 15071 1897 15087 1931
rect 15139 1897 15155 1931
rect 15189 1897 15205 1931
rect 15257 1897 15273 1931
rect 15307 1897 15323 1931
rect 15375 1897 15391 1931
rect 15425 1897 15441 1931
rect 15693 1913 15731 1947
rect 15765 1913 15803 1947
rect 15837 1913 15875 1947
rect 15909 1913 15947 1947
rect 15981 1913 16019 1947
rect 16053 1913 16091 1947
rect 16125 1913 16163 1947
rect 16197 1913 16235 1947
rect 16269 1913 16307 1947
rect 16341 1913 16379 1947
rect 16788 1897 16800 1931
rect 16834 1897 16846 1931
rect 16902 1897 16918 1931
rect 16952 1897 16968 1931
rect 17020 1897 17036 1931
rect 17070 1897 17086 1931
rect 17138 1897 17154 1931
rect 17188 1897 17204 1931
rect 17256 1897 17272 1931
rect 17306 1897 17322 1931
rect 17374 1897 17390 1931
rect 17424 1897 17440 1931
rect 17492 1897 17508 1931
rect 17542 1897 17558 1931
rect 17610 1897 17626 1931
rect 17660 1897 17676 1931
rect 17728 1897 17744 1931
rect 17778 1897 17794 1931
rect 17846 1897 17862 1931
rect 17896 1897 17912 1931
rect 17964 1897 17980 1931
rect 18014 1897 18030 1931
rect 18082 1897 18098 1931
rect 18132 1897 18148 1931
rect 18200 1897 18216 1931
rect 18250 1897 18266 1931
rect 18318 1897 18334 1931
rect 18368 1897 18384 1931
rect 18436 1897 18452 1931
rect 18486 1897 18502 1931
rect 18554 1897 18570 1931
rect 18604 1897 18620 1931
rect 18672 1897 18688 1931
rect 18722 1897 18738 1931
rect 18790 1897 18806 1931
rect 18840 1897 18856 1931
rect 18908 1897 18924 1931
rect 18958 1897 18974 1931
rect 19026 1897 19042 1931
rect 19076 1897 19092 1931
rect 19144 1897 19160 1931
rect 19194 1897 19210 1931
rect 19262 1897 19278 1931
rect 19312 1897 19328 1931
rect 19380 1897 19396 1931
rect 19430 1897 19446 1931
rect 19498 1897 19514 1931
rect 19548 1897 19564 1931
rect 19816 1913 19854 1947
rect 19888 1913 19926 1947
rect 19960 1913 19998 1947
rect 20032 1913 20070 1947
rect 20104 1913 20142 1947
rect 20176 1913 20214 1947
rect 20248 1913 20286 1947
rect 20320 1913 20358 1947
rect 20392 1913 20430 1947
rect 20464 1913 20502 1947
rect 20911 1897 20923 1931
rect 20957 1897 20969 1931
rect 21025 1897 21041 1931
rect 21075 1897 21091 1931
rect 21143 1897 21159 1931
rect 21193 1897 21209 1931
rect 21261 1897 21277 1931
rect 21311 1897 21327 1931
rect 21379 1897 21395 1931
rect 21429 1897 21445 1931
rect 21497 1897 21513 1931
rect 21547 1897 21563 1931
rect 21615 1897 21631 1931
rect 21665 1897 21681 1931
rect 21733 1897 21749 1931
rect 21783 1897 21799 1931
rect 21851 1897 21867 1931
rect 21901 1897 21917 1931
rect 21969 1897 21985 1931
rect 22019 1897 22035 1931
rect 22087 1897 22103 1931
rect 22137 1897 22153 1931
rect 22205 1897 22221 1931
rect 22255 1897 22271 1931
rect 22323 1897 22339 1931
rect 22373 1897 22389 1931
rect 22441 1897 22457 1931
rect 22491 1897 22507 1931
rect 22559 1897 22575 1931
rect 22609 1897 22625 1931
rect 22677 1897 22693 1931
rect 22727 1897 22743 1931
rect 22795 1897 22811 1931
rect 22845 1897 22861 1931
rect 22913 1897 22929 1931
rect 22963 1897 22979 1931
rect 23031 1897 23047 1931
rect 23081 1897 23097 1931
rect 23149 1897 23165 1931
rect 23199 1897 23215 1931
rect 23267 1897 23283 1931
rect 23317 1897 23333 1931
rect 23385 1897 23401 1931
rect 23435 1897 23451 1931
rect 23503 1897 23519 1931
rect 23553 1897 23569 1931
rect 23621 1897 23637 1931
rect 23671 1897 23687 1931
rect 23939 1913 23977 1947
rect 24011 1913 24049 1947
rect 24083 1913 24121 1947
rect 24155 1913 24193 1947
rect 24227 1913 24265 1947
rect 24299 1913 24337 1947
rect 24371 1913 24409 1947
rect 24443 1913 24481 1947
rect 24515 1913 24553 1947
rect 24587 1913 24625 1947
rect 15693 1839 15731 1873
rect 15765 1839 15803 1873
rect 15837 1839 15875 1873
rect 15909 1839 15947 1873
rect 15981 1839 16019 1873
rect 16053 1839 16091 1873
rect 16125 1839 16163 1873
rect 16197 1839 16235 1873
rect 16269 1839 16307 1873
rect 16341 1839 16379 1873
rect 19816 1839 19854 1873
rect 19888 1839 19926 1873
rect 19960 1839 19998 1873
rect 20032 1839 20070 1873
rect 20104 1839 20142 1873
rect 20176 1839 20214 1873
rect 20248 1839 20286 1873
rect 20320 1839 20358 1873
rect 20392 1839 20430 1873
rect 20464 1839 20502 1873
rect 23939 1839 23977 1873
rect 24011 1839 24049 1873
rect 24083 1839 24121 1873
rect 24155 1839 24193 1873
rect 24227 1839 24265 1873
rect 24299 1839 24337 1873
rect 24371 1839 24409 1873
rect 24443 1839 24481 1873
rect 24515 1839 24553 1873
rect 24587 1839 24625 1873
rect 4703 1515 4836 1549
rect 4710 1429 4792 1461
rect 4718 1427 4792 1429
rect 10762 1427 10778 1461
rect 4696 1339 4792 1373
rect 10762 1339 10858 1373
rect 4696 1277 4730 1339
rect 10824 1277 10858 1339
rect 4810 1178 4844 1194
rect 4810 586 4844 602
rect 4928 1178 4962 1194
rect 4928 586 4962 602
rect 5046 1178 5080 1194
rect 5046 586 5080 602
rect 5164 1178 5198 1194
rect 5164 586 5198 602
rect 5282 1178 5316 1194
rect 5282 586 5316 602
rect 5400 1178 5434 1194
rect 5400 586 5434 602
rect 5518 1178 5552 1194
rect 5518 586 5552 602
rect 5636 1178 5670 1194
rect 5636 586 5670 602
rect 5754 1178 5788 1194
rect 5754 586 5788 602
rect 5872 1178 5906 1194
rect 5872 586 5906 602
rect 5990 1178 6024 1194
rect 5990 586 6024 602
rect 6108 1178 6142 1194
rect 6108 586 6142 602
rect 6226 1178 6260 1194
rect 6226 586 6260 602
rect 6344 1178 6378 1194
rect 6344 586 6378 602
rect 6462 1178 6496 1194
rect 6462 586 6496 602
rect 6580 1178 6614 1194
rect 6580 586 6614 602
rect 6698 1178 6732 1194
rect 6698 586 6732 602
rect 6816 1178 6850 1194
rect 6816 586 6850 602
rect 6934 1178 6968 1194
rect 6934 586 6968 602
rect 7052 1178 7086 1194
rect 7052 586 7086 602
rect 7170 1178 7204 1194
rect 7170 586 7204 602
rect 7288 1178 7322 1194
rect 7288 586 7322 602
rect 7406 1178 7440 1194
rect 7406 586 7440 602
rect 7524 1178 7558 1194
rect 7524 586 7558 602
rect 7642 1178 7676 1194
rect 7642 586 7676 602
rect 7760 1178 7794 1194
rect 7760 586 7794 602
rect 7878 1178 7912 1194
rect 7878 586 7912 602
rect 7996 1178 8030 1194
rect 7996 586 8030 602
rect 8114 1178 8148 1194
rect 8114 586 8148 602
rect 8232 1178 8266 1194
rect 8232 586 8266 602
rect 8350 1178 8384 1194
rect 8350 586 8384 602
rect 8468 1178 8502 1194
rect 8468 586 8502 602
rect 8586 1178 8620 1194
rect 8586 586 8620 602
rect 8704 1178 8738 1194
rect 8704 586 8738 602
rect 8822 1178 8856 1194
rect 8822 586 8856 602
rect 8940 1178 8974 1194
rect 8940 586 8974 602
rect 9058 1178 9092 1194
rect 9058 586 9092 602
rect 9176 1178 9210 1194
rect 9176 586 9210 602
rect 9294 1178 9328 1194
rect 9294 586 9328 602
rect 9412 1178 9446 1194
rect 9412 586 9446 602
rect 9530 1178 9564 1194
rect 9530 586 9564 602
rect 9648 1178 9682 1194
rect 9648 586 9682 602
rect 9766 1178 9800 1194
rect 9766 586 9800 602
rect 9884 1178 9918 1194
rect 9884 586 9918 602
rect 10002 1178 10036 1194
rect 10002 586 10036 602
rect 10120 1178 10154 1194
rect 10120 586 10154 602
rect 10238 1178 10272 1194
rect 10238 586 10272 602
rect 10356 1178 10390 1194
rect 10356 586 10390 602
rect 10474 1178 10508 1194
rect 10474 586 10508 602
rect 10592 1178 10626 1194
rect 10592 586 10626 602
rect 10710 1178 10744 1194
rect 10710 586 10744 602
rect 4853 509 4869 543
rect 4903 509 4919 543
rect 4971 509 4987 543
rect 5021 509 5037 543
rect 5089 509 5105 543
rect 5139 509 5155 543
rect 5207 509 5223 543
rect 5257 509 5273 543
rect 5325 509 5341 543
rect 5375 509 5391 543
rect 5443 509 5459 543
rect 5493 509 5509 543
rect 5561 509 5577 543
rect 5611 509 5627 543
rect 5679 509 5695 543
rect 5729 509 5745 543
rect 5797 509 5813 543
rect 5847 509 5863 543
rect 5915 509 5931 543
rect 5965 509 5981 543
rect 6033 509 6049 543
rect 6083 509 6099 543
rect 6151 509 6167 543
rect 6201 509 6217 543
rect 6269 509 6285 543
rect 6319 509 6335 543
rect 6387 509 6403 543
rect 6437 509 6453 543
rect 6505 509 6521 543
rect 6555 509 6571 543
rect 6623 509 6639 543
rect 6673 509 6689 543
rect 6741 509 6757 543
rect 6791 509 6807 543
rect 6859 509 6875 543
rect 6909 509 6925 543
rect 6977 509 6993 543
rect 7027 509 7043 543
rect 7095 509 7111 543
rect 7145 509 7161 543
rect 7213 509 7229 543
rect 7263 509 7279 543
rect 7331 509 7347 543
rect 7381 509 7397 543
rect 7449 509 7465 543
rect 7499 509 7515 543
rect 7567 509 7583 543
rect 7617 509 7633 543
rect 7685 509 7701 543
rect 7735 509 7751 543
rect 7803 509 7819 543
rect 7853 509 7869 543
rect 7921 509 7937 543
rect 7971 509 7987 543
rect 8039 509 8055 543
rect 8089 509 8105 543
rect 8157 509 8173 543
rect 8207 509 8223 543
rect 8275 509 8291 543
rect 8325 509 8341 543
rect 8393 509 8409 543
rect 8443 509 8459 543
rect 8511 509 8527 543
rect 8561 509 8577 543
rect 8629 509 8645 543
rect 8679 509 8695 543
rect 8747 509 8763 543
rect 8797 509 8813 543
rect 8865 509 8881 543
rect 8915 509 8931 543
rect 8983 509 8999 543
rect 9033 509 9049 543
rect 9101 509 9117 543
rect 9151 509 9167 543
rect 9219 509 9235 543
rect 9269 509 9285 543
rect 9337 509 9353 543
rect 9387 509 9403 543
rect 9455 509 9471 543
rect 9505 509 9521 543
rect 9573 509 9589 543
rect 9623 509 9639 543
rect 9691 509 9707 543
rect 9741 509 9757 543
rect 9809 509 9825 543
rect 9859 509 9875 543
rect 9927 509 9943 543
rect 9977 509 9993 543
rect 10045 509 10061 543
rect 10095 509 10111 543
rect 10163 509 10179 543
rect 10213 509 10229 543
rect 10281 509 10297 543
rect 10331 509 10347 543
rect 10399 509 10415 543
rect 10449 509 10465 543
rect 10517 509 10533 543
rect 10567 509 10583 543
rect 10635 509 10651 543
rect 10685 509 10701 543
rect 4853 401 4869 435
rect 4903 401 4919 435
rect 4971 401 4987 435
rect 5021 401 5037 435
rect 5089 401 5105 435
rect 5139 401 5155 435
rect 5207 401 5223 435
rect 5257 401 5273 435
rect 5325 401 5341 435
rect 5375 401 5391 435
rect 5443 401 5459 435
rect 5493 401 5509 435
rect 5561 401 5577 435
rect 5611 401 5627 435
rect 5679 401 5695 435
rect 5729 401 5745 435
rect 5797 401 5813 435
rect 5847 401 5863 435
rect 5915 401 5931 435
rect 5965 401 5981 435
rect 6033 401 6049 435
rect 6083 401 6099 435
rect 6151 401 6167 435
rect 6201 401 6217 435
rect 6269 401 6285 435
rect 6319 401 6335 435
rect 6387 401 6403 435
rect 6437 401 6453 435
rect 6505 401 6521 435
rect 6555 401 6571 435
rect 6623 401 6639 435
rect 6673 401 6689 435
rect 6741 401 6757 435
rect 6791 401 6807 435
rect 6859 401 6875 435
rect 6909 401 6925 435
rect 6977 401 6993 435
rect 7027 401 7043 435
rect 7095 401 7111 435
rect 7145 401 7161 435
rect 7213 401 7229 435
rect 7263 401 7279 435
rect 7331 401 7347 435
rect 7381 401 7397 435
rect 7449 401 7465 435
rect 7499 401 7515 435
rect 7567 401 7583 435
rect 7617 401 7633 435
rect 7685 401 7701 435
rect 7735 401 7751 435
rect 7803 401 7819 435
rect 7853 401 7869 435
rect 7921 401 7937 435
rect 7971 401 7987 435
rect 8039 401 8055 435
rect 8089 401 8105 435
rect 8157 401 8173 435
rect 8207 401 8223 435
rect 8275 401 8291 435
rect 8325 401 8341 435
rect 8393 401 8409 435
rect 8443 401 8459 435
rect 8511 401 8527 435
rect 8561 401 8577 435
rect 8629 401 8645 435
rect 8679 401 8695 435
rect 8747 401 8763 435
rect 8797 401 8813 435
rect 8865 401 8881 435
rect 8915 401 8931 435
rect 8983 401 8999 435
rect 9033 401 9049 435
rect 9101 401 9117 435
rect 9151 401 9167 435
rect 9219 401 9235 435
rect 9269 401 9285 435
rect 9337 401 9353 435
rect 9387 401 9403 435
rect 9455 401 9471 435
rect 9505 401 9521 435
rect 9573 401 9589 435
rect 9623 401 9639 435
rect 9691 401 9707 435
rect 9741 401 9757 435
rect 9809 401 9825 435
rect 9859 401 9875 435
rect 9927 401 9943 435
rect 9977 401 9993 435
rect 10045 401 10061 435
rect 10095 401 10111 435
rect 10163 401 10179 435
rect 10213 401 10229 435
rect 10281 401 10297 435
rect 10331 401 10347 435
rect 10399 401 10415 435
rect 10449 401 10465 435
rect 10517 401 10533 435
rect 10567 401 10583 435
rect 10635 401 10651 435
rect 10685 401 10701 435
rect 4810 342 4844 358
rect 4810 -250 4844 -234
rect 4928 342 4962 358
rect 4928 -250 4962 -234
rect 5046 342 5080 358
rect 5046 -250 5080 -234
rect 5164 342 5198 358
rect 5164 -250 5198 -234
rect 5282 342 5316 358
rect 5282 -250 5316 -234
rect 5400 342 5434 358
rect 5400 -250 5434 -234
rect 5518 342 5552 358
rect 5518 -250 5552 -234
rect 5636 342 5670 358
rect 5636 -250 5670 -234
rect 5754 342 5788 358
rect 5754 -250 5788 -234
rect 5872 342 5906 358
rect 5872 -250 5906 -234
rect 5990 342 6024 358
rect 5990 -250 6024 -234
rect 6108 342 6142 358
rect 6108 -250 6142 -234
rect 6226 342 6260 358
rect 6226 -250 6260 -234
rect 6344 342 6378 358
rect 6344 -250 6378 -234
rect 6462 342 6496 358
rect 6462 -250 6496 -234
rect 6580 342 6614 358
rect 6580 -250 6614 -234
rect 6698 342 6732 358
rect 6698 -250 6732 -234
rect 6816 342 6850 358
rect 6816 -250 6850 -234
rect 6934 342 6968 358
rect 6934 -250 6968 -234
rect 7052 342 7086 358
rect 7052 -250 7086 -234
rect 7170 342 7204 358
rect 7170 -250 7204 -234
rect 7288 342 7322 358
rect 7288 -250 7322 -234
rect 7406 342 7440 358
rect 7406 -250 7440 -234
rect 7524 342 7558 358
rect 7524 -250 7558 -234
rect 7642 342 7676 358
rect 7642 -250 7676 -234
rect 7760 342 7794 358
rect 7760 -250 7794 -234
rect 7878 342 7912 358
rect 7878 -250 7912 -234
rect 7996 342 8030 358
rect 7996 -250 8030 -234
rect 8114 342 8148 358
rect 8114 -250 8148 -234
rect 8232 342 8266 358
rect 8232 -250 8266 -234
rect 8350 342 8384 358
rect 8350 -250 8384 -234
rect 8468 342 8502 358
rect 8468 -250 8502 -234
rect 8586 342 8620 358
rect 8586 -250 8620 -234
rect 8704 342 8738 358
rect 8704 -250 8738 -234
rect 8822 342 8856 358
rect 8822 -250 8856 -234
rect 8940 342 8974 358
rect 8940 -250 8974 -234
rect 9058 342 9092 358
rect 9058 -250 9092 -234
rect 9176 342 9210 358
rect 9176 -250 9210 -234
rect 9294 342 9328 358
rect 9294 -250 9328 -234
rect 9412 342 9446 358
rect 9412 -250 9446 -234
rect 9530 342 9564 358
rect 9530 -250 9564 -234
rect 9648 342 9682 358
rect 9648 -250 9682 -234
rect 9766 342 9800 358
rect 9766 -250 9800 -234
rect 9884 342 9918 358
rect 9884 -250 9918 -234
rect 10002 342 10036 358
rect 10002 -250 10036 -234
rect 10120 342 10154 358
rect 10120 -250 10154 -234
rect 10238 342 10272 358
rect 10238 -250 10272 -234
rect 10356 342 10390 358
rect 10356 -250 10390 -234
rect 10474 342 10508 358
rect 10474 -250 10508 -234
rect 10592 342 10626 358
rect 10592 -250 10626 -234
rect 10710 342 10744 358
rect 10710 -250 10744 -234
rect 4696 -395 4730 -333
rect 15693 1765 15731 1799
rect 15765 1765 15803 1799
rect 15837 1765 15875 1799
rect 15909 1765 15947 1799
rect 15981 1765 16019 1799
rect 16053 1765 16091 1799
rect 16125 1765 16163 1799
rect 16197 1765 16235 1799
rect 16269 1765 16307 1799
rect 16341 1765 16379 1799
rect 15693 1691 15731 1725
rect 15765 1691 15803 1725
rect 15837 1691 15875 1725
rect 15909 1691 15947 1725
rect 15981 1691 16019 1725
rect 16053 1691 16091 1725
rect 16125 1691 16163 1725
rect 16197 1691 16235 1725
rect 16269 1691 16307 1725
rect 16341 1691 16379 1725
rect 15693 1617 15731 1651
rect 15765 1617 15803 1651
rect 15837 1617 15875 1651
rect 15909 1617 15947 1651
rect 15981 1617 16019 1651
rect 16053 1617 16091 1651
rect 16125 1617 16163 1651
rect 16197 1617 16235 1651
rect 16269 1617 16307 1651
rect 16341 1617 16379 1651
rect 15693 1543 15731 1577
rect 15765 1543 15803 1577
rect 15837 1543 15875 1577
rect 15909 1543 15947 1577
rect 15981 1543 16019 1577
rect 16053 1543 16091 1577
rect 16125 1543 16163 1577
rect 16197 1543 16235 1577
rect 16269 1543 16307 1577
rect 16341 1543 16379 1577
rect 15693 1469 15731 1503
rect 15765 1469 15803 1503
rect 15837 1469 15875 1503
rect 15909 1469 15947 1503
rect 15981 1469 16019 1503
rect 16053 1469 16091 1503
rect 16125 1469 16163 1503
rect 16197 1469 16235 1503
rect 16269 1469 16307 1503
rect 16341 1469 16379 1503
rect 15693 1395 15731 1429
rect 15765 1395 15803 1429
rect 15837 1395 15875 1429
rect 15909 1395 15947 1429
rect 15981 1395 16019 1429
rect 16053 1395 16091 1429
rect 16125 1395 16163 1429
rect 16197 1395 16235 1429
rect 16269 1395 16307 1429
rect 16341 1395 16379 1429
rect 15693 1321 15731 1355
rect 15765 1321 15803 1355
rect 15837 1321 15875 1355
rect 15909 1321 15947 1355
rect 15981 1321 16019 1355
rect 16053 1321 16091 1355
rect 16125 1321 16163 1355
rect 16197 1321 16235 1355
rect 16269 1321 16307 1355
rect 16341 1321 16379 1355
rect 15693 1247 15731 1281
rect 15765 1247 15803 1281
rect 15837 1247 15875 1281
rect 15909 1247 15947 1281
rect 15981 1247 16019 1281
rect 16053 1247 16091 1281
rect 16125 1247 16163 1281
rect 16197 1247 16235 1281
rect 16269 1247 16307 1281
rect 16341 1247 16379 1281
rect 19816 1765 19854 1799
rect 19888 1765 19926 1799
rect 19960 1765 19998 1799
rect 20032 1765 20070 1799
rect 20104 1765 20142 1799
rect 20176 1765 20214 1799
rect 20248 1765 20286 1799
rect 20320 1765 20358 1799
rect 20392 1765 20430 1799
rect 20464 1765 20502 1799
rect 19816 1691 19854 1725
rect 19888 1691 19926 1725
rect 19960 1691 19998 1725
rect 20032 1691 20070 1725
rect 20104 1691 20142 1725
rect 20176 1691 20214 1725
rect 20248 1691 20286 1725
rect 20320 1691 20358 1725
rect 20392 1691 20430 1725
rect 20464 1691 20502 1725
rect 19816 1617 19854 1651
rect 19888 1617 19926 1651
rect 19960 1617 19998 1651
rect 20032 1617 20070 1651
rect 20104 1617 20142 1651
rect 20176 1617 20214 1651
rect 20248 1617 20286 1651
rect 20320 1617 20358 1651
rect 20392 1617 20430 1651
rect 20464 1617 20502 1651
rect 19816 1543 19854 1577
rect 19888 1543 19926 1577
rect 19960 1543 19998 1577
rect 20032 1543 20070 1577
rect 20104 1543 20142 1577
rect 20176 1543 20214 1577
rect 20248 1543 20286 1577
rect 20320 1543 20358 1577
rect 20392 1543 20430 1577
rect 20464 1543 20502 1577
rect 19816 1469 19854 1503
rect 19888 1469 19926 1503
rect 19960 1469 19998 1503
rect 20032 1469 20070 1503
rect 20104 1469 20142 1503
rect 20176 1469 20214 1503
rect 20248 1469 20286 1503
rect 20320 1469 20358 1503
rect 20392 1469 20430 1503
rect 20464 1469 20502 1503
rect 19816 1395 19854 1429
rect 19888 1395 19926 1429
rect 19960 1395 19998 1429
rect 20032 1395 20070 1429
rect 20104 1395 20142 1429
rect 20176 1395 20214 1429
rect 20248 1395 20286 1429
rect 20320 1395 20358 1429
rect 20392 1395 20430 1429
rect 20464 1395 20502 1429
rect 19816 1321 19854 1355
rect 19888 1321 19926 1355
rect 19960 1321 19998 1355
rect 20032 1321 20070 1355
rect 20104 1321 20142 1355
rect 20176 1321 20214 1355
rect 20248 1321 20286 1355
rect 20320 1321 20358 1355
rect 20392 1321 20430 1355
rect 20464 1321 20502 1355
rect 19816 1247 19854 1281
rect 19888 1247 19926 1281
rect 19960 1247 19998 1281
rect 20032 1247 20070 1281
rect 20104 1247 20142 1281
rect 20176 1247 20214 1281
rect 20248 1247 20286 1281
rect 20320 1247 20358 1281
rect 20392 1247 20430 1281
rect 20464 1247 20502 1281
rect 23939 1765 23977 1799
rect 24011 1765 24049 1799
rect 24083 1765 24121 1799
rect 24155 1765 24193 1799
rect 24227 1765 24265 1799
rect 24299 1765 24337 1799
rect 24371 1765 24409 1799
rect 24443 1765 24481 1799
rect 24515 1765 24553 1799
rect 24587 1765 24625 1799
rect 23939 1691 23977 1725
rect 24011 1691 24049 1725
rect 24083 1691 24121 1725
rect 24155 1691 24193 1725
rect 24227 1691 24265 1725
rect 24299 1691 24337 1725
rect 24371 1691 24409 1725
rect 24443 1691 24481 1725
rect 24515 1691 24553 1725
rect 24587 1691 24625 1725
rect 23939 1617 23977 1651
rect 24011 1617 24049 1651
rect 24083 1617 24121 1651
rect 24155 1617 24193 1651
rect 24227 1617 24265 1651
rect 24299 1617 24337 1651
rect 24371 1617 24409 1651
rect 24443 1617 24481 1651
rect 24515 1617 24553 1651
rect 24587 1617 24625 1651
rect 23939 1543 23977 1577
rect 24011 1543 24049 1577
rect 24083 1543 24121 1577
rect 24155 1543 24193 1577
rect 24227 1543 24265 1577
rect 24299 1543 24337 1577
rect 24371 1543 24409 1577
rect 24443 1543 24481 1577
rect 24515 1543 24553 1577
rect 24587 1543 24625 1577
rect 23939 1469 23977 1503
rect 24011 1469 24049 1503
rect 24083 1469 24121 1503
rect 24155 1469 24193 1503
rect 24227 1469 24265 1503
rect 24299 1469 24337 1503
rect 24371 1469 24409 1503
rect 24443 1469 24481 1503
rect 24515 1469 24553 1503
rect 24587 1469 24625 1503
rect 23939 1395 23977 1429
rect 24011 1395 24049 1429
rect 24083 1395 24121 1429
rect 24155 1395 24193 1429
rect 24227 1395 24265 1429
rect 24299 1395 24337 1429
rect 24371 1395 24409 1429
rect 24443 1395 24481 1429
rect 24515 1395 24553 1429
rect 24587 1395 24625 1429
rect 23939 1321 23977 1355
rect 24011 1321 24049 1355
rect 24083 1321 24121 1355
rect 24155 1321 24193 1355
rect 24227 1321 24265 1355
rect 24299 1321 24337 1355
rect 24371 1321 24409 1355
rect 24443 1321 24481 1355
rect 24515 1321 24553 1355
rect 24587 1321 24625 1355
rect 23939 1247 23977 1281
rect 24011 1247 24049 1281
rect 24083 1247 24121 1281
rect 24155 1247 24193 1281
rect 24227 1247 24265 1281
rect 24299 1247 24337 1281
rect 24371 1247 24409 1281
rect 24443 1247 24481 1281
rect 24515 1247 24553 1281
rect 24587 1247 24625 1281
rect 10824 -395 10858 -333
rect 4696 -429 4776 -395
rect 10786 -429 10858 -395
rect 4709 -513 4776 -483
rect 4715 -517 4776 -513
rect 10786 -517 10794 -483
rect 4706 -605 4776 -571
rect 10786 -605 10794 -571
rect 4696 -711 4792 -677
rect 10762 -711 10858 -677
rect 4696 -773 4730 -711
rect 10824 -773 10858 -711
rect 4810 -872 4844 -856
rect 4810 -1464 4844 -1448
rect 4928 -872 4962 -856
rect 4928 -1464 4962 -1448
rect 5046 -872 5080 -856
rect 5046 -1464 5080 -1448
rect 5164 -872 5198 -856
rect 5164 -1464 5198 -1448
rect 5282 -872 5316 -856
rect 5282 -1464 5316 -1448
rect 5400 -872 5434 -856
rect 5400 -1464 5434 -1448
rect 5518 -872 5552 -856
rect 5518 -1464 5552 -1448
rect 5636 -872 5670 -856
rect 5636 -1464 5670 -1448
rect 5754 -872 5788 -856
rect 5754 -1464 5788 -1448
rect 5872 -872 5906 -856
rect 5872 -1464 5906 -1448
rect 5990 -872 6024 -856
rect 5990 -1464 6024 -1448
rect 6108 -872 6142 -856
rect 6108 -1464 6142 -1448
rect 6226 -872 6260 -856
rect 6226 -1464 6260 -1448
rect 6344 -872 6378 -856
rect 6344 -1464 6378 -1448
rect 6462 -872 6496 -856
rect 6462 -1464 6496 -1448
rect 6580 -872 6614 -856
rect 6580 -1464 6614 -1448
rect 6698 -872 6732 -856
rect 6698 -1464 6732 -1448
rect 6816 -872 6850 -856
rect 6816 -1464 6850 -1448
rect 6934 -872 6968 -856
rect 6934 -1464 6968 -1448
rect 7052 -872 7086 -856
rect 7052 -1464 7086 -1448
rect 7170 -872 7204 -856
rect 7170 -1464 7204 -1448
rect 7288 -872 7322 -856
rect 7288 -1464 7322 -1448
rect 7406 -872 7440 -856
rect 7406 -1464 7440 -1448
rect 7524 -872 7558 -856
rect 7524 -1464 7558 -1448
rect 7642 -872 7676 -856
rect 7642 -1464 7676 -1448
rect 7760 -872 7794 -856
rect 7760 -1464 7794 -1448
rect 7878 -872 7912 -856
rect 7878 -1464 7912 -1448
rect 7996 -872 8030 -856
rect 7996 -1464 8030 -1448
rect 8114 -872 8148 -856
rect 8114 -1464 8148 -1448
rect 8232 -872 8266 -856
rect 8232 -1464 8266 -1448
rect 8350 -872 8384 -856
rect 8350 -1464 8384 -1448
rect 8468 -872 8502 -856
rect 8468 -1464 8502 -1448
rect 8586 -872 8620 -856
rect 8586 -1464 8620 -1448
rect 8704 -872 8738 -856
rect 8704 -1464 8738 -1448
rect 8822 -872 8856 -856
rect 8822 -1464 8856 -1448
rect 8940 -872 8974 -856
rect 8940 -1464 8974 -1448
rect 9058 -872 9092 -856
rect 9058 -1464 9092 -1448
rect 9176 -872 9210 -856
rect 9176 -1464 9210 -1448
rect 9294 -872 9328 -856
rect 9294 -1464 9328 -1448
rect 9412 -872 9446 -856
rect 9412 -1464 9446 -1448
rect 9530 -872 9564 -856
rect 9530 -1464 9564 -1448
rect 9648 -872 9682 -856
rect 9648 -1464 9682 -1448
rect 9766 -872 9800 -856
rect 9766 -1464 9800 -1448
rect 9884 -872 9918 -856
rect 9884 -1464 9918 -1448
rect 10002 -872 10036 -856
rect 10002 -1464 10036 -1448
rect 10120 -872 10154 -856
rect 10120 -1464 10154 -1448
rect 10238 -872 10272 -856
rect 10238 -1464 10272 -1448
rect 10356 -872 10390 -856
rect 10356 -1464 10390 -1448
rect 10474 -872 10508 -856
rect 10474 -1464 10508 -1448
rect 10592 -872 10626 -856
rect 10592 -1464 10626 -1448
rect 10710 -872 10744 -856
rect 10710 -1464 10744 -1448
rect 4853 -1541 4869 -1507
rect 4903 -1541 4919 -1507
rect 4971 -1541 4987 -1507
rect 5021 -1541 5037 -1507
rect 5089 -1541 5105 -1507
rect 5139 -1541 5155 -1507
rect 5207 -1541 5223 -1507
rect 5257 -1541 5273 -1507
rect 5325 -1541 5341 -1507
rect 5375 -1541 5391 -1507
rect 5443 -1541 5459 -1507
rect 5493 -1541 5509 -1507
rect 5561 -1541 5577 -1507
rect 5611 -1541 5627 -1507
rect 5679 -1541 5695 -1507
rect 5729 -1541 5745 -1507
rect 5797 -1541 5813 -1507
rect 5847 -1541 5863 -1507
rect 5915 -1541 5931 -1507
rect 5965 -1541 5981 -1507
rect 6033 -1541 6049 -1507
rect 6083 -1541 6099 -1507
rect 6151 -1541 6167 -1507
rect 6201 -1541 6217 -1507
rect 6269 -1541 6285 -1507
rect 6319 -1541 6335 -1507
rect 6387 -1541 6403 -1507
rect 6437 -1541 6453 -1507
rect 6505 -1541 6521 -1507
rect 6555 -1541 6571 -1507
rect 6623 -1541 6639 -1507
rect 6673 -1541 6689 -1507
rect 6741 -1541 6757 -1507
rect 6791 -1541 6807 -1507
rect 6859 -1541 6875 -1507
rect 6909 -1541 6925 -1507
rect 6977 -1541 6993 -1507
rect 7027 -1541 7043 -1507
rect 7095 -1541 7111 -1507
rect 7145 -1541 7161 -1507
rect 7213 -1541 7229 -1507
rect 7263 -1541 7279 -1507
rect 7331 -1541 7347 -1507
rect 7381 -1541 7397 -1507
rect 7449 -1541 7465 -1507
rect 7499 -1541 7515 -1507
rect 7567 -1541 7583 -1507
rect 7617 -1541 7633 -1507
rect 7685 -1541 7701 -1507
rect 7735 -1541 7751 -1507
rect 7803 -1541 7819 -1507
rect 7853 -1541 7869 -1507
rect 7921 -1541 7937 -1507
rect 7971 -1541 7987 -1507
rect 8039 -1541 8055 -1507
rect 8089 -1541 8105 -1507
rect 8157 -1541 8173 -1507
rect 8207 -1541 8223 -1507
rect 8275 -1541 8291 -1507
rect 8325 -1541 8341 -1507
rect 8393 -1541 8409 -1507
rect 8443 -1541 8459 -1507
rect 8511 -1541 8527 -1507
rect 8561 -1541 8577 -1507
rect 8629 -1541 8645 -1507
rect 8679 -1541 8695 -1507
rect 8747 -1541 8763 -1507
rect 8797 -1541 8813 -1507
rect 8865 -1541 8881 -1507
rect 8915 -1541 8931 -1507
rect 8983 -1541 8999 -1507
rect 9033 -1541 9049 -1507
rect 9101 -1541 9117 -1507
rect 9151 -1541 9167 -1507
rect 9219 -1541 9235 -1507
rect 9269 -1541 9285 -1507
rect 9337 -1541 9353 -1507
rect 9387 -1541 9403 -1507
rect 9455 -1541 9471 -1507
rect 9505 -1541 9521 -1507
rect 9573 -1541 9589 -1507
rect 9623 -1541 9639 -1507
rect 9691 -1541 9707 -1507
rect 9741 -1541 9757 -1507
rect 9809 -1541 9825 -1507
rect 9859 -1541 9875 -1507
rect 9927 -1541 9943 -1507
rect 9977 -1541 9993 -1507
rect 10045 -1541 10061 -1507
rect 10095 -1541 10111 -1507
rect 10163 -1541 10179 -1507
rect 10213 -1541 10229 -1507
rect 10281 -1541 10297 -1507
rect 10331 -1541 10347 -1507
rect 10399 -1541 10415 -1507
rect 10449 -1541 10465 -1507
rect 10517 -1541 10533 -1507
rect 10567 -1541 10583 -1507
rect 10635 -1541 10651 -1507
rect 10685 -1541 10701 -1507
rect 4853 -1649 4869 -1615
rect 4903 -1649 4919 -1615
rect 4971 -1649 4987 -1615
rect 5021 -1649 5037 -1615
rect 5089 -1649 5105 -1615
rect 5139 -1649 5155 -1615
rect 5207 -1649 5223 -1615
rect 5257 -1649 5273 -1615
rect 5325 -1649 5341 -1615
rect 5375 -1649 5391 -1615
rect 5443 -1649 5459 -1615
rect 5493 -1649 5509 -1615
rect 5561 -1649 5577 -1615
rect 5611 -1649 5627 -1615
rect 5679 -1649 5695 -1615
rect 5729 -1649 5745 -1615
rect 5797 -1649 5813 -1615
rect 5847 -1649 5863 -1615
rect 5915 -1649 5931 -1615
rect 5965 -1649 5981 -1615
rect 6033 -1649 6049 -1615
rect 6083 -1649 6099 -1615
rect 6151 -1649 6167 -1615
rect 6201 -1649 6217 -1615
rect 6269 -1649 6285 -1615
rect 6319 -1649 6335 -1615
rect 6387 -1649 6403 -1615
rect 6437 -1649 6453 -1615
rect 6505 -1649 6521 -1615
rect 6555 -1649 6571 -1615
rect 6623 -1649 6639 -1615
rect 6673 -1649 6689 -1615
rect 6741 -1649 6757 -1615
rect 6791 -1649 6807 -1615
rect 6859 -1649 6875 -1615
rect 6909 -1649 6925 -1615
rect 6977 -1649 6993 -1615
rect 7027 -1649 7043 -1615
rect 7095 -1649 7111 -1615
rect 7145 -1649 7161 -1615
rect 7213 -1649 7229 -1615
rect 7263 -1649 7279 -1615
rect 7331 -1649 7347 -1615
rect 7381 -1649 7397 -1615
rect 7449 -1649 7465 -1615
rect 7499 -1649 7515 -1615
rect 7567 -1649 7583 -1615
rect 7617 -1649 7633 -1615
rect 7685 -1649 7701 -1615
rect 7735 -1649 7751 -1615
rect 7803 -1649 7819 -1615
rect 7853 -1649 7869 -1615
rect 7921 -1649 7937 -1615
rect 7971 -1649 7987 -1615
rect 8039 -1649 8055 -1615
rect 8089 -1649 8105 -1615
rect 8157 -1649 8173 -1615
rect 8207 -1649 8223 -1615
rect 8275 -1649 8291 -1615
rect 8325 -1649 8341 -1615
rect 8393 -1649 8409 -1615
rect 8443 -1649 8459 -1615
rect 8511 -1649 8527 -1615
rect 8561 -1649 8577 -1615
rect 8629 -1649 8645 -1615
rect 8679 -1649 8695 -1615
rect 8747 -1649 8763 -1615
rect 8797 -1649 8813 -1615
rect 8865 -1649 8881 -1615
rect 8915 -1649 8931 -1615
rect 8983 -1649 8999 -1615
rect 9033 -1649 9049 -1615
rect 9101 -1649 9117 -1615
rect 9151 -1649 9167 -1615
rect 9219 -1649 9235 -1615
rect 9269 -1649 9285 -1615
rect 9337 -1649 9353 -1615
rect 9387 -1649 9403 -1615
rect 9455 -1649 9471 -1615
rect 9505 -1649 9521 -1615
rect 9573 -1649 9589 -1615
rect 9623 -1649 9639 -1615
rect 9691 -1649 9707 -1615
rect 9741 -1649 9757 -1615
rect 9809 -1649 9825 -1615
rect 9859 -1649 9875 -1615
rect 9927 -1649 9943 -1615
rect 9977 -1649 9993 -1615
rect 10045 -1649 10061 -1615
rect 10095 -1649 10111 -1615
rect 10163 -1649 10179 -1615
rect 10213 -1649 10229 -1615
rect 10281 -1649 10297 -1615
rect 10331 -1649 10347 -1615
rect 10399 -1649 10415 -1615
rect 10449 -1649 10465 -1615
rect 10517 -1649 10533 -1615
rect 10567 -1649 10583 -1615
rect 10635 -1649 10651 -1615
rect 10685 -1649 10701 -1615
rect 4810 -1708 4844 -1692
rect 4810 -2300 4844 -2284
rect 4928 -1708 4962 -1692
rect 4928 -2300 4962 -2284
rect 5046 -1708 5080 -1692
rect 5046 -2300 5080 -2284
rect 5164 -1708 5198 -1692
rect 5164 -2300 5198 -2284
rect 5282 -1708 5316 -1692
rect 5282 -2300 5316 -2284
rect 5400 -1708 5434 -1692
rect 5400 -2300 5434 -2284
rect 5518 -1708 5552 -1692
rect 5518 -2300 5552 -2284
rect 5636 -1708 5670 -1692
rect 5636 -2300 5670 -2284
rect 5754 -1708 5788 -1692
rect 5754 -2300 5788 -2284
rect 5872 -1708 5906 -1692
rect 5872 -2300 5906 -2284
rect 5990 -1708 6024 -1692
rect 5990 -2300 6024 -2284
rect 6108 -1708 6142 -1692
rect 6108 -2300 6142 -2284
rect 6226 -1708 6260 -1692
rect 6226 -2300 6260 -2284
rect 6344 -1708 6378 -1692
rect 6344 -2300 6378 -2284
rect 6462 -1708 6496 -1692
rect 6462 -2300 6496 -2284
rect 6580 -1708 6614 -1692
rect 6580 -2300 6614 -2284
rect 6698 -1708 6732 -1692
rect 6698 -2300 6732 -2284
rect 6816 -1708 6850 -1692
rect 6816 -2300 6850 -2284
rect 6934 -1708 6968 -1692
rect 6934 -2300 6968 -2284
rect 7052 -1708 7086 -1692
rect 7052 -2300 7086 -2284
rect 7170 -1708 7204 -1692
rect 7170 -2300 7204 -2284
rect 7288 -1708 7322 -1692
rect 7288 -2300 7322 -2284
rect 7406 -1708 7440 -1692
rect 7406 -2300 7440 -2284
rect 7524 -1708 7558 -1692
rect 7524 -2300 7558 -2284
rect 7642 -1708 7676 -1692
rect 7642 -2300 7676 -2284
rect 7760 -1708 7794 -1692
rect 7760 -2300 7794 -2284
rect 7878 -1708 7912 -1692
rect 7878 -2300 7912 -2284
rect 7996 -1708 8030 -1692
rect 7996 -2300 8030 -2284
rect 8114 -1708 8148 -1692
rect 8114 -2300 8148 -2284
rect 8232 -1708 8266 -1692
rect 8232 -2300 8266 -2284
rect 8350 -1708 8384 -1692
rect 8350 -2300 8384 -2284
rect 8468 -1708 8502 -1692
rect 8468 -2300 8502 -2284
rect 8586 -1708 8620 -1692
rect 8586 -2300 8620 -2284
rect 8704 -1708 8738 -1692
rect 8704 -2300 8738 -2284
rect 8822 -1708 8856 -1692
rect 8822 -2300 8856 -2284
rect 8940 -1708 8974 -1692
rect 8940 -2300 8974 -2284
rect 9058 -1708 9092 -1692
rect 9058 -2300 9092 -2284
rect 9176 -1708 9210 -1692
rect 9176 -2300 9210 -2284
rect 9294 -1708 9328 -1692
rect 9294 -2300 9328 -2284
rect 9412 -1708 9446 -1692
rect 9412 -2300 9446 -2284
rect 9530 -1708 9564 -1692
rect 9530 -2300 9564 -2284
rect 9648 -1708 9682 -1692
rect 9648 -2300 9682 -2284
rect 9766 -1708 9800 -1692
rect 9766 -2300 9800 -2284
rect 9884 -1708 9918 -1692
rect 9884 -2300 9918 -2284
rect 10002 -1708 10036 -1692
rect 10002 -2300 10036 -2284
rect 10120 -1708 10154 -1692
rect 10120 -2300 10154 -2284
rect 10238 -1708 10272 -1692
rect 10238 -2300 10272 -2284
rect 10356 -1708 10390 -1692
rect 10356 -2300 10390 -2284
rect 10474 -1708 10508 -1692
rect 10474 -2300 10508 -2284
rect 10592 -1708 10626 -1692
rect 10592 -2300 10626 -2284
rect 10710 -1708 10744 -1692
rect 10710 -2300 10744 -2284
rect 4696 -2445 4730 -2383
rect 10824 -2445 10858 -2383
rect 4696 -2479 4776 -2445
rect 10786 -2479 10858 -2445
rect 4703 -2564 4776 -2533
rect 4709 -2567 4776 -2564
rect 10786 -2567 10794 -2533
rect 4711 -2651 4776 -2621
rect 4714 -2655 4776 -2651
rect 10786 -2655 10794 -2621
rect 4696 -2761 4792 -2727
rect 10762 -2761 10858 -2727
rect 4696 -2823 4730 -2761
rect 10824 -2823 10858 -2761
rect 4810 -2922 4844 -2906
rect 4810 -3514 4844 -3498
rect 4928 -2922 4962 -2906
rect 4928 -3514 4962 -3498
rect 5046 -2922 5080 -2906
rect 5046 -3514 5080 -3498
rect 5164 -2922 5198 -2906
rect 5164 -3514 5198 -3498
rect 5282 -2922 5316 -2906
rect 5282 -3514 5316 -3498
rect 5400 -2922 5434 -2906
rect 5400 -3514 5434 -3498
rect 5518 -2922 5552 -2906
rect 5518 -3514 5552 -3498
rect 5636 -2922 5670 -2906
rect 5636 -3514 5670 -3498
rect 5754 -2922 5788 -2906
rect 5754 -3514 5788 -3498
rect 5872 -2922 5906 -2906
rect 5872 -3514 5906 -3498
rect 5990 -2922 6024 -2906
rect 5990 -3514 6024 -3498
rect 6108 -2922 6142 -2906
rect 6108 -3514 6142 -3498
rect 6226 -2922 6260 -2906
rect 6226 -3514 6260 -3498
rect 6344 -2922 6378 -2906
rect 6344 -3514 6378 -3498
rect 6462 -2922 6496 -2906
rect 6462 -3514 6496 -3498
rect 6580 -2922 6614 -2906
rect 6580 -3514 6614 -3498
rect 6698 -2922 6732 -2906
rect 6698 -3514 6732 -3498
rect 6816 -2922 6850 -2906
rect 6816 -3514 6850 -3498
rect 6934 -2922 6968 -2906
rect 6934 -3514 6968 -3498
rect 7052 -2922 7086 -2906
rect 7052 -3514 7086 -3498
rect 7170 -2922 7204 -2906
rect 7170 -3514 7204 -3498
rect 7288 -2922 7322 -2906
rect 7288 -3514 7322 -3498
rect 7406 -2922 7440 -2906
rect 7406 -3514 7440 -3498
rect 7524 -2922 7558 -2906
rect 7524 -3514 7558 -3498
rect 7642 -2922 7676 -2906
rect 7642 -3514 7676 -3498
rect 7760 -2922 7794 -2906
rect 7760 -3514 7794 -3498
rect 7878 -2922 7912 -2906
rect 7878 -3514 7912 -3498
rect 7996 -2922 8030 -2906
rect 7996 -3514 8030 -3498
rect 8114 -2922 8148 -2906
rect 8114 -3514 8148 -3498
rect 8232 -2922 8266 -2906
rect 8232 -3514 8266 -3498
rect 8350 -2922 8384 -2906
rect 8350 -3514 8384 -3498
rect 8468 -2922 8502 -2906
rect 8468 -3514 8502 -3498
rect 8586 -2922 8620 -2906
rect 8586 -3514 8620 -3498
rect 8704 -2922 8738 -2906
rect 8704 -3514 8738 -3498
rect 8822 -2922 8856 -2906
rect 8822 -3514 8856 -3498
rect 8940 -2922 8974 -2906
rect 8940 -3514 8974 -3498
rect 9058 -2922 9092 -2906
rect 9058 -3514 9092 -3498
rect 9176 -2922 9210 -2906
rect 9176 -3514 9210 -3498
rect 9294 -2922 9328 -2906
rect 9294 -3514 9328 -3498
rect 9412 -2922 9446 -2906
rect 9412 -3514 9446 -3498
rect 9530 -2922 9564 -2906
rect 9530 -3514 9564 -3498
rect 9648 -2922 9682 -2906
rect 9648 -3514 9682 -3498
rect 9766 -2922 9800 -2906
rect 9766 -3514 9800 -3498
rect 9884 -2922 9918 -2906
rect 9884 -3514 9918 -3498
rect 10002 -2922 10036 -2906
rect 10002 -3514 10036 -3498
rect 10120 -2922 10154 -2906
rect 10120 -3514 10154 -3498
rect 10238 -2922 10272 -2906
rect 10238 -3514 10272 -3498
rect 10356 -2922 10390 -2906
rect 10356 -3514 10390 -3498
rect 10474 -2922 10508 -2906
rect 10474 -3514 10508 -3498
rect 10592 -2922 10626 -2906
rect 10592 -3514 10626 -3498
rect 10710 -2922 10744 -2906
rect 10710 -3514 10744 -3498
rect 4853 -3591 4869 -3557
rect 4903 -3591 4919 -3557
rect 4971 -3591 4987 -3557
rect 5021 -3591 5037 -3557
rect 5089 -3591 5105 -3557
rect 5139 -3591 5155 -3557
rect 5207 -3591 5223 -3557
rect 5257 -3591 5273 -3557
rect 5325 -3591 5341 -3557
rect 5375 -3591 5391 -3557
rect 5443 -3591 5459 -3557
rect 5493 -3591 5509 -3557
rect 5561 -3591 5577 -3557
rect 5611 -3591 5627 -3557
rect 5679 -3591 5695 -3557
rect 5729 -3591 5745 -3557
rect 5797 -3591 5813 -3557
rect 5847 -3591 5863 -3557
rect 5915 -3591 5931 -3557
rect 5965 -3591 5981 -3557
rect 6033 -3591 6049 -3557
rect 6083 -3591 6099 -3557
rect 6151 -3591 6167 -3557
rect 6201 -3591 6217 -3557
rect 6269 -3591 6285 -3557
rect 6319 -3591 6335 -3557
rect 6387 -3591 6403 -3557
rect 6437 -3591 6453 -3557
rect 6505 -3591 6521 -3557
rect 6555 -3591 6571 -3557
rect 6623 -3591 6639 -3557
rect 6673 -3591 6689 -3557
rect 6741 -3591 6757 -3557
rect 6791 -3591 6807 -3557
rect 6859 -3591 6875 -3557
rect 6909 -3591 6925 -3557
rect 6977 -3591 6993 -3557
rect 7027 -3591 7043 -3557
rect 7095 -3591 7111 -3557
rect 7145 -3591 7161 -3557
rect 7213 -3591 7229 -3557
rect 7263 -3591 7279 -3557
rect 7331 -3591 7347 -3557
rect 7381 -3591 7397 -3557
rect 7449 -3591 7465 -3557
rect 7499 -3591 7515 -3557
rect 7567 -3591 7583 -3557
rect 7617 -3591 7633 -3557
rect 7685 -3591 7701 -3557
rect 7735 -3591 7751 -3557
rect 7803 -3591 7819 -3557
rect 7853 -3591 7869 -3557
rect 7921 -3591 7937 -3557
rect 7971 -3591 7987 -3557
rect 8039 -3591 8055 -3557
rect 8089 -3591 8105 -3557
rect 8157 -3591 8173 -3557
rect 8207 -3591 8223 -3557
rect 8275 -3591 8291 -3557
rect 8325 -3591 8341 -3557
rect 8393 -3591 8409 -3557
rect 8443 -3591 8459 -3557
rect 8511 -3591 8527 -3557
rect 8561 -3591 8577 -3557
rect 8629 -3591 8645 -3557
rect 8679 -3591 8695 -3557
rect 8747 -3591 8763 -3557
rect 8797 -3591 8813 -3557
rect 8865 -3591 8881 -3557
rect 8915 -3591 8931 -3557
rect 8983 -3591 8999 -3557
rect 9033 -3591 9049 -3557
rect 9101 -3591 9117 -3557
rect 9151 -3591 9167 -3557
rect 9219 -3591 9235 -3557
rect 9269 -3591 9285 -3557
rect 9337 -3591 9353 -3557
rect 9387 -3591 9403 -3557
rect 9455 -3591 9471 -3557
rect 9505 -3591 9521 -3557
rect 9573 -3591 9589 -3557
rect 9623 -3591 9639 -3557
rect 9691 -3591 9707 -3557
rect 9741 -3591 9757 -3557
rect 9809 -3591 9825 -3557
rect 9859 -3591 9875 -3557
rect 9927 -3591 9943 -3557
rect 9977 -3591 9993 -3557
rect 10045 -3591 10061 -3557
rect 10095 -3591 10111 -3557
rect 10163 -3591 10179 -3557
rect 10213 -3591 10229 -3557
rect 10281 -3591 10297 -3557
rect 10331 -3591 10347 -3557
rect 10399 -3591 10415 -3557
rect 10449 -3591 10465 -3557
rect 10517 -3591 10533 -3557
rect 10567 -3591 10583 -3557
rect 10635 -3591 10651 -3557
rect 10685 -3591 10701 -3557
rect 4853 -3699 4869 -3665
rect 4903 -3699 4919 -3665
rect 4971 -3699 4987 -3665
rect 5021 -3699 5037 -3665
rect 5089 -3699 5105 -3665
rect 5139 -3699 5155 -3665
rect 5207 -3699 5223 -3665
rect 5257 -3699 5273 -3665
rect 5325 -3699 5341 -3665
rect 5375 -3699 5391 -3665
rect 5443 -3699 5459 -3665
rect 5493 -3699 5509 -3665
rect 5561 -3699 5577 -3665
rect 5611 -3699 5627 -3665
rect 5679 -3699 5695 -3665
rect 5729 -3699 5745 -3665
rect 5797 -3699 5813 -3665
rect 5847 -3699 5863 -3665
rect 5915 -3699 5931 -3665
rect 5965 -3699 5981 -3665
rect 6033 -3699 6049 -3665
rect 6083 -3699 6099 -3665
rect 6151 -3699 6167 -3665
rect 6201 -3699 6217 -3665
rect 6269 -3699 6285 -3665
rect 6319 -3699 6335 -3665
rect 6387 -3699 6403 -3665
rect 6437 -3699 6453 -3665
rect 6505 -3699 6521 -3665
rect 6555 -3699 6571 -3665
rect 6623 -3699 6639 -3665
rect 6673 -3699 6689 -3665
rect 6741 -3699 6757 -3665
rect 6791 -3699 6807 -3665
rect 6859 -3699 6875 -3665
rect 6909 -3699 6925 -3665
rect 6977 -3699 6993 -3665
rect 7027 -3699 7043 -3665
rect 7095 -3699 7111 -3665
rect 7145 -3699 7161 -3665
rect 7213 -3699 7229 -3665
rect 7263 -3699 7279 -3665
rect 7331 -3699 7347 -3665
rect 7381 -3699 7397 -3665
rect 7449 -3699 7465 -3665
rect 7499 -3699 7515 -3665
rect 7567 -3699 7583 -3665
rect 7617 -3699 7633 -3665
rect 7685 -3699 7701 -3665
rect 7735 -3699 7751 -3665
rect 7803 -3699 7819 -3665
rect 7853 -3699 7869 -3665
rect 7921 -3699 7937 -3665
rect 7971 -3699 7987 -3665
rect 8039 -3699 8055 -3665
rect 8089 -3699 8105 -3665
rect 8157 -3699 8173 -3665
rect 8207 -3699 8223 -3665
rect 8275 -3699 8291 -3665
rect 8325 -3699 8341 -3665
rect 8393 -3699 8409 -3665
rect 8443 -3699 8459 -3665
rect 8511 -3699 8527 -3665
rect 8561 -3699 8577 -3665
rect 8629 -3699 8645 -3665
rect 8679 -3699 8695 -3665
rect 8747 -3699 8763 -3665
rect 8797 -3699 8813 -3665
rect 8865 -3699 8881 -3665
rect 8915 -3699 8931 -3665
rect 8983 -3699 8999 -3665
rect 9033 -3699 9049 -3665
rect 9101 -3699 9117 -3665
rect 9151 -3699 9167 -3665
rect 9219 -3699 9235 -3665
rect 9269 -3699 9285 -3665
rect 9337 -3699 9353 -3665
rect 9387 -3699 9403 -3665
rect 9455 -3699 9471 -3665
rect 9505 -3699 9521 -3665
rect 9573 -3699 9589 -3665
rect 9623 -3699 9639 -3665
rect 9691 -3699 9707 -3665
rect 9741 -3699 9757 -3665
rect 9809 -3699 9825 -3665
rect 9859 -3699 9875 -3665
rect 9927 -3699 9943 -3665
rect 9977 -3699 9993 -3665
rect 10045 -3699 10061 -3665
rect 10095 -3699 10111 -3665
rect 10163 -3699 10179 -3665
rect 10213 -3699 10229 -3665
rect 10281 -3699 10297 -3665
rect 10331 -3699 10347 -3665
rect 10399 -3699 10415 -3665
rect 10449 -3699 10465 -3665
rect 10517 -3699 10533 -3665
rect 10567 -3699 10583 -3665
rect 10635 -3699 10651 -3665
rect 10685 -3699 10701 -3665
rect 4810 -3758 4844 -3742
rect 4810 -4350 4844 -4334
rect 4928 -3758 4962 -3742
rect 4928 -4350 4962 -4334
rect 5046 -3758 5080 -3742
rect 5046 -4350 5080 -4334
rect 5164 -3758 5198 -3742
rect 5164 -4350 5198 -4334
rect 5282 -3758 5316 -3742
rect 5282 -4350 5316 -4334
rect 5400 -3758 5434 -3742
rect 5400 -4350 5434 -4334
rect 5518 -3758 5552 -3742
rect 5518 -4350 5552 -4334
rect 5636 -3758 5670 -3742
rect 5636 -4350 5670 -4334
rect 5754 -3758 5788 -3742
rect 5754 -4350 5788 -4334
rect 5872 -3758 5906 -3742
rect 5872 -4350 5906 -4334
rect 5990 -3758 6024 -3742
rect 5990 -4350 6024 -4334
rect 6108 -3758 6142 -3742
rect 6108 -4350 6142 -4334
rect 6226 -3758 6260 -3742
rect 6226 -4350 6260 -4334
rect 6344 -3758 6378 -3742
rect 6344 -4350 6378 -4334
rect 6462 -3758 6496 -3742
rect 6462 -4350 6496 -4334
rect 6580 -3758 6614 -3742
rect 6580 -4350 6614 -4334
rect 6698 -3758 6732 -3742
rect 6698 -4350 6732 -4334
rect 6816 -3758 6850 -3742
rect 6816 -4350 6850 -4334
rect 6934 -3758 6968 -3742
rect 6934 -4350 6968 -4334
rect 7052 -3758 7086 -3742
rect 7052 -4350 7086 -4334
rect 7170 -3758 7204 -3742
rect 7170 -4350 7204 -4334
rect 7288 -3758 7322 -3742
rect 7288 -4350 7322 -4334
rect 7406 -3758 7440 -3742
rect 7406 -4350 7440 -4334
rect 7524 -3758 7558 -3742
rect 7524 -4350 7558 -4334
rect 7642 -3758 7676 -3742
rect 7642 -4350 7676 -4334
rect 7760 -3758 7794 -3742
rect 7760 -4350 7794 -4334
rect 7878 -3758 7912 -3742
rect 7878 -4350 7912 -4334
rect 7996 -3758 8030 -3742
rect 7996 -4350 8030 -4334
rect 8114 -3758 8148 -3742
rect 8114 -4350 8148 -4334
rect 8232 -3758 8266 -3742
rect 8232 -4350 8266 -4334
rect 8350 -3758 8384 -3742
rect 8350 -4350 8384 -4334
rect 8468 -3758 8502 -3742
rect 8468 -4350 8502 -4334
rect 8586 -3758 8620 -3742
rect 8586 -4350 8620 -4334
rect 8704 -3758 8738 -3742
rect 8704 -4350 8738 -4334
rect 8822 -3758 8856 -3742
rect 8822 -4350 8856 -4334
rect 8940 -3758 8974 -3742
rect 8940 -4350 8974 -4334
rect 9058 -3758 9092 -3742
rect 9058 -4350 9092 -4334
rect 9176 -3758 9210 -3742
rect 9176 -4350 9210 -4334
rect 9294 -3758 9328 -3742
rect 9294 -4350 9328 -4334
rect 9412 -3758 9446 -3742
rect 9412 -4350 9446 -4334
rect 9530 -3758 9564 -3742
rect 9530 -4350 9564 -4334
rect 9648 -3758 9682 -3742
rect 9648 -4350 9682 -4334
rect 9766 -3758 9800 -3742
rect 9766 -4350 9800 -4334
rect 9884 -3758 9918 -3742
rect 9884 -4350 9918 -4334
rect 10002 -3758 10036 -3742
rect 10002 -4350 10036 -4334
rect 10120 -3758 10154 -3742
rect 10120 -4350 10154 -4334
rect 10238 -3758 10272 -3742
rect 10238 -4350 10272 -4334
rect 10356 -3758 10390 -3742
rect 10356 -4350 10390 -4334
rect 10474 -3758 10508 -3742
rect 10474 -4350 10508 -4334
rect 10592 -3758 10626 -3742
rect 10592 -4350 10626 -4334
rect 10710 -3758 10744 -3742
rect 10710 -4350 10744 -4334
rect 4696 -4495 4730 -4433
rect 10824 -4495 10858 -4433
rect 4696 -4529 4768 -4495
rect 10778 -4529 10858 -4495
rect 4709 -4591 4768 -4583
rect 4714 -4617 4768 -4591
rect 10778 -4617 10808 -4583
rect 4707 -4701 4768 -4671
rect 4719 -4705 4768 -4701
rect 10778 -4705 10808 -4671
rect 4853 -5641 4869 -5607
rect 4903 -5641 4919 -5607
rect 4971 -5641 4987 -5607
rect 5021 -5641 5037 -5607
rect 5089 -5641 5105 -5607
rect 5139 -5641 5155 -5607
rect 5207 -5641 5223 -5607
rect 5257 -5641 5273 -5607
rect 5325 -5641 5341 -5607
rect 5375 -5641 5391 -5607
rect 5443 -5641 5459 -5607
rect 5493 -5641 5509 -5607
rect 5561 -5641 5577 -5607
rect 5611 -5641 5627 -5607
rect 5679 -5641 5695 -5607
rect 5729 -5641 5745 -5607
rect 5797 -5641 5813 -5607
rect 5847 -5641 5863 -5607
rect 5915 -5641 5931 -5607
rect 5965 -5641 5981 -5607
rect 6033 -5641 6049 -5607
rect 6083 -5641 6099 -5607
rect 6151 -5641 6167 -5607
rect 6201 -5641 6217 -5607
rect 6269 -5641 6285 -5607
rect 6319 -5641 6335 -5607
rect 6387 -5641 6403 -5607
rect 6437 -5641 6453 -5607
rect 6505 -5641 6521 -5607
rect 6555 -5641 6571 -5607
rect 6623 -5641 6639 -5607
rect 6673 -5641 6689 -5607
rect 6741 -5641 6757 -5607
rect 6791 -5641 6807 -5607
rect 6859 -5641 6875 -5607
rect 6909 -5641 6925 -5607
rect 6977 -5641 6993 -5607
rect 7027 -5641 7043 -5607
rect 7095 -5641 7111 -5607
rect 7145 -5641 7161 -5607
rect 7213 -5641 7229 -5607
rect 7263 -5641 7279 -5607
rect 7331 -5641 7347 -5607
rect 7381 -5641 7397 -5607
rect 7449 -5641 7465 -5607
rect 7499 -5641 7515 -5607
rect 7567 -5641 7583 -5607
rect 7617 -5641 7633 -5607
rect 7685 -5641 7701 -5607
rect 7735 -5641 7751 -5607
rect 7803 -5641 7819 -5607
rect 7853 -5641 7869 -5607
rect 7921 -5641 7937 -5607
rect 7971 -5641 7987 -5607
rect 8039 -5641 8055 -5607
rect 8089 -5641 8105 -5607
rect 8157 -5641 8173 -5607
rect 8207 -5641 8223 -5607
rect 8275 -5641 8291 -5607
rect 8325 -5641 8341 -5607
rect 8393 -5641 8409 -5607
rect 8443 -5641 8459 -5607
rect 8511 -5641 8527 -5607
rect 8561 -5641 8577 -5607
rect 8629 -5641 8645 -5607
rect 8679 -5641 8695 -5607
rect 8747 -5641 8763 -5607
rect 8797 -5641 8813 -5607
rect 8865 -5641 8881 -5607
rect 8915 -5641 8931 -5607
rect 8983 -5641 8999 -5607
rect 9033 -5641 9049 -5607
rect 9101 -5641 9117 -5607
rect 9151 -5641 9167 -5607
rect 9219 -5641 9235 -5607
rect 9269 -5641 9285 -5607
rect 9337 -5641 9353 -5607
rect 9387 -5641 9403 -5607
rect 9455 -5641 9471 -5607
rect 9505 -5641 9521 -5607
rect 9573 -5641 9589 -5607
rect 9623 -5641 9639 -5607
rect 9691 -5641 9707 -5607
rect 9741 -5641 9757 -5607
rect 9809 -5641 9825 -5607
rect 9859 -5641 9875 -5607
rect 9927 -5641 9943 -5607
rect 9977 -5641 9993 -5607
rect 10045 -5641 10061 -5607
rect 10095 -5641 10111 -5607
rect 10163 -5641 10179 -5607
rect 10213 -5641 10229 -5607
rect 10281 -5641 10297 -5607
rect 10331 -5641 10347 -5607
rect 10399 -5641 10415 -5607
rect 10449 -5641 10465 -5607
rect 10517 -5641 10533 -5607
rect 10567 -5641 10583 -5607
rect 10635 -5641 10651 -5607
rect 10685 -5641 10701 -5607
rect 4853 -5749 4869 -5715
rect 4903 -5749 4919 -5715
rect 4971 -5749 4987 -5715
rect 5021 -5749 5037 -5715
rect 5089 -5749 5105 -5715
rect 5139 -5749 5155 -5715
rect 5207 -5749 5223 -5715
rect 5257 -5749 5273 -5715
rect 5325 -5749 5341 -5715
rect 5375 -5749 5391 -5715
rect 5443 -5749 5459 -5715
rect 5493 -5749 5509 -5715
rect 5561 -5749 5577 -5715
rect 5611 -5749 5627 -5715
rect 5679 -5749 5695 -5715
rect 5729 -5749 5745 -5715
rect 5797 -5749 5813 -5715
rect 5847 -5749 5863 -5715
rect 5915 -5749 5931 -5715
rect 5965 -5749 5981 -5715
rect 6033 -5749 6049 -5715
rect 6083 -5749 6099 -5715
rect 6151 -5749 6167 -5715
rect 6201 -5749 6217 -5715
rect 6269 -5749 6285 -5715
rect 6319 -5749 6335 -5715
rect 6387 -5749 6403 -5715
rect 6437 -5749 6453 -5715
rect 6505 -5749 6521 -5715
rect 6555 -5749 6571 -5715
rect 6623 -5749 6639 -5715
rect 6673 -5749 6689 -5715
rect 6741 -5749 6757 -5715
rect 6791 -5749 6807 -5715
rect 6859 -5749 6875 -5715
rect 6909 -5749 6925 -5715
rect 6977 -5749 6993 -5715
rect 7027 -5749 7043 -5715
rect 7095 -5749 7111 -5715
rect 7145 -5749 7161 -5715
rect 7213 -5749 7229 -5715
rect 7263 -5749 7279 -5715
rect 7331 -5749 7347 -5715
rect 7381 -5749 7397 -5715
rect 7449 -5749 7465 -5715
rect 7499 -5749 7515 -5715
rect 7567 -5749 7583 -5715
rect 7617 -5749 7633 -5715
rect 7685 -5749 7701 -5715
rect 7735 -5749 7751 -5715
rect 7803 -5749 7819 -5715
rect 7853 -5749 7869 -5715
rect 7921 -5749 7937 -5715
rect 7971 -5749 7987 -5715
rect 8039 -5749 8055 -5715
rect 8089 -5749 8105 -5715
rect 8157 -5749 8173 -5715
rect 8207 -5749 8223 -5715
rect 8275 -5749 8291 -5715
rect 8325 -5749 8341 -5715
rect 8393 -5749 8409 -5715
rect 8443 -5749 8459 -5715
rect 8511 -5749 8527 -5715
rect 8561 -5749 8577 -5715
rect 8629 -5749 8645 -5715
rect 8679 -5749 8695 -5715
rect 8747 -5749 8763 -5715
rect 8797 -5749 8813 -5715
rect 8865 -5749 8881 -5715
rect 8915 -5749 8931 -5715
rect 8983 -5749 8999 -5715
rect 9033 -5749 9049 -5715
rect 9101 -5749 9117 -5715
rect 9151 -5749 9167 -5715
rect 9219 -5749 9235 -5715
rect 9269 -5749 9285 -5715
rect 9337 -5749 9353 -5715
rect 9387 -5749 9403 -5715
rect 9455 -5749 9471 -5715
rect 9505 -5749 9521 -5715
rect 9573 -5749 9589 -5715
rect 9623 -5749 9639 -5715
rect 9691 -5749 9707 -5715
rect 9741 -5749 9757 -5715
rect 9809 -5749 9825 -5715
rect 9859 -5749 9875 -5715
rect 9927 -5749 9943 -5715
rect 9977 -5749 9993 -5715
rect 10045 -5749 10061 -5715
rect 10095 -5749 10111 -5715
rect 10163 -5749 10179 -5715
rect 10213 -5749 10229 -5715
rect 10281 -5749 10297 -5715
rect 10331 -5749 10347 -5715
rect 10399 -5749 10415 -5715
rect 10449 -5749 10465 -5715
rect 10517 -5749 10533 -5715
rect 10567 -5749 10583 -5715
rect 10635 -5749 10651 -5715
rect 10685 -5749 10701 -5715
rect 4776 -6667 4792 -6633
rect 10762 -6667 10778 -6633
rect 4776 -6755 4792 -6721
rect 10762 -6755 10778 -6721
rect 4132 -7159 4170 -7125
rect 4204 -7159 4242 -7125
rect 4276 -7159 4314 -7125
rect 4348 -7159 4386 -7125
rect 4420 -7159 4458 -7125
rect 4492 -7159 4530 -7125
rect 4564 -7159 4602 -7125
rect 4636 -7159 4674 -7125
rect 4708 -7159 4746 -7125
rect 4780 -7159 4818 -7125
rect 4852 -7159 4890 -7125
rect 4924 -7159 4962 -7125
rect 4996 -7159 5034 -7125
rect 5068 -7159 5106 -7125
rect 5140 -7159 5178 -7125
rect 5212 -7159 5250 -7125
rect 5284 -7159 5322 -7125
rect 5356 -7159 5394 -7125
rect 5428 -7159 5466 -7125
rect 5500 -7159 5538 -7125
rect 4132 -7233 4170 -7199
rect 4204 -7233 4242 -7199
rect 4276 -7233 4314 -7199
rect 4348 -7233 4386 -7199
rect 4420 -7233 4458 -7199
rect 4492 -7233 4530 -7199
rect 4564 -7233 4602 -7199
rect 4636 -7233 4674 -7199
rect 4708 -7233 4746 -7199
rect 4780 -7233 4818 -7199
rect 4852 -7233 4890 -7199
rect 4924 -7233 4962 -7199
rect 4996 -7233 5034 -7199
rect 5068 -7233 5106 -7199
rect 5140 -7233 5178 -7199
rect 5212 -7233 5250 -7199
rect 5284 -7233 5322 -7199
rect 5356 -7233 5394 -7199
rect 5428 -7233 5466 -7199
rect 5500 -7233 5538 -7199
rect 4132 -7307 4170 -7273
rect 4204 -7307 4242 -7273
rect 4276 -7307 4314 -7273
rect 4348 -7307 4386 -7273
rect 4420 -7307 4458 -7273
rect 4492 -7307 4530 -7273
rect 4564 -7307 4602 -7273
rect 4636 -7307 4674 -7273
rect 4708 -7307 4746 -7273
rect 4780 -7307 4818 -7273
rect 4852 -7307 4890 -7273
rect 4924 -7307 4962 -7273
rect 4996 -7307 5034 -7273
rect 5068 -7307 5106 -7273
rect 5140 -7307 5178 -7273
rect 5212 -7307 5250 -7273
rect 5284 -7307 5322 -7273
rect 5356 -7307 5394 -7273
rect 5428 -7307 5466 -7273
rect 5500 -7307 5538 -7273
rect 4132 -7381 4170 -7347
rect 4204 -7381 4242 -7347
rect 4276 -7381 4314 -7347
rect 4348 -7381 4386 -7347
rect 4420 -7381 4458 -7347
rect 4492 -7381 4530 -7347
rect 4564 -7381 4602 -7347
rect 4636 -7381 4674 -7347
rect 4708 -7381 4746 -7347
rect 4780 -7381 4818 -7347
rect 4852 -7381 4890 -7347
rect 4924 -7381 4962 -7347
rect 4996 -7381 5034 -7347
rect 5068 -7381 5106 -7347
rect 5140 -7381 5178 -7347
rect 5212 -7381 5250 -7347
rect 5284 -7381 5322 -7347
rect 5356 -7381 5394 -7347
rect 5428 -7381 5466 -7347
rect 5500 -7381 5538 -7347
rect 4132 -7455 4170 -7421
rect 4204 -7455 4242 -7421
rect 4276 -7455 4314 -7421
rect 4348 -7455 4386 -7421
rect 4420 -7455 4458 -7421
rect 4492 -7455 4530 -7421
rect 4564 -7455 4602 -7421
rect 4636 -7455 4674 -7421
rect 4708 -7455 4746 -7421
rect 4780 -7455 4818 -7421
rect 4852 -7455 4890 -7421
rect 4924 -7455 4962 -7421
rect 4996 -7455 5034 -7421
rect 5068 -7455 5106 -7421
rect 5140 -7455 5178 -7421
rect 5212 -7455 5250 -7421
rect 5284 -7455 5322 -7421
rect 5356 -7455 5394 -7421
rect 5428 -7455 5466 -7421
rect 5500 -7455 5538 -7421
rect 4132 -7529 4170 -7495
rect 4204 -7529 4242 -7495
rect 4276 -7529 4314 -7495
rect 4348 -7529 4386 -7495
rect 4420 -7529 4458 -7495
rect 4492 -7529 4530 -7495
rect 4564 -7529 4602 -7495
rect 4636 -7529 4674 -7495
rect 4708 -7529 4746 -7495
rect 4780 -7529 4818 -7495
rect 4852 -7529 4890 -7495
rect 4924 -7529 4962 -7495
rect 4996 -7529 5034 -7495
rect 5068 -7529 5106 -7495
rect 5140 -7529 5178 -7495
rect 5212 -7529 5250 -7495
rect 5284 -7529 5322 -7495
rect 5356 -7529 5394 -7495
rect 5428 -7529 5466 -7495
rect 5500 -7529 5538 -7495
rect 4132 -7603 4170 -7569
rect 4204 -7603 4242 -7569
rect 4276 -7603 4314 -7569
rect 4348 -7603 4386 -7569
rect 4420 -7603 4458 -7569
rect 4492 -7603 4530 -7569
rect 4564 -7603 4602 -7569
rect 4636 -7603 4674 -7569
rect 4708 -7603 4746 -7569
rect 4780 -7603 4818 -7569
rect 4852 -7603 4890 -7569
rect 4924 -7603 4962 -7569
rect 4996 -7603 5034 -7569
rect 5068 -7603 5106 -7569
rect 5140 -7603 5178 -7569
rect 5212 -7603 5250 -7569
rect 5284 -7603 5322 -7569
rect 5356 -7603 5394 -7569
rect 5428 -7603 5466 -7569
rect 5500 -7603 5538 -7569
rect 4132 -7677 4170 -7643
rect 4204 -7677 4242 -7643
rect 4276 -7677 4314 -7643
rect 4348 -7677 4386 -7643
rect 4420 -7677 4458 -7643
rect 4492 -7677 4530 -7643
rect 4564 -7677 4602 -7643
rect 4636 -7677 4674 -7643
rect 4708 -7677 4746 -7643
rect 4780 -7677 4818 -7643
rect 4852 -7677 4890 -7643
rect 4924 -7677 4962 -7643
rect 4996 -7677 5034 -7643
rect 5068 -7677 5106 -7643
rect 5140 -7677 5178 -7643
rect 5212 -7677 5250 -7643
rect 5284 -7677 5322 -7643
rect 5356 -7677 5394 -7643
rect 5428 -7677 5466 -7643
rect 5500 -7677 5538 -7643
rect 4132 -7751 4170 -7717
rect 4204 -7751 4242 -7717
rect 4276 -7751 4314 -7717
rect 4348 -7751 4386 -7717
rect 4420 -7751 4458 -7717
rect 4492 -7751 4530 -7717
rect 4564 -7751 4602 -7717
rect 4636 -7751 4674 -7717
rect 4708 -7751 4746 -7717
rect 4780 -7751 4818 -7717
rect 4852 -7751 4890 -7717
rect 4924 -7751 4962 -7717
rect 4996 -7751 5034 -7717
rect 5068 -7751 5106 -7717
rect 5140 -7751 5178 -7717
rect 5212 -7751 5250 -7717
rect 5284 -7751 5322 -7717
rect 5356 -7751 5394 -7717
rect 5428 -7751 5466 -7717
rect 5500 -7751 5538 -7717
rect 9868 -7223 9906 -7189
rect 9940 -7223 9978 -7189
rect 10012 -7223 10050 -7189
rect 10084 -7223 10122 -7189
rect 10156 -7223 10194 -7189
rect 10228 -7223 10266 -7189
rect 10300 -7223 10337 -7189
rect 10771 -7225 10777 -7191
rect 11087 -7225 11093 -7191
rect 11403 -7225 11409 -7191
rect 11719 -7225 11725 -7191
rect 12035 -7225 12041 -7191
rect 12351 -7225 12357 -7191
rect 9868 -7297 9906 -7263
rect 9940 -7297 9978 -7263
rect 10012 -7297 10050 -7263
rect 10084 -7297 10122 -7263
rect 10156 -7297 10194 -7263
rect 10228 -7297 10266 -7263
rect 10300 -7297 10337 -7263
rect 10421 -7264 10455 -7234
rect 10421 -7337 10455 -7298
rect 9868 -7371 9906 -7337
rect 9940 -7371 9978 -7337
rect 10012 -7371 10050 -7337
rect 10084 -7371 10122 -7337
rect 10156 -7371 10194 -7337
rect 10228 -7371 10266 -7337
rect 10300 -7371 10337 -7337
rect 10421 -7410 10455 -7371
rect 9868 -7445 9906 -7411
rect 9940 -7445 9978 -7411
rect 10012 -7445 10050 -7411
rect 10084 -7445 10122 -7411
rect 10156 -7445 10194 -7411
rect 10228 -7445 10266 -7411
rect 10300 -7445 10337 -7411
rect 10421 -7483 10455 -7444
rect 9868 -7519 9906 -7485
rect 9940 -7519 9978 -7485
rect 10012 -7519 10050 -7485
rect 10084 -7519 10122 -7485
rect 10156 -7519 10194 -7485
rect 10228 -7519 10266 -7485
rect 10300 -7519 10337 -7485
rect 10421 -7556 10455 -7517
rect 9868 -7593 9906 -7559
rect 9940 -7593 9978 -7559
rect 10012 -7593 10050 -7559
rect 10084 -7593 10122 -7559
rect 10156 -7593 10194 -7559
rect 10228 -7593 10266 -7559
rect 10300 -7593 10337 -7559
rect 9868 -7667 9906 -7633
rect 9940 -7667 9978 -7633
rect 10012 -7667 10050 -7633
rect 10084 -7667 10122 -7633
rect 10156 -7667 10194 -7633
rect 10228 -7667 10266 -7633
rect 10300 -7667 10337 -7633
rect 10421 -7655 10455 -7590
rect 10737 -7264 10771 -7225
rect 11053 -7264 11087 -7225
rect 10851 -7377 10885 -7361
rect 10851 -7519 10885 -7503
rect 10939 -7377 10973 -7361
rect 10939 -7519 10973 -7503
rect 11369 -7264 11403 -7225
rect 10737 -7649 10771 -7593
rect 11167 -7377 11201 -7361
rect 11167 -7519 11201 -7503
rect 11255 -7377 11289 -7361
rect 11255 -7519 11289 -7503
rect 11685 -7264 11719 -7225
rect 11053 -7649 11087 -7593
rect 11483 -7377 11517 -7361
rect 11483 -7519 11517 -7503
rect 11571 -7377 11605 -7361
rect 11571 -7519 11605 -7503
rect 12001 -7264 12035 -7225
rect 11369 -7649 11403 -7593
rect 11799 -7377 11833 -7361
rect 11799 -7519 11833 -7503
rect 11887 -7377 11921 -7361
rect 11887 -7519 11921 -7503
rect 12317 -7264 12351 -7225
rect 11685 -7649 11719 -7593
rect 12115 -7377 12149 -7361
rect 12115 -7519 12149 -7503
rect 12203 -7377 12237 -7361
rect 12203 -7519 12237 -7503
rect 12001 -7649 12035 -7593
rect 12317 -7649 12351 -7593
rect 10737 -7655 10747 -7649
rect 9868 -7741 9906 -7707
rect 9940 -7741 9978 -7707
rect 10012 -7741 10050 -7707
rect 10084 -7741 10122 -7707
rect 10156 -7741 10194 -7707
rect 10228 -7741 10266 -7707
rect 10300 -7741 10337 -7707
rect 4132 -7825 4170 -7791
rect 4204 -7825 4242 -7791
rect 4276 -7825 4314 -7791
rect 4348 -7825 4386 -7791
rect 4420 -7825 4458 -7791
rect 4492 -7825 4530 -7791
rect 4564 -7825 4602 -7791
rect 4636 -7825 4674 -7791
rect 4708 -7825 4746 -7791
rect 4780 -7825 4818 -7791
rect 4852 -7825 4890 -7791
rect 4924 -7825 4962 -7791
rect 4996 -7825 5034 -7791
rect 5068 -7825 5106 -7791
rect 5140 -7825 5178 -7791
rect 5212 -7825 5250 -7791
rect 5284 -7825 5322 -7791
rect 5356 -7825 5394 -7791
rect 5428 -7825 5466 -7791
rect 5500 -7825 5538 -7791
rect 9868 -7815 9906 -7781
rect 9940 -7815 9978 -7781
rect 10012 -7815 10050 -7781
rect 10084 -7815 10122 -7781
rect 10156 -7815 10194 -7781
rect 10228 -7815 10266 -7781
rect 10300 -7815 10338 -7781
rect 10372 -7815 10410 -7781
rect 10444 -7815 10482 -7781
rect 10516 -7815 10554 -7781
rect 4132 -7899 4170 -7865
rect 4204 -7899 4242 -7865
rect 4276 -7899 4314 -7865
rect 4348 -7899 4386 -7865
rect 4420 -7899 4458 -7865
rect 4492 -7899 4530 -7865
rect 4564 -7899 4602 -7865
rect 4636 -7899 4674 -7865
rect 4708 -7899 4746 -7865
rect 4780 -7899 4818 -7865
rect 4852 -7899 4890 -7865
rect 4924 -7899 4962 -7865
rect 4996 -7899 5034 -7865
rect 5068 -7899 5106 -7865
rect 5140 -7899 5178 -7865
rect 5212 -7899 5250 -7865
rect 5284 -7899 5322 -7865
rect 5356 -7899 5394 -7865
rect 5428 -7899 5466 -7865
rect 5500 -7899 5538 -7865
rect 5919 -7875 5935 -7841
rect 5969 -7875 5985 -7841
rect 6037 -7875 6053 -7841
rect 6087 -7875 6103 -7841
rect 6155 -7875 6171 -7841
rect 6205 -7875 6221 -7841
rect 6273 -7875 6289 -7841
rect 6323 -7875 6339 -7841
rect 6391 -7875 6407 -7841
rect 6441 -7875 6457 -7841
rect 6509 -7875 6525 -7841
rect 6559 -7875 6575 -7841
rect 6627 -7875 6643 -7841
rect 6677 -7875 6693 -7841
rect 6745 -7875 6761 -7841
rect 6795 -7875 6811 -7841
rect 6863 -7875 6879 -7841
rect 6913 -7875 6929 -7841
rect 6981 -7875 6997 -7841
rect 7031 -7875 7047 -7841
rect 7099 -7875 7115 -7841
rect 7149 -7875 7165 -7841
rect 7217 -7875 7233 -7841
rect 7267 -7875 7283 -7841
rect 7335 -7875 7351 -7841
rect 7385 -7875 7401 -7841
rect 7453 -7875 7469 -7841
rect 7503 -7875 7519 -7841
rect 7571 -7875 7587 -7841
rect 7621 -7875 7637 -7841
rect 7917 -7875 7933 -7841
rect 7967 -7875 7983 -7841
rect 8035 -7875 8051 -7841
rect 8085 -7875 8101 -7841
rect 8153 -7875 8169 -7841
rect 8203 -7875 8219 -7841
rect 8271 -7875 8287 -7841
rect 8321 -7875 8337 -7841
rect 8389 -7875 8405 -7841
rect 8439 -7875 8455 -7841
rect 8507 -7875 8523 -7841
rect 8557 -7875 8573 -7841
rect 8625 -7875 8641 -7841
rect 8675 -7875 8691 -7841
rect 8743 -7875 8759 -7841
rect 8793 -7875 8809 -7841
rect 8861 -7875 8877 -7841
rect 8911 -7875 8927 -7841
rect 8979 -7875 8995 -7841
rect 9029 -7875 9045 -7841
rect 9097 -7875 9113 -7841
rect 9147 -7875 9163 -7841
rect 9215 -7875 9231 -7841
rect 9265 -7875 9281 -7841
rect 9333 -7875 9349 -7841
rect 9383 -7875 9399 -7841
rect 9451 -7875 9467 -7841
rect 9501 -7875 9517 -7841
rect 9569 -7875 9585 -7841
rect 9619 -7875 9635 -7841
rect 9868 -7889 9906 -7855
rect 9940 -7889 9978 -7855
rect 10012 -7889 10050 -7855
rect 10084 -7889 10122 -7855
rect 10156 -7889 10194 -7855
rect 10228 -7889 10266 -7855
rect 10300 -7889 10338 -7855
rect 10372 -7889 10410 -7855
rect 10444 -7889 10482 -7855
rect 10516 -7889 10554 -7855
rect 4132 -7973 4170 -7939
rect 4204 -7973 4242 -7939
rect 4276 -7973 4314 -7939
rect 4348 -7973 4386 -7939
rect 4420 -7973 4458 -7939
rect 4492 -7973 4530 -7939
rect 4564 -7973 4602 -7939
rect 4636 -7973 4674 -7939
rect 4708 -7973 4746 -7939
rect 4780 -7973 4818 -7939
rect 4852 -7973 4890 -7939
rect 4924 -7973 4962 -7939
rect 4996 -7973 5034 -7939
rect 5068 -7973 5106 -7939
rect 5140 -7973 5178 -7939
rect 5212 -7973 5250 -7939
rect 5284 -7973 5322 -7939
rect 5356 -7973 5394 -7939
rect 5428 -7973 5466 -7939
rect 5500 -7973 5538 -7939
rect 5919 -7983 5935 -7949
rect 5969 -7983 5985 -7949
rect 6037 -7983 6053 -7949
rect 6087 -7983 6103 -7949
rect 6155 -7983 6171 -7949
rect 6205 -7983 6221 -7949
rect 6273 -7983 6289 -7949
rect 6323 -7983 6339 -7949
rect 6391 -7983 6407 -7949
rect 6441 -7983 6457 -7949
rect 6509 -7983 6525 -7949
rect 6559 -7983 6575 -7949
rect 6627 -7983 6643 -7949
rect 6677 -7983 6693 -7949
rect 6745 -7983 6761 -7949
rect 6795 -7983 6811 -7949
rect 6863 -7983 6879 -7949
rect 6913 -7983 6929 -7949
rect 6981 -7983 6997 -7949
rect 7031 -7983 7047 -7949
rect 7099 -7983 7115 -7949
rect 7149 -7983 7165 -7949
rect 7217 -7983 7233 -7949
rect 7267 -7983 7283 -7949
rect 7335 -7983 7351 -7949
rect 7385 -7983 7401 -7949
rect 7453 -7983 7469 -7949
rect 7503 -7983 7519 -7949
rect 7571 -7983 7587 -7949
rect 7621 -7983 7637 -7949
rect 7917 -7983 7933 -7949
rect 7967 -7983 7983 -7949
rect 8035 -7983 8051 -7949
rect 8085 -7983 8101 -7949
rect 8153 -7983 8169 -7949
rect 8203 -7983 8219 -7949
rect 8271 -7983 8287 -7949
rect 8321 -7983 8337 -7949
rect 8389 -7983 8405 -7949
rect 8439 -7983 8455 -7949
rect 8507 -7983 8523 -7949
rect 8557 -7983 8573 -7949
rect 8625 -7983 8641 -7949
rect 8675 -7983 8691 -7949
rect 8743 -7983 8759 -7949
rect 8793 -7983 8809 -7949
rect 8861 -7983 8877 -7949
rect 8911 -7983 8927 -7949
rect 8979 -7983 8995 -7949
rect 9029 -7983 9045 -7949
rect 9097 -7983 9113 -7949
rect 9147 -7983 9163 -7949
rect 9215 -7983 9231 -7949
rect 9265 -7983 9281 -7949
rect 9333 -7983 9349 -7949
rect 9383 -7983 9399 -7949
rect 9451 -7983 9467 -7949
rect 9501 -7983 9517 -7949
rect 9569 -7983 9585 -7949
rect 9619 -7983 9635 -7949
rect 9868 -7963 9906 -7929
rect 9940 -7963 9978 -7929
rect 10012 -7963 10050 -7929
rect 10084 -7963 10122 -7929
rect 10156 -7963 10194 -7929
rect 10228 -7963 10266 -7929
rect 10300 -7963 10338 -7929
rect 10372 -7963 10410 -7929
rect 10444 -7963 10482 -7929
rect 4132 -8047 4170 -8013
rect 4204 -8047 4242 -8013
rect 4276 -8047 4314 -8013
rect 4348 -8047 4386 -8013
rect 4420 -8047 4458 -8013
rect 4492 -8047 4530 -8013
rect 4564 -8047 4602 -8013
rect 4636 -8047 4674 -8013
rect 4708 -8047 4746 -8013
rect 4780 -8047 4818 -8013
rect 4852 -8047 4890 -8013
rect 4924 -8047 4962 -8013
rect 4996 -8047 5034 -8013
rect 5068 -8047 5106 -8013
rect 5140 -8047 5178 -8013
rect 5212 -8047 5250 -8013
rect 5284 -8047 5322 -8013
rect 5356 -8047 5394 -8013
rect 5428 -8047 5466 -8013
rect 5500 -8047 5538 -8013
rect 4132 -8121 4170 -8087
rect 4204 -8121 4242 -8087
rect 4276 -8121 4314 -8087
rect 4348 -8121 4386 -8087
rect 4420 -8121 4458 -8087
rect 4492 -8121 4530 -8087
rect 4564 -8121 4602 -8087
rect 4636 -8121 4674 -8087
rect 4708 -8121 4746 -8087
rect 4780 -8121 4818 -8087
rect 4852 -8121 4890 -8087
rect 4924 -8121 4962 -8087
rect 4996 -8121 5034 -8087
rect 5068 -8121 5106 -8087
rect 5140 -8121 5178 -8087
rect 5212 -8121 5250 -8087
rect 5284 -8121 5322 -8087
rect 5356 -8121 5394 -8087
rect 5428 -8121 5466 -8087
rect 5500 -8121 5538 -8087
rect 4132 -8195 4170 -8161
rect 4204 -8195 4242 -8161
rect 4276 -8195 4314 -8161
rect 4348 -8195 4386 -8161
rect 4420 -8195 4458 -8161
rect 4492 -8195 4530 -8161
rect 4564 -8195 4602 -8161
rect 4636 -8195 4674 -8161
rect 4708 -8195 4746 -8161
rect 4780 -8195 4818 -8161
rect 4852 -8195 4890 -8161
rect 4924 -8195 4962 -8161
rect 4996 -8195 5034 -8161
rect 5068 -8195 5106 -8161
rect 5140 -8195 5178 -8161
rect 5212 -8195 5250 -8161
rect 5284 -8195 5322 -8161
rect 5356 -8195 5394 -8161
rect 5428 -8195 5466 -8161
rect 5500 -8195 5538 -8161
rect 4132 -8269 4170 -8235
rect 4204 -8269 4242 -8235
rect 4276 -8269 4314 -8235
rect 4348 -8269 4386 -8235
rect 4420 -8269 4458 -8235
rect 4492 -8269 4530 -8235
rect 4564 -8269 4602 -8235
rect 4636 -8269 4674 -8235
rect 4708 -8269 4746 -8235
rect 4780 -8269 4818 -8235
rect 4852 -8269 4890 -8235
rect 4924 -8269 4962 -8235
rect 4996 -8269 5034 -8235
rect 5068 -8269 5106 -8235
rect 5140 -8269 5178 -8235
rect 5212 -8269 5250 -8235
rect 5284 -8269 5322 -8235
rect 5356 -8269 5394 -8235
rect 5428 -8269 5466 -8235
rect 5500 -8269 5538 -8235
rect 4132 -8343 4170 -8309
rect 4204 -8343 4242 -8309
rect 4276 -8343 4314 -8309
rect 4348 -8343 4386 -8309
rect 4420 -8343 4458 -8309
rect 4492 -8343 4530 -8309
rect 4564 -8343 4602 -8309
rect 4636 -8343 4674 -8309
rect 4708 -8343 4746 -8309
rect 4780 -8343 4818 -8309
rect 4852 -8343 4890 -8309
rect 4924 -8343 4962 -8309
rect 4996 -8343 5034 -8309
rect 5068 -8343 5106 -8309
rect 5140 -8343 5178 -8309
rect 5212 -8343 5250 -8309
rect 5284 -8343 5322 -8309
rect 5356 -8343 5394 -8309
rect 5428 -8343 5466 -8309
rect 5500 -8343 5538 -8309
rect 4132 -8417 4170 -8383
rect 4204 -8417 4242 -8383
rect 4276 -8417 4314 -8383
rect 4348 -8417 4386 -8383
rect 4420 -8417 4458 -8383
rect 4492 -8417 4530 -8383
rect 4564 -8417 4602 -8383
rect 4636 -8417 4674 -8383
rect 4708 -8417 4746 -8383
rect 4780 -8417 4818 -8383
rect 4852 -8417 4890 -8383
rect 4924 -8417 4962 -8383
rect 4996 -8417 5034 -8383
rect 5068 -8417 5106 -8383
rect 5140 -8417 5178 -8383
rect 5212 -8417 5250 -8383
rect 5284 -8417 5322 -8383
rect 5356 -8417 5394 -8383
rect 5428 -8417 5466 -8383
rect 5500 -8417 5538 -8383
rect 4132 -8491 4170 -8457
rect 4204 -8491 4242 -8457
rect 4276 -8491 4314 -8457
rect 4348 -8491 4386 -8457
rect 4420 -8491 4458 -8457
rect 4492 -8491 4530 -8457
rect 4564 -8491 4602 -8457
rect 4636 -8491 4674 -8457
rect 4708 -8491 4746 -8457
rect 4780 -8491 4818 -8457
rect 4852 -8491 4890 -8457
rect 4924 -8491 4962 -8457
rect 4996 -8491 5034 -8457
rect 5068 -8491 5106 -8457
rect 5140 -8491 5178 -8457
rect 5212 -8491 5250 -8457
rect 5284 -8491 5322 -8457
rect 5356 -8491 5394 -8457
rect 5428 -8491 5466 -8457
rect 5500 -8491 5538 -8457
rect 4132 -8565 4170 -8531
rect 4204 -8565 4242 -8531
rect 4276 -8565 4314 -8531
rect 4348 -8565 4386 -8531
rect 4420 -8565 4458 -8531
rect 4492 -8565 4530 -8531
rect 4564 -8565 4602 -8531
rect 4636 -8565 4674 -8531
rect 4708 -8565 4746 -8531
rect 4780 -8565 4818 -8531
rect 4852 -8565 4890 -8531
rect 4924 -8565 4962 -8531
rect 4996 -8565 5034 -8531
rect 5068 -8565 5106 -8531
rect 5140 -8565 5178 -8531
rect 5212 -8565 5250 -8531
rect 5284 -8565 5322 -8531
rect 5356 -8565 5394 -8531
rect 5428 -8565 5466 -8531
rect 5500 -8565 5538 -8531
rect 9868 -8037 9906 -8003
rect 9940 -8037 9978 -8003
rect 10012 -8037 10050 -8003
rect 10084 -8037 10122 -8003
rect 10156 -8037 10194 -8003
rect 10228 -8037 10266 -8003
rect 10300 -8037 10338 -8003
rect 10372 -8037 10410 -8003
rect 10444 -8037 10482 -8003
rect 9868 -8111 9906 -8077
rect 9940 -8111 9978 -8077
rect 10012 -8111 10050 -8077
rect 10084 -8111 10122 -8077
rect 10156 -8111 10194 -8077
rect 10228 -8111 10266 -8077
rect 10300 -8111 10338 -8077
rect 10372 -8111 10410 -8077
rect 10444 -8111 10482 -8077
rect 9868 -8185 9906 -8151
rect 9940 -8185 9978 -8151
rect 10012 -8185 10050 -8151
rect 10084 -8185 10122 -8151
rect 10156 -8185 10194 -8151
rect 10228 -8185 10266 -8151
rect 10300 -8185 10338 -8151
rect 10372 -8185 10410 -8151
rect 10444 -8185 10482 -8151
rect 12728 -8175 12744 -8141
rect 12802 -8175 12818 -8141
rect 12876 -8175 12892 -8141
rect 12950 -8175 12966 -8141
rect 13024 -8175 13040 -8141
rect 13098 -8175 13114 -8141
rect 13172 -8175 13188 -8141
rect 13246 -8175 13262 -8141
rect 13320 -8175 13336 -8141
rect 13394 -8175 13410 -8141
rect 13468 -8175 13484 -8141
rect 13542 -8175 13558 -8141
rect 13616 -8175 13632 -8141
rect 13690 -8175 13706 -8141
rect 13764 -8175 13780 -8141
rect 13838 -8175 13854 -8141
rect 13912 -8175 13928 -8141
rect 13986 -8175 14002 -8141
rect 14060 -8175 14076 -8141
rect 14134 -8175 14150 -8141
rect 14208 -8175 14224 -8141
rect 14282 -8175 14298 -8141
rect 14356 -8175 14372 -8141
rect 14430 -8175 14446 -8141
rect 14504 -8175 14520 -8141
rect 14578 -8175 14594 -8141
rect 14652 -8175 14668 -8141
rect 14726 -8175 14742 -8141
rect 14800 -8175 14816 -8141
rect 14874 -8175 14890 -8141
rect 14948 -8175 14964 -8141
rect 15022 -8175 15038 -8141
rect 15096 -8175 15112 -8141
rect 15170 -8175 15186 -8141
rect 15244 -8175 15260 -8141
rect 15318 -8175 15334 -8141
rect 15392 -8175 15408 -8141
rect 15466 -8175 15482 -8141
rect 15540 -8175 15556 -8141
rect 15614 -8175 15630 -8141
rect 15688 -8175 15704 -8141
rect 15762 -8175 15778 -8141
rect 15836 -8175 15852 -8141
rect 15910 -8175 15926 -8141
rect 15984 -8175 16000 -8141
rect 16058 -8175 16074 -8141
rect 16132 -8175 16148 -8141
rect 16206 -8175 16222 -8141
rect 16280 -8175 16296 -8141
rect 16354 -8175 16370 -8141
rect 16428 -8175 16444 -8141
rect 16502 -8175 16518 -8141
rect 16576 -8175 16592 -8141
rect 16650 -8175 16666 -8141
rect 16724 -8175 16740 -8141
rect 16798 -8175 16814 -8141
rect 16872 -8175 16888 -8141
rect 16946 -8175 16962 -8141
rect 17020 -8175 17036 -8141
rect 17094 -8175 17110 -8141
rect 17168 -8175 17184 -8141
rect 17242 -8175 17258 -8141
rect 17316 -8175 17332 -8141
rect 17390 -8175 17406 -8141
rect 17464 -8175 17480 -8141
rect 17538 -8175 17554 -8141
rect 17612 -8175 17628 -8141
rect 17686 -8175 17702 -8141
rect 17760 -8175 17776 -8141
rect 17834 -8175 17850 -8141
rect 17908 -8175 17924 -8141
rect 17982 -8175 17998 -8141
rect 18056 -8175 18072 -8141
rect 18130 -8175 18146 -8141
rect 18204 -8175 18220 -8141
rect 18278 -8175 18294 -8141
rect 18352 -8175 18368 -8141
rect 18426 -8175 18442 -8141
rect 18500 -8175 18516 -8141
rect 18574 -8175 18590 -8141
rect 18648 -8175 18664 -8141
rect 18722 -8175 18738 -8141
rect 18796 -8175 18812 -8141
rect 18870 -8175 18886 -8141
rect 18944 -8175 18960 -8141
rect 19018 -8175 19034 -8141
rect 19092 -8175 19108 -8141
rect 19166 -8175 19182 -8141
rect 19240 -8175 19256 -8141
rect 19314 -8175 19330 -8141
rect 19388 -8175 19404 -8141
rect 19462 -8175 19478 -8141
rect 19536 -8175 19552 -8141
rect 19610 -8175 19626 -8141
rect 19684 -8175 19700 -8141
rect 19758 -8175 19774 -8141
rect 19832 -8175 19848 -8141
rect 19906 -8175 19922 -8141
rect 19980 -8175 19996 -8141
rect 20054 -8175 20070 -8141
rect 20128 -8175 20144 -8141
rect 20202 -8175 20218 -8141
rect 20276 -8175 20292 -8141
rect 20350 -8175 20366 -8141
rect 20424 -8175 20440 -8141
rect 20498 -8175 20514 -8141
rect 20572 -8175 20588 -8141
rect 20646 -8175 20662 -8141
rect 20720 -8175 20736 -8141
rect 20794 -8175 20810 -8141
rect 20868 -8175 20884 -8141
rect 20942 -8175 20958 -8141
rect 21016 -8175 21032 -8141
rect 21090 -8175 21106 -8141
rect 21164 -8175 21180 -8141
rect 21238 -8175 21254 -8141
rect 21312 -8175 21328 -8141
rect 21386 -8175 21402 -8141
rect 21460 -8175 21476 -8141
rect 21534 -8175 21550 -8141
rect 21608 -8175 21624 -8141
rect 21682 -8175 21698 -8141
rect 21756 -8175 21772 -8141
rect 21830 -8175 21846 -8141
rect 21904 -8175 21920 -8141
rect 21978 -8175 21994 -8141
rect 22052 -8175 22068 -8141
rect 22126 -8175 22142 -8141
rect 22200 -8175 22216 -8141
rect 22274 -8175 22290 -8141
rect 22348 -8175 22364 -8141
rect 22422 -8175 22438 -8141
rect 22496 -8175 22512 -8141
rect 22570 -8175 22586 -8141
rect 22644 -8175 22660 -8141
rect 22718 -8175 22734 -8141
rect 22792 -8175 22808 -8141
rect 22866 -8175 22882 -8141
rect 22940 -8175 22956 -8141
rect 23014 -8175 23030 -8141
rect 23088 -8175 23104 -8141
rect 23162 -8175 23178 -8141
rect 23236 -8175 23252 -8141
rect 23310 -8175 23326 -8141
rect 23384 -8175 23400 -8141
rect 23458 -8175 23474 -8141
rect 23532 -8175 23548 -8141
rect 23606 -8175 23622 -8141
rect 9868 -8259 9906 -8225
rect 9940 -8259 9978 -8225
rect 10012 -8259 10050 -8225
rect 10084 -8259 10122 -8225
rect 10156 -8259 10194 -8225
rect 10228 -8259 10266 -8225
rect 10300 -8259 10338 -8225
rect 10372 -8259 10410 -8225
rect 10444 -8259 10482 -8225
rect 12728 -8283 12744 -8249
rect 12802 -8283 12818 -8249
rect 12876 -8283 12892 -8249
rect 12950 -8283 12966 -8249
rect 13024 -8283 13040 -8249
rect 13098 -8283 13114 -8249
rect 13172 -8283 13188 -8249
rect 13246 -8283 13262 -8249
rect 13320 -8283 13336 -8249
rect 13394 -8283 13410 -8249
rect 13468 -8283 13484 -8249
rect 13542 -8283 13558 -8249
rect 13616 -8283 13632 -8249
rect 13690 -8283 13706 -8249
rect 13764 -8283 13780 -8249
rect 13838 -8283 13854 -8249
rect 13912 -8283 13928 -8249
rect 13986 -8283 14002 -8249
rect 14060 -8283 14076 -8249
rect 14134 -8283 14150 -8249
rect 14208 -8283 14224 -8249
rect 14282 -8283 14298 -8249
rect 14356 -8283 14372 -8249
rect 14430 -8283 14446 -8249
rect 14504 -8283 14520 -8249
rect 14578 -8283 14594 -8249
rect 14652 -8283 14668 -8249
rect 14726 -8283 14742 -8249
rect 14800 -8283 14816 -8249
rect 14874 -8283 14890 -8249
rect 14948 -8283 14964 -8249
rect 15022 -8283 15038 -8249
rect 15096 -8283 15112 -8249
rect 15170 -8283 15186 -8249
rect 15244 -8283 15260 -8249
rect 15318 -8283 15334 -8249
rect 15392 -8283 15408 -8249
rect 15466 -8283 15482 -8249
rect 15540 -8283 15556 -8249
rect 15614 -8283 15630 -8249
rect 15688 -8283 15704 -8249
rect 15762 -8283 15778 -8249
rect 15836 -8283 15852 -8249
rect 15910 -8283 15926 -8249
rect 15984 -8283 16000 -8249
rect 16058 -8283 16074 -8249
rect 16132 -8283 16148 -8249
rect 16206 -8283 16222 -8249
rect 16280 -8283 16296 -8249
rect 16354 -8283 16370 -8249
rect 16428 -8283 16444 -8249
rect 16502 -8283 16518 -8249
rect 16576 -8283 16592 -8249
rect 16650 -8283 16666 -8249
rect 16724 -8283 16740 -8249
rect 16798 -8283 16814 -8249
rect 16872 -8283 16888 -8249
rect 16946 -8283 16962 -8249
rect 17020 -8283 17036 -8249
rect 17094 -8283 17110 -8249
rect 17168 -8283 17184 -8249
rect 17242 -8283 17258 -8249
rect 17316 -8283 17332 -8249
rect 17390 -8283 17406 -8249
rect 17464 -8283 17480 -8249
rect 17538 -8283 17554 -8249
rect 17612 -8283 17628 -8249
rect 17686 -8283 17702 -8249
rect 17760 -8283 17776 -8249
rect 17834 -8283 17850 -8249
rect 17908 -8283 17924 -8249
rect 17982 -8283 17998 -8249
rect 18056 -8283 18072 -8249
rect 18130 -8283 18146 -8249
rect 18204 -8283 18220 -8249
rect 18278 -8283 18294 -8249
rect 18352 -8283 18368 -8249
rect 18426 -8283 18442 -8249
rect 18500 -8283 18516 -8249
rect 18574 -8283 18590 -8249
rect 18648 -8283 18664 -8249
rect 18722 -8283 18738 -8249
rect 18796 -8283 18812 -8249
rect 18870 -8283 18886 -8249
rect 18944 -8283 18960 -8249
rect 19018 -8283 19034 -8249
rect 19092 -8283 19108 -8249
rect 19166 -8283 19182 -8249
rect 19240 -8283 19256 -8249
rect 19314 -8283 19330 -8249
rect 19388 -8283 19404 -8249
rect 19462 -8283 19478 -8249
rect 19536 -8283 19552 -8249
rect 19610 -8283 19626 -8249
rect 19684 -8283 19700 -8249
rect 19758 -8283 19774 -8249
rect 19832 -8283 19848 -8249
rect 19906 -8283 19922 -8249
rect 19980 -8283 19996 -8249
rect 20054 -8283 20070 -8249
rect 20128 -8283 20144 -8249
rect 20202 -8283 20218 -8249
rect 20276 -8283 20292 -8249
rect 20350 -8283 20366 -8249
rect 20424 -8283 20440 -8249
rect 20498 -8283 20514 -8249
rect 20572 -8283 20588 -8249
rect 20646 -8283 20662 -8249
rect 20720 -8283 20736 -8249
rect 20794 -8283 20810 -8249
rect 20868 -8283 20884 -8249
rect 20942 -8283 20958 -8249
rect 21016 -8283 21032 -8249
rect 21090 -8283 21106 -8249
rect 21164 -8283 21180 -8249
rect 21238 -8283 21254 -8249
rect 21312 -8283 21328 -8249
rect 21386 -8283 21402 -8249
rect 21460 -8283 21476 -8249
rect 21534 -8283 21550 -8249
rect 21608 -8283 21624 -8249
rect 21682 -8283 21698 -8249
rect 21756 -8283 21772 -8249
rect 21830 -8283 21846 -8249
rect 21904 -8283 21920 -8249
rect 21978 -8283 21994 -8249
rect 22052 -8283 22068 -8249
rect 22126 -8283 22142 -8249
rect 22200 -8283 22216 -8249
rect 22274 -8283 22290 -8249
rect 22348 -8283 22364 -8249
rect 22422 -8283 22438 -8249
rect 22496 -8283 22512 -8249
rect 22570 -8283 22586 -8249
rect 22644 -8283 22660 -8249
rect 22718 -8283 22734 -8249
rect 22792 -8283 22808 -8249
rect 22866 -8283 22882 -8249
rect 22940 -8283 22956 -8249
rect 23014 -8283 23030 -8249
rect 23088 -8283 23104 -8249
rect 23162 -8283 23178 -8249
rect 23236 -8283 23252 -8249
rect 23310 -8283 23326 -8249
rect 23384 -8283 23400 -8249
rect 23458 -8283 23474 -8249
rect 23532 -8283 23548 -8249
rect 23606 -8283 23622 -8249
rect 9868 -8333 9906 -8299
rect 9940 -8333 9978 -8299
rect 10012 -8333 10050 -8299
rect 10084 -8333 10122 -8299
rect 10156 -8333 10194 -8299
rect 10228 -8333 10266 -8299
rect 10300 -8333 10338 -8299
rect 10372 -8333 10410 -8299
rect 10444 -8333 10482 -8299
rect 10516 -8333 10554 -8299
rect 9868 -8407 9906 -8373
rect 9940 -8407 9978 -8373
rect 10012 -8407 10050 -8373
rect 10084 -8407 10122 -8373
rect 10156 -8407 10194 -8373
rect 10228 -8407 10266 -8373
rect 10300 -8407 10338 -8373
rect 10372 -8407 10410 -8373
rect 10444 -8407 10482 -8373
rect 10516 -8407 10554 -8373
rect 9868 -8481 9906 -8447
rect 9940 -8481 9978 -8447
rect 10012 -8481 10050 -8447
rect 10084 -8481 10122 -8447
rect 10156 -8481 10194 -8447
rect 10228 -8481 10266 -8447
rect 10300 -8481 10338 -8447
rect 10372 -8481 10410 -8447
rect 10444 -8481 10482 -8447
rect 10516 -8481 10554 -8447
rect 9868 -8555 9906 -8521
rect 9940 -8555 9978 -8521
rect 10012 -8555 10050 -8521
rect 10084 -8555 10122 -8521
rect 10156 -8555 10194 -8521
rect 10228 -8555 10266 -8521
rect 10300 -8555 10338 -8521
rect 10372 -8555 10410 -8521
rect 10444 -8555 10482 -8521
rect 10516 -8555 10554 -8521
rect 9868 -8629 9906 -8595
rect 9940 -8629 9978 -8595
rect 10012 -8629 10050 -8595
rect 10084 -8629 10122 -8595
rect 10156 -8629 10194 -8595
rect 10228 -8629 10266 -8595
rect 10300 -8629 10338 -8595
rect 10372 -8629 10410 -8595
rect 10444 -8629 10482 -8595
rect 10516 -8629 10554 -8595
rect 9868 -8703 9906 -8669
rect 9940 -8703 9978 -8669
rect 10012 -8703 10050 -8669
rect 10084 -8703 10122 -8669
rect 10156 -8703 10194 -8669
rect 10228 -8703 10266 -8669
rect 10300 -8703 10338 -8669
rect 10372 -8703 10410 -8669
rect 10444 -8703 10482 -8669
rect 10516 -8703 10554 -8669
rect 4020 -9712 4060 -9678
rect 4094 -9712 4134 -9678
rect 4168 -9712 4208 -9678
rect 4242 -9712 4282 -9678
rect 4316 -9712 4356 -9678
rect 4390 -9712 4430 -9678
rect 4464 -9712 4504 -9678
rect 4538 -9712 4578 -9678
rect 4612 -9712 4652 -9678
rect 4686 -9712 4726 -9678
rect 4760 -9712 4800 -9678
rect 4834 -9712 4874 -9678
rect 4908 -9712 4948 -9678
rect 4982 -9712 5022 -9678
rect 5056 -9712 5096 -9678
rect 5130 -9712 5170 -9678
rect 5204 -9712 5244 -9678
rect 5278 -9712 5318 -9678
rect 5352 -9712 5392 -9678
rect 5426 -9712 5466 -9678
rect 5500 -9712 5540 -9678
rect 5574 -9712 5614 -9678
rect 5648 -9712 5688 -9678
rect 5722 -9712 5762 -9678
rect 5796 -9712 5836 -9678
rect 5870 -9712 5910 -9678
rect 5944 -9712 5984 -9678
rect 6018 -9712 6058 -9678
rect 6092 -9712 6132 -9678
rect 6166 -9712 6206 -9678
rect 6240 -9712 6280 -9678
rect 6314 -9712 6354 -9678
rect 6388 -9712 6428 -9678
rect 6462 -9712 6502 -9678
rect 6536 -9712 6576 -9678
rect 6610 -9712 6650 -9678
rect 6684 -9712 6724 -9678
rect 6758 -9712 6798 -9678
rect 6832 -9712 6872 -9678
rect 6906 -9712 6946 -9678
rect 6980 -9712 7020 -9678
rect 7054 -9712 7094 -9678
rect 7128 -9712 7168 -9678
rect 7202 -9712 7242 -9678
rect 7276 -9712 7316 -9678
rect 7350 -9712 7390 -9678
rect 7424 -9712 7464 -9678
rect 7498 -9712 7538 -9678
rect 7572 -9712 7612 -9678
rect 7646 -9712 7686 -9678
rect 7720 -9712 7760 -9678
rect 7794 -9712 7834 -9678
rect 7868 -9712 7908 -9678
rect 7942 -9712 7982 -9678
rect 8016 -9712 8056 -9678
rect 8090 -9712 8130 -9678
rect 8164 -9712 8204 -9678
rect 8238 -9712 8278 -9678
rect 8312 -9712 8352 -9678
rect 8386 -9712 8426 -9678
rect 8460 -9712 8500 -9678
rect 8534 -9712 8574 -9678
rect 8608 -9712 8648 -9678
rect 8682 -9712 8722 -9678
rect 8756 -9712 8796 -9678
rect 8830 -9712 8870 -9678
rect 8904 -9712 8944 -9678
rect 8978 -9712 9018 -9678
rect 9052 -9712 9092 -9678
rect 9126 -9712 9166 -9678
rect 9200 -9712 9240 -9678
rect 9274 -9712 9314 -9678
rect 9348 -9712 9388 -9678
rect 9422 -9712 9462 -9678
rect 9496 -9712 9536 -9678
rect 9570 -9712 9610 -9678
rect 9644 -9712 9684 -9678
rect 9718 -9712 9758 -9678
rect 9792 -9712 9832 -9678
rect 9866 -9712 9906 -9678
rect 9940 -9712 9980 -9678
rect 10014 -9712 10054 -9678
rect 10088 -9712 10128 -9678
rect 10162 -9712 10202 -9678
rect 10236 -9712 10276 -9678
rect 10310 -9712 10350 -9678
rect 10384 -9712 10424 -9678
rect 10458 -9712 10498 -9678
rect 10532 -9712 10572 -9678
rect 10606 -9712 10646 -9678
rect 10680 -9712 10720 -9678
rect 10754 -9712 10794 -9678
rect 10828 -9712 10868 -9678
rect 10902 -9712 10942 -9678
rect 10976 -9712 11016 -9678
rect 11050 -9712 11090 -9678
rect 11124 -9712 11164 -9678
rect 11198 -9712 11238 -9678
rect 11272 -9712 11312 -9678
rect 11346 -9712 11386 -9678
rect 11420 -9712 11460 -9678
rect 11494 -9712 11534 -9678
rect 11568 -9712 11608 -9678
rect 11642 -9712 11682 -9678
rect 11716 -9712 11756 -9678
rect 11790 -9712 11830 -9678
rect 11864 -9712 11904 -9678
rect 11938 -9712 11978 -9678
rect 12012 -9712 12052 -9678
rect 12086 -9712 12126 -9678
rect 12160 -9712 12200 -9678
rect 12234 -9712 12274 -9678
rect 12308 -9712 12348 -9678
rect 12382 -9712 12422 -9678
rect 12456 -9712 12496 -9678
rect 12530 -9712 12570 -9678
rect 12604 -9712 12644 -9678
rect 12678 -9712 12718 -9678
rect 12752 -9712 12792 -9678
rect 12826 -9712 12866 -9678
rect 12900 -9712 12940 -9678
rect 12974 -9712 13014 -9678
rect 13048 -9712 13088 -9678
rect 13122 -9712 13162 -9678
rect 13196 -9712 13236 -9678
rect 13270 -9712 13310 -9678
rect 13344 -9712 13384 -9678
rect 13418 -9712 13458 -9678
rect 13492 -9712 13532 -9678
rect 13566 -9712 13606 -9678
rect 13640 -9712 13680 -9678
rect 13714 -9712 13754 -9678
rect 13788 -9712 13828 -9678
rect 13862 -9712 13902 -9678
rect 13936 -9712 13976 -9678
rect 14010 -9712 14050 -9678
rect 14084 -9712 14124 -9678
rect 14158 -9712 14198 -9678
rect 14232 -9712 14272 -9678
rect 14306 -9712 14346 -9678
rect 14380 -9712 14420 -9678
rect 14454 -9712 14494 -9678
rect 14528 -9712 14568 -9678
rect 14602 -9712 14642 -9678
rect 14676 -9712 14716 -9678
rect 14750 -9712 14790 -9678
rect 14824 -9712 14864 -9678
rect 14898 -9712 14938 -9678
rect 14972 -9712 15012 -9678
rect 15046 -9712 15086 -9678
rect 15120 -9712 15160 -9678
rect 15194 -9712 15234 -9678
rect 15268 -9712 15308 -9678
rect 15342 -9712 15382 -9678
rect 15416 -9712 15456 -9678
rect 15490 -9712 15530 -9678
rect 15564 -9712 15604 -9678
rect 15638 -9712 15678 -9678
rect 15712 -9712 15752 -9678
rect 15786 -9712 15826 -9678
rect 15860 -9712 15900 -9678
rect 15934 -9712 15974 -9678
rect 16008 -9712 16048 -9678
rect 16082 -9712 16122 -9678
rect 16156 -9712 16196 -9678
rect 16230 -9712 16270 -9678
rect 16304 -9712 16344 -9678
rect 16378 -9712 16418 -9678
rect 16452 -9712 16492 -9678
rect 16526 -9712 16566 -9678
rect 16600 -9712 16640 -9678
rect 16674 -9712 16714 -9678
rect 16748 -9712 16788 -9678
rect 16822 -9712 16862 -9678
rect 16896 -9712 16936 -9678
rect 16970 -9712 17010 -9678
rect 17044 -9712 17084 -9678
rect 17118 -9712 17158 -9678
rect 17192 -9712 17232 -9678
rect 17266 -9712 17306 -9678
rect 17340 -9712 17380 -9678
rect 17414 -9712 17454 -9678
rect 17488 -9712 17528 -9678
rect 17562 -9712 17602 -9678
rect 17636 -9712 17676 -9678
rect 17710 -9712 17750 -9678
rect 17784 -9712 17824 -9678
rect 17858 -9712 17898 -9678
rect 17932 -9712 17972 -9678
rect 18006 -9712 18046 -9678
rect 18080 -9712 18120 -9678
rect 18154 -9712 18194 -9678
rect 18228 -9712 18268 -9678
rect 18302 -9712 18342 -9678
rect 18376 -9712 18416 -9678
rect 18450 -9712 18490 -9678
rect 18524 -9712 18564 -9678
rect 18598 -9712 18638 -9678
rect 18672 -9712 18712 -9678
rect 18746 -9712 18786 -9678
rect 18820 -9712 18860 -9678
rect 18894 -9712 18934 -9678
rect 18968 -9712 19008 -9678
rect 19042 -9712 19082 -9678
rect 19116 -9712 19156 -9678
rect 19190 -9712 19230 -9678
rect 19264 -9712 19304 -9678
rect 19338 -9712 19378 -9678
rect 19412 -9712 19452 -9678
rect 19486 -9712 19526 -9678
rect 19560 -9712 19600 -9678
rect 19634 -9712 19674 -9678
rect 19708 -9712 19748 -9678
rect 19782 -9712 19822 -9678
rect 19856 -9712 19896 -9678
rect 19930 -9712 19970 -9678
rect 20004 -9712 20044 -9678
rect 20078 -9712 20118 -9678
rect 20152 -9712 20192 -9678
rect 20226 -9712 20266 -9678
rect 20300 -9712 20340 -9678
rect 20374 -9712 20414 -9678
rect 20448 -9712 20488 -9678
rect 20522 -9712 20562 -9678
rect 20596 -9712 20636 -9678
rect 20670 -9712 20710 -9678
rect 20744 -9712 20784 -9678
rect 20818 -9712 20858 -9678
rect 20892 -9712 20932 -9678
rect 20966 -9712 21006 -9678
rect 21040 -9712 21080 -9678
rect 21114 -9712 21154 -9678
rect 21188 -9712 21228 -9678
rect 21262 -9712 21302 -9678
rect 21336 -9712 21376 -9678
rect 21410 -9712 21450 -9678
rect 21484 -9712 21524 -9678
rect 21558 -9712 21598 -9678
rect 21632 -9712 21672 -9678
rect 21706 -9712 21746 -9678
rect 21780 -9712 21820 -9678
rect 21854 -9712 21894 -9678
rect 21928 -9712 21968 -9678
rect 22002 -9712 22042 -9678
rect 22076 -9712 22116 -9678
rect 22150 -9712 22190 -9678
rect 22224 -9712 22264 -9678
rect 22298 -9712 22338 -9678
rect 22372 -9712 22412 -9678
rect 22446 -9712 22486 -9678
rect 22520 -9712 22560 -9678
rect 22594 -9712 22634 -9678
rect 22668 -9712 22708 -9678
rect 22742 -9712 22782 -9678
rect 22816 -9712 22856 -9678
rect 22890 -9712 22930 -9678
rect 22964 -9712 23004 -9678
rect 23038 -9712 23078 -9678
rect 23112 -9712 23152 -9678
rect 23186 -9712 23226 -9678
rect 23260 -9712 23300 -9678
rect 23334 -9712 23374 -9678
rect 23408 -9712 23448 -9678
rect 23482 -9712 23522 -9678
rect 23556 -9712 23596 -9678
rect 23630 -9712 23670 -9678
rect 23704 -9712 23744 -9678
rect 23778 -9712 23818 -9678
rect 23852 -9712 23892 -9678
rect 23926 -9712 23966 -9678
rect 24000 -9712 24040 -9678
rect 24074 -9712 24114 -9678
rect 24148 -9712 24188 -9678
rect 24222 -9712 24262 -9678
rect 24296 -9712 24336 -9678
rect 24370 -9712 24410 -9678
rect 24444 -9712 24484 -9678
rect 24518 -9712 24558 -9678
rect 24592 -9712 24632 -9678
rect 24666 -9712 24706 -9678
rect 24740 -9712 24780 -9678
rect 24814 -9712 24854 -9678
rect 24888 -9712 24928 -9678
rect 24962 -9712 25002 -9678
rect 25036 -9712 25076 -9678
rect 25110 -9712 25150 -9678
rect 25184 -9712 26250 -9678
rect 4020 -9786 4060 -9752
rect 4094 -9786 4134 -9752
rect 4168 -9786 4208 -9752
rect 4242 -9786 4282 -9752
rect 4316 -9786 4356 -9752
rect 4390 -9786 4430 -9752
rect 4464 -9786 4504 -9752
rect 4538 -9786 4578 -9752
rect 4612 -9786 4652 -9752
rect 4686 -9786 4726 -9752
rect 4760 -9786 4800 -9752
rect 4834 -9786 4874 -9752
rect 4908 -9786 4948 -9752
rect 4982 -9786 5022 -9752
rect 5056 -9786 5096 -9752
rect 5130 -9786 5170 -9752
rect 5204 -9786 5244 -9752
rect 5278 -9786 5318 -9752
rect 5352 -9786 5392 -9752
rect 5426 -9786 5466 -9752
rect 5500 -9786 5540 -9752
rect 5574 -9786 5614 -9752
rect 5648 -9786 5688 -9752
rect 5722 -9786 5762 -9752
rect 5796 -9786 5836 -9752
rect 5870 -9786 5910 -9752
rect 5944 -9786 5984 -9752
rect 6018 -9786 6058 -9752
rect 6092 -9786 6132 -9752
rect 6166 -9786 6206 -9752
rect 6240 -9786 6280 -9752
rect 6314 -9786 6354 -9752
rect 6388 -9786 6428 -9752
rect 6462 -9786 6502 -9752
rect 6536 -9786 6576 -9752
rect 6610 -9786 6650 -9752
rect 6684 -9786 6724 -9752
rect 6758 -9786 6798 -9752
rect 6832 -9786 6872 -9752
rect 6906 -9786 6946 -9752
rect 6980 -9786 7020 -9752
rect 7054 -9786 7094 -9752
rect 7128 -9786 7168 -9752
rect 7202 -9786 7242 -9752
rect 7276 -9786 7316 -9752
rect 7350 -9786 7390 -9752
rect 7424 -9786 7464 -9752
rect 7498 -9786 7538 -9752
rect 7572 -9786 7612 -9752
rect 7646 -9786 7686 -9752
rect 7720 -9786 7760 -9752
rect 7794 -9786 7834 -9752
rect 7868 -9786 7908 -9752
rect 7942 -9786 7982 -9752
rect 8016 -9786 8056 -9752
rect 8090 -9786 8130 -9752
rect 8164 -9786 8204 -9752
rect 8238 -9786 8278 -9752
rect 8312 -9786 8352 -9752
rect 8386 -9786 8426 -9752
rect 8460 -9786 8500 -9752
rect 8534 -9786 8574 -9752
rect 8608 -9786 8648 -9752
rect 8682 -9786 8722 -9752
rect 8756 -9786 8796 -9752
rect 8830 -9786 8870 -9752
rect 8904 -9786 8944 -9752
rect 8978 -9786 9018 -9752
rect 9052 -9786 9092 -9752
rect 9126 -9786 9166 -9752
rect 9200 -9786 9240 -9752
rect 9274 -9786 9314 -9752
rect 9348 -9786 9388 -9752
rect 9422 -9786 9462 -9752
rect 9496 -9786 9536 -9752
rect 9570 -9786 9610 -9752
rect 9644 -9786 9684 -9752
rect 9718 -9786 9758 -9752
rect 9792 -9786 9832 -9752
rect 9866 -9786 9906 -9752
rect 9940 -9786 9980 -9752
rect 10014 -9786 10054 -9752
rect 10088 -9786 10128 -9752
rect 10162 -9786 10202 -9752
rect 10236 -9786 10276 -9752
rect 10310 -9786 10350 -9752
rect 10384 -9786 10424 -9752
rect 10458 -9786 10498 -9752
rect 10532 -9786 10572 -9752
rect 10606 -9786 10646 -9752
rect 10680 -9786 10720 -9752
rect 10754 -9786 10794 -9752
rect 10828 -9786 10868 -9752
rect 10902 -9786 10942 -9752
rect 10976 -9786 11016 -9752
rect 11050 -9786 11090 -9752
rect 11124 -9786 11164 -9752
rect 11198 -9786 11238 -9752
rect 11272 -9786 11312 -9752
rect 11346 -9786 11386 -9752
rect 11420 -9786 11460 -9752
rect 11494 -9786 11534 -9752
rect 11568 -9786 11608 -9752
rect 11642 -9786 11682 -9752
rect 11716 -9786 11756 -9752
rect 11790 -9786 11830 -9752
rect 11864 -9786 11904 -9752
rect 11938 -9786 11978 -9752
rect 12012 -9786 12052 -9752
rect 12086 -9786 12126 -9752
rect 12160 -9786 12200 -9752
rect 12234 -9786 12274 -9752
rect 12308 -9786 12348 -9752
rect 12382 -9786 12422 -9752
rect 12456 -9786 12496 -9752
rect 12530 -9786 12570 -9752
rect 12604 -9786 12644 -9752
rect 12678 -9786 12718 -9752
rect 12752 -9786 12792 -9752
rect 12826 -9786 12866 -9752
rect 12900 -9786 12940 -9752
rect 12974 -9786 13014 -9752
rect 13048 -9786 13088 -9752
rect 13122 -9786 13162 -9752
rect 13196 -9786 13236 -9752
rect 13270 -9786 13310 -9752
rect 13344 -9786 13384 -9752
rect 13418 -9786 13458 -9752
rect 13492 -9786 13532 -9752
rect 13566 -9786 13606 -9752
rect 13640 -9786 13680 -9752
rect 13714 -9786 13754 -9752
rect 13788 -9786 13828 -9752
rect 13862 -9786 13902 -9752
rect 13936 -9786 13976 -9752
rect 14010 -9786 14050 -9752
rect 14084 -9786 14124 -9752
rect 14158 -9786 14198 -9752
rect 14232 -9786 14272 -9752
rect 14306 -9786 14346 -9752
rect 14380 -9786 14420 -9752
rect 14454 -9786 14494 -9752
rect 14528 -9786 14568 -9752
rect 14602 -9786 14642 -9752
rect 14676 -9786 14716 -9752
rect 14750 -9786 14790 -9752
rect 14824 -9786 14864 -9752
rect 14898 -9786 14938 -9752
rect 14972 -9786 15012 -9752
rect 15046 -9786 15086 -9752
rect 15120 -9786 15160 -9752
rect 15194 -9786 15234 -9752
rect 15268 -9786 15308 -9752
rect 15342 -9786 15382 -9752
rect 15416 -9786 15456 -9752
rect 15490 -9786 15530 -9752
rect 15564 -9786 15604 -9752
rect 15638 -9786 15678 -9752
rect 15712 -9786 15752 -9752
rect 15786 -9786 15826 -9752
rect 15860 -9786 15900 -9752
rect 15934 -9786 15974 -9752
rect 16008 -9786 16048 -9752
rect 16082 -9786 16122 -9752
rect 16156 -9786 16196 -9752
rect 16230 -9786 16270 -9752
rect 16304 -9786 16344 -9752
rect 16378 -9786 16418 -9752
rect 16452 -9786 16492 -9752
rect 16526 -9786 16566 -9752
rect 16600 -9786 16640 -9752
rect 16674 -9786 16714 -9752
rect 16748 -9786 16788 -9752
rect 16822 -9786 16862 -9752
rect 16896 -9786 16936 -9752
rect 16970 -9786 17010 -9752
rect 17044 -9786 17084 -9752
rect 17118 -9786 17158 -9752
rect 17192 -9786 17232 -9752
rect 17266 -9786 17306 -9752
rect 17340 -9786 17380 -9752
rect 17414 -9786 17454 -9752
rect 17488 -9786 17528 -9752
rect 17562 -9786 17602 -9752
rect 17636 -9786 17676 -9752
rect 17710 -9786 17750 -9752
rect 17784 -9786 17824 -9752
rect 17858 -9786 17898 -9752
rect 17932 -9786 17972 -9752
rect 18006 -9786 18046 -9752
rect 18080 -9786 18120 -9752
rect 18154 -9786 18194 -9752
rect 18228 -9786 18268 -9752
rect 18302 -9786 18342 -9752
rect 18376 -9786 18416 -9752
rect 18450 -9786 18490 -9752
rect 18524 -9786 18564 -9752
rect 18598 -9786 18638 -9752
rect 18672 -9786 18712 -9752
rect 18746 -9786 18786 -9752
rect 18820 -9786 18860 -9752
rect 18894 -9786 18934 -9752
rect 18968 -9786 19008 -9752
rect 19042 -9786 19082 -9752
rect 19116 -9786 19156 -9752
rect 19190 -9786 19230 -9752
rect 19264 -9786 19304 -9752
rect 19338 -9786 19378 -9752
rect 19412 -9786 19452 -9752
rect 19486 -9786 19526 -9752
rect 19560 -9786 19600 -9752
rect 19634 -9786 19674 -9752
rect 19708 -9786 19748 -9752
rect 19782 -9786 19822 -9752
rect 19856 -9786 19896 -9752
rect 19930 -9786 19970 -9752
rect 20004 -9786 20044 -9752
rect 20078 -9786 20118 -9752
rect 20152 -9786 20192 -9752
rect 20226 -9786 20266 -9752
rect 20300 -9786 20340 -9752
rect 20374 -9786 20414 -9752
rect 20448 -9786 20488 -9752
rect 20522 -9786 20562 -9752
rect 20596 -9786 20636 -9752
rect 20670 -9786 20710 -9752
rect 20744 -9786 20784 -9752
rect 20818 -9786 20858 -9752
rect 20892 -9786 20932 -9752
rect 20966 -9786 21006 -9752
rect 21040 -9786 21080 -9752
rect 21114 -9786 21154 -9752
rect 21188 -9786 21228 -9752
rect 21262 -9786 21302 -9752
rect 21336 -9786 21376 -9752
rect 21410 -9786 21450 -9752
rect 21484 -9786 21524 -9752
rect 21558 -9786 21598 -9752
rect 21632 -9786 21672 -9752
rect 21706 -9786 21746 -9752
rect 21780 -9786 21820 -9752
rect 21854 -9786 21894 -9752
rect 21928 -9786 21968 -9752
rect 22002 -9786 22042 -9752
rect 22076 -9786 22116 -9752
rect 22150 -9786 22190 -9752
rect 22224 -9786 22264 -9752
rect 22298 -9786 22338 -9752
rect 22372 -9786 22412 -9752
rect 22446 -9786 22486 -9752
rect 22520 -9786 22560 -9752
rect 22594 -9786 22634 -9752
rect 22668 -9786 22708 -9752
rect 22742 -9786 22782 -9752
rect 22816 -9786 22856 -9752
rect 22890 -9786 22930 -9752
rect 22964 -9786 23004 -9752
rect 23038 -9786 23078 -9752
rect 23112 -9786 23152 -9752
rect 23186 -9786 23226 -9752
rect 23260 -9786 23300 -9752
rect 23334 -9786 23374 -9752
rect 23408 -9786 23448 -9752
rect 23482 -9786 23522 -9752
rect 23556 -9786 23596 -9752
rect 23630 -9786 23670 -9752
rect 23704 -9786 23744 -9752
rect 23778 -9786 23818 -9752
rect 23852 -9786 23892 -9752
rect 23926 -9786 23966 -9752
rect 24000 -9786 24040 -9752
rect 24074 -9786 24114 -9752
rect 24148 -9786 24188 -9752
rect 24222 -9786 24262 -9752
rect 24296 -9786 24336 -9752
rect 24370 -9786 24410 -9752
rect 24444 -9786 24484 -9752
rect 24518 -9786 24558 -9752
rect 24592 -9786 24632 -9752
rect 24666 -9786 24706 -9752
rect 24740 -9786 24780 -9752
rect 24814 -9786 24854 -9752
rect 24888 -9786 24928 -9752
rect 24962 -9786 25002 -9752
rect 25036 -9786 25076 -9752
rect 25110 -9786 25150 -9752
rect 25184 -9786 26250 -9752
rect 4020 -9860 4060 -9826
rect 4094 -9860 4134 -9826
rect 4168 -9860 4208 -9826
rect 4242 -9860 4282 -9826
rect 4316 -9860 4356 -9826
rect 4390 -9860 4430 -9826
rect 4464 -9860 4504 -9826
rect 4538 -9860 4578 -9826
rect 4612 -9860 4652 -9826
rect 4686 -9860 4726 -9826
rect 4760 -9860 4800 -9826
rect 4834 -9860 4874 -9826
rect 4908 -9860 4948 -9826
rect 4982 -9860 5022 -9826
rect 5056 -9860 5096 -9826
rect 5130 -9860 5170 -9826
rect 5204 -9860 5244 -9826
rect 5278 -9860 5318 -9826
rect 5352 -9860 5392 -9826
rect 5426 -9860 5466 -9826
rect 5500 -9860 5540 -9826
rect 5574 -9860 5614 -9826
rect 5648 -9860 5688 -9826
rect 5722 -9860 5762 -9826
rect 5796 -9860 5836 -9826
rect 5870 -9860 5910 -9826
rect 5944 -9860 5984 -9826
rect 6018 -9860 6058 -9826
rect 6092 -9860 6132 -9826
rect 6166 -9860 6206 -9826
rect 6240 -9860 6280 -9826
rect 6314 -9860 6354 -9826
rect 6388 -9860 6428 -9826
rect 6462 -9860 6502 -9826
rect 6536 -9860 6576 -9826
rect 6610 -9860 6650 -9826
rect 6684 -9860 6724 -9826
rect 6758 -9860 6798 -9826
rect 6832 -9860 6872 -9826
rect 6906 -9860 6946 -9826
rect 6980 -9860 7020 -9826
rect 7054 -9860 7094 -9826
rect 7128 -9860 7168 -9826
rect 7202 -9860 7242 -9826
rect 7276 -9860 7316 -9826
rect 7350 -9860 7390 -9826
rect 7424 -9860 7464 -9826
rect 7498 -9860 7538 -9826
rect 7572 -9860 7612 -9826
rect 7646 -9860 7686 -9826
rect 7720 -9860 7760 -9826
rect 7794 -9860 7834 -9826
rect 7868 -9860 7908 -9826
rect 7942 -9860 7982 -9826
rect 8016 -9860 8056 -9826
rect 8090 -9860 8130 -9826
rect 8164 -9860 8204 -9826
rect 8238 -9860 8278 -9826
rect 8312 -9860 8352 -9826
rect 8386 -9860 8426 -9826
rect 8460 -9860 8500 -9826
rect 8534 -9860 8574 -9826
rect 8608 -9860 8648 -9826
rect 8682 -9860 8722 -9826
rect 8756 -9860 8796 -9826
rect 8830 -9860 8870 -9826
rect 8904 -9860 8944 -9826
rect 8978 -9860 9018 -9826
rect 9052 -9860 9092 -9826
rect 9126 -9860 9166 -9826
rect 9200 -9860 9240 -9826
rect 9274 -9860 9314 -9826
rect 9348 -9860 9388 -9826
rect 9422 -9860 9462 -9826
rect 9496 -9860 9536 -9826
rect 9570 -9860 9610 -9826
rect 9644 -9860 9684 -9826
rect 9718 -9860 9758 -9826
rect 9792 -9860 9832 -9826
rect 9866 -9860 9906 -9826
rect 9940 -9860 9980 -9826
rect 10014 -9860 10054 -9826
rect 10088 -9860 10128 -9826
rect 10162 -9860 10202 -9826
rect 10236 -9860 10276 -9826
rect 10310 -9860 10350 -9826
rect 10384 -9860 10424 -9826
rect 10458 -9860 10498 -9826
rect 10532 -9860 10572 -9826
rect 10606 -9860 10646 -9826
rect 10680 -9860 10720 -9826
rect 10754 -9860 10794 -9826
rect 10828 -9860 10868 -9826
rect 10902 -9860 10942 -9826
rect 10976 -9860 11016 -9826
rect 11050 -9860 11090 -9826
rect 11124 -9860 11164 -9826
rect 11198 -9860 11238 -9826
rect 11272 -9860 11312 -9826
rect 11346 -9860 11386 -9826
rect 11420 -9860 11460 -9826
rect 11494 -9860 11534 -9826
rect 11568 -9860 11608 -9826
rect 11642 -9860 11682 -9826
rect 11716 -9860 11756 -9826
rect 11790 -9860 11830 -9826
rect 11864 -9860 11904 -9826
rect 11938 -9860 11978 -9826
rect 12012 -9860 12052 -9826
rect 12086 -9860 12126 -9826
rect 12160 -9860 12200 -9826
rect 12234 -9860 12274 -9826
rect 12308 -9860 12348 -9826
rect 12382 -9860 12422 -9826
rect 12456 -9860 12496 -9826
rect 12530 -9860 12570 -9826
rect 12604 -9860 12644 -9826
rect 12678 -9860 12718 -9826
rect 12752 -9860 12792 -9826
rect 12826 -9860 12866 -9826
rect 12900 -9860 12940 -9826
rect 12974 -9860 13014 -9826
rect 13048 -9860 13088 -9826
rect 13122 -9860 13162 -9826
rect 13196 -9860 13236 -9826
rect 13270 -9860 13310 -9826
rect 13344 -9860 13384 -9826
rect 13418 -9860 13458 -9826
rect 13492 -9860 13532 -9826
rect 13566 -9860 13606 -9826
rect 13640 -9860 13680 -9826
rect 13714 -9860 13754 -9826
rect 13788 -9860 13828 -9826
rect 13862 -9860 13902 -9826
rect 13936 -9860 13976 -9826
rect 14010 -9860 14050 -9826
rect 14084 -9860 14124 -9826
rect 14158 -9860 14198 -9826
rect 14232 -9860 14272 -9826
rect 14306 -9860 14346 -9826
rect 14380 -9860 14420 -9826
rect 14454 -9860 14494 -9826
rect 14528 -9860 14568 -9826
rect 14602 -9860 14642 -9826
rect 14676 -9860 14716 -9826
rect 14750 -9860 14790 -9826
rect 14824 -9860 14864 -9826
rect 14898 -9860 14938 -9826
rect 14972 -9860 15012 -9826
rect 15046 -9860 15086 -9826
rect 15120 -9860 15160 -9826
rect 15194 -9860 15234 -9826
rect 15268 -9860 15308 -9826
rect 15342 -9860 15382 -9826
rect 15416 -9860 15456 -9826
rect 15490 -9860 15530 -9826
rect 15564 -9860 15604 -9826
rect 15638 -9860 15678 -9826
rect 15712 -9860 15752 -9826
rect 15786 -9860 15826 -9826
rect 15860 -9860 15900 -9826
rect 15934 -9860 15974 -9826
rect 16008 -9860 16048 -9826
rect 16082 -9860 16122 -9826
rect 16156 -9860 16196 -9826
rect 16230 -9860 16270 -9826
rect 16304 -9860 16344 -9826
rect 16378 -9860 16418 -9826
rect 16452 -9860 16492 -9826
rect 16526 -9860 16566 -9826
rect 16600 -9860 16640 -9826
rect 16674 -9860 16714 -9826
rect 16748 -9860 16788 -9826
rect 16822 -9860 16862 -9826
rect 16896 -9860 16936 -9826
rect 16970 -9860 17010 -9826
rect 17044 -9860 17084 -9826
rect 17118 -9860 17158 -9826
rect 17192 -9860 17232 -9826
rect 17266 -9860 17306 -9826
rect 17340 -9860 17380 -9826
rect 17414 -9860 17454 -9826
rect 17488 -9860 17528 -9826
rect 17562 -9860 17602 -9826
rect 17636 -9860 17676 -9826
rect 17710 -9860 17750 -9826
rect 17784 -9860 17824 -9826
rect 17858 -9860 17898 -9826
rect 17932 -9860 17972 -9826
rect 18006 -9860 18046 -9826
rect 18080 -9860 18120 -9826
rect 18154 -9860 18194 -9826
rect 18228 -9860 18268 -9826
rect 18302 -9860 18342 -9826
rect 18376 -9860 18416 -9826
rect 18450 -9860 18490 -9826
rect 18524 -9860 18564 -9826
rect 18598 -9860 18638 -9826
rect 18672 -9860 18712 -9826
rect 18746 -9860 18786 -9826
rect 18820 -9860 18860 -9826
rect 18894 -9860 18934 -9826
rect 18968 -9860 19008 -9826
rect 19042 -9860 19082 -9826
rect 19116 -9860 19156 -9826
rect 19190 -9860 19230 -9826
rect 19264 -9860 19304 -9826
rect 19338 -9860 19378 -9826
rect 19412 -9860 19452 -9826
rect 19486 -9860 19526 -9826
rect 19560 -9860 19600 -9826
rect 19634 -9860 19674 -9826
rect 19708 -9860 19748 -9826
rect 19782 -9860 19822 -9826
rect 19856 -9860 19896 -9826
rect 19930 -9860 19970 -9826
rect 20004 -9860 20044 -9826
rect 20078 -9860 20118 -9826
rect 20152 -9860 20192 -9826
rect 20226 -9860 20266 -9826
rect 20300 -9860 20340 -9826
rect 20374 -9860 20414 -9826
rect 20448 -9860 20488 -9826
rect 20522 -9860 20562 -9826
rect 20596 -9860 20636 -9826
rect 20670 -9860 20710 -9826
rect 20744 -9860 20784 -9826
rect 20818 -9860 20858 -9826
rect 20892 -9860 20932 -9826
rect 20966 -9860 21006 -9826
rect 21040 -9860 21080 -9826
rect 21114 -9860 21154 -9826
rect 21188 -9860 21228 -9826
rect 21262 -9860 21302 -9826
rect 21336 -9860 21376 -9826
rect 21410 -9860 21450 -9826
rect 21484 -9860 21524 -9826
rect 21558 -9860 21598 -9826
rect 21632 -9860 21672 -9826
rect 21706 -9860 21746 -9826
rect 21780 -9860 21820 -9826
rect 21854 -9860 21894 -9826
rect 21928 -9860 21968 -9826
rect 22002 -9860 22042 -9826
rect 22076 -9860 22116 -9826
rect 22150 -9860 22190 -9826
rect 22224 -9860 22264 -9826
rect 22298 -9860 22338 -9826
rect 22372 -9860 22412 -9826
rect 22446 -9860 22486 -9826
rect 22520 -9860 22560 -9826
rect 22594 -9860 22634 -9826
rect 22668 -9860 22708 -9826
rect 22742 -9860 22782 -9826
rect 22816 -9860 22856 -9826
rect 22890 -9860 22930 -9826
rect 22964 -9860 23004 -9826
rect 23038 -9860 23078 -9826
rect 23112 -9860 23152 -9826
rect 23186 -9860 23226 -9826
rect 23260 -9860 23300 -9826
rect 23334 -9860 23374 -9826
rect 23408 -9860 23448 -9826
rect 23482 -9860 23522 -9826
rect 23556 -9860 23596 -9826
rect 23630 -9860 23670 -9826
rect 23704 -9860 23744 -9826
rect 23778 -9860 23818 -9826
rect 23852 -9860 23892 -9826
rect 23926 -9860 23966 -9826
rect 24000 -9860 24040 -9826
rect 24074 -9860 24114 -9826
rect 24148 -9860 24188 -9826
rect 24222 -9860 24262 -9826
rect 24296 -9860 24336 -9826
rect 24370 -9860 24410 -9826
rect 24444 -9860 24484 -9826
rect 24518 -9860 24558 -9826
rect 24592 -9860 24632 -9826
rect 24666 -9860 24706 -9826
rect 24740 -9860 24780 -9826
rect 24814 -9860 24854 -9826
rect 24888 -9860 24928 -9826
rect 24962 -9860 25002 -9826
rect 25036 -9860 25076 -9826
rect 25110 -9860 25150 -9826
rect 25184 -9860 26250 -9826
rect 4020 -9934 4060 -9900
rect 4094 -9934 4134 -9900
rect 4168 -9934 4208 -9900
rect 4242 -9934 4282 -9900
rect 4316 -9934 4356 -9900
rect 4390 -9934 4430 -9900
rect 4464 -9934 4504 -9900
rect 4538 -9934 4578 -9900
rect 4612 -9934 4652 -9900
rect 4686 -9934 4726 -9900
rect 4760 -9934 4800 -9900
rect 4834 -9934 4874 -9900
rect 4908 -9934 4948 -9900
rect 4982 -9934 5022 -9900
rect 5056 -9934 5096 -9900
rect 5130 -9934 5170 -9900
rect 5204 -9934 5244 -9900
rect 5278 -9934 5318 -9900
rect 5352 -9934 5392 -9900
rect 5426 -9934 5466 -9900
rect 5500 -9934 5540 -9900
rect 5574 -9934 5614 -9900
rect 5648 -9934 5688 -9900
rect 5722 -9934 5762 -9900
rect 5796 -9934 5836 -9900
rect 5870 -9934 5910 -9900
rect 5944 -9934 5984 -9900
rect 6018 -9934 6058 -9900
rect 6092 -9934 6132 -9900
rect 6166 -9934 6206 -9900
rect 6240 -9934 6280 -9900
rect 6314 -9934 6354 -9900
rect 6388 -9934 6428 -9900
rect 6462 -9934 6502 -9900
rect 6536 -9934 6576 -9900
rect 6610 -9934 6650 -9900
rect 6684 -9934 6724 -9900
rect 6758 -9934 6798 -9900
rect 6832 -9934 6872 -9900
rect 6906 -9934 6946 -9900
rect 6980 -9934 7020 -9900
rect 7054 -9934 7094 -9900
rect 7128 -9934 7168 -9900
rect 7202 -9934 7242 -9900
rect 7276 -9934 7316 -9900
rect 7350 -9934 7390 -9900
rect 7424 -9934 7464 -9900
rect 7498 -9934 7538 -9900
rect 7572 -9934 7612 -9900
rect 7646 -9934 7686 -9900
rect 7720 -9934 7760 -9900
rect 7794 -9934 7834 -9900
rect 7868 -9934 7908 -9900
rect 7942 -9934 7982 -9900
rect 8016 -9934 8056 -9900
rect 8090 -9934 8130 -9900
rect 8164 -9934 8204 -9900
rect 8238 -9934 8278 -9900
rect 8312 -9934 8352 -9900
rect 8386 -9934 8426 -9900
rect 8460 -9934 8500 -9900
rect 8534 -9934 8574 -9900
rect 8608 -9934 8648 -9900
rect 8682 -9934 8722 -9900
rect 8756 -9934 8796 -9900
rect 8830 -9934 8870 -9900
rect 8904 -9934 8944 -9900
rect 8978 -9934 9018 -9900
rect 9052 -9934 9092 -9900
rect 9126 -9934 9166 -9900
rect 9200 -9934 9240 -9900
rect 9274 -9934 9314 -9900
rect 9348 -9934 9388 -9900
rect 9422 -9934 9462 -9900
rect 9496 -9934 9536 -9900
rect 9570 -9934 9610 -9900
rect 9644 -9934 9684 -9900
rect 9718 -9934 9758 -9900
rect 9792 -9934 9832 -9900
rect 9866 -9934 9906 -9900
rect 9940 -9934 9980 -9900
rect 10014 -9934 10054 -9900
rect 10088 -9934 10128 -9900
rect 10162 -9934 10202 -9900
rect 10236 -9934 10276 -9900
rect 10310 -9934 10350 -9900
rect 10384 -9934 10424 -9900
rect 10458 -9934 10498 -9900
rect 10532 -9934 10572 -9900
rect 10606 -9934 10646 -9900
rect 10680 -9934 10720 -9900
rect 10754 -9934 10794 -9900
rect 10828 -9934 10868 -9900
rect 10902 -9934 10942 -9900
rect 10976 -9934 11016 -9900
rect 11050 -9934 11090 -9900
rect 11124 -9934 11164 -9900
rect 11198 -9934 11238 -9900
rect 11272 -9934 11312 -9900
rect 11346 -9934 11386 -9900
rect 11420 -9934 11460 -9900
rect 11494 -9934 11534 -9900
rect 11568 -9934 11608 -9900
rect 11642 -9934 11682 -9900
rect 11716 -9934 11756 -9900
rect 11790 -9934 11830 -9900
rect 11864 -9934 11904 -9900
rect 11938 -9934 11978 -9900
rect 12012 -9934 12052 -9900
rect 12086 -9934 12126 -9900
rect 12160 -9934 12200 -9900
rect 12234 -9934 12274 -9900
rect 12308 -9934 12348 -9900
rect 12382 -9934 12422 -9900
rect 12456 -9934 12496 -9900
rect 12530 -9934 12570 -9900
rect 12604 -9934 12644 -9900
rect 12678 -9934 12718 -9900
rect 12752 -9934 12792 -9900
rect 12826 -9934 12866 -9900
rect 12900 -9934 12940 -9900
rect 12974 -9934 13014 -9900
rect 13048 -9934 13088 -9900
rect 13122 -9934 13162 -9900
rect 13196 -9934 13236 -9900
rect 13270 -9934 13310 -9900
rect 13344 -9934 13384 -9900
rect 13418 -9934 13458 -9900
rect 13492 -9934 13532 -9900
rect 13566 -9934 13606 -9900
rect 13640 -9934 13680 -9900
rect 13714 -9934 13754 -9900
rect 13788 -9934 13828 -9900
rect 13862 -9934 13902 -9900
rect 13936 -9934 13976 -9900
rect 14010 -9934 14050 -9900
rect 14084 -9934 14124 -9900
rect 14158 -9934 14198 -9900
rect 14232 -9934 14272 -9900
rect 14306 -9934 14346 -9900
rect 14380 -9934 14420 -9900
rect 14454 -9934 14494 -9900
rect 14528 -9934 14568 -9900
rect 14602 -9934 14642 -9900
rect 14676 -9934 14716 -9900
rect 14750 -9934 14790 -9900
rect 14824 -9934 14864 -9900
rect 14898 -9934 14938 -9900
rect 14972 -9934 15012 -9900
rect 15046 -9934 15086 -9900
rect 15120 -9934 15160 -9900
rect 15194 -9934 15234 -9900
rect 15268 -9934 15308 -9900
rect 15342 -9934 15382 -9900
rect 15416 -9934 15456 -9900
rect 15490 -9934 15530 -9900
rect 15564 -9934 15604 -9900
rect 15638 -9934 15678 -9900
rect 15712 -9934 15752 -9900
rect 15786 -9934 15826 -9900
rect 15860 -9934 15900 -9900
rect 15934 -9934 15974 -9900
rect 16008 -9934 16048 -9900
rect 16082 -9934 16122 -9900
rect 16156 -9934 16196 -9900
rect 16230 -9934 16270 -9900
rect 16304 -9934 16344 -9900
rect 16378 -9934 16418 -9900
rect 16452 -9934 16492 -9900
rect 16526 -9934 16566 -9900
rect 16600 -9934 16640 -9900
rect 16674 -9934 16714 -9900
rect 16748 -9934 16788 -9900
rect 16822 -9934 16862 -9900
rect 16896 -9934 16936 -9900
rect 16970 -9934 17010 -9900
rect 17044 -9934 17084 -9900
rect 17118 -9934 17158 -9900
rect 17192 -9934 17232 -9900
rect 17266 -9934 17306 -9900
rect 17340 -9934 17380 -9900
rect 17414 -9934 17454 -9900
rect 17488 -9934 17528 -9900
rect 17562 -9934 17602 -9900
rect 17636 -9934 17676 -9900
rect 17710 -9934 17750 -9900
rect 17784 -9934 17824 -9900
rect 17858 -9934 17898 -9900
rect 17932 -9934 17972 -9900
rect 18006 -9934 18046 -9900
rect 18080 -9934 18120 -9900
rect 18154 -9934 18194 -9900
rect 18228 -9934 18268 -9900
rect 18302 -9934 18342 -9900
rect 18376 -9934 18416 -9900
rect 18450 -9934 18490 -9900
rect 18524 -9934 18564 -9900
rect 18598 -9934 18638 -9900
rect 18672 -9934 18712 -9900
rect 18746 -9934 18786 -9900
rect 18820 -9934 18860 -9900
rect 18894 -9934 18934 -9900
rect 18968 -9934 19008 -9900
rect 19042 -9934 19082 -9900
rect 19116 -9934 19156 -9900
rect 19190 -9934 19230 -9900
rect 19264 -9934 19304 -9900
rect 19338 -9934 19378 -9900
rect 19412 -9934 19452 -9900
rect 19486 -9934 19526 -9900
rect 19560 -9934 19600 -9900
rect 19634 -9934 19674 -9900
rect 19708 -9934 19748 -9900
rect 19782 -9934 19822 -9900
rect 19856 -9934 19896 -9900
rect 19930 -9934 19970 -9900
rect 20004 -9934 20044 -9900
rect 20078 -9934 20118 -9900
rect 20152 -9934 20192 -9900
rect 20226 -9934 20266 -9900
rect 20300 -9934 20340 -9900
rect 20374 -9934 20414 -9900
rect 20448 -9934 20488 -9900
rect 20522 -9934 20562 -9900
rect 20596 -9934 20636 -9900
rect 20670 -9934 20710 -9900
rect 20744 -9934 20784 -9900
rect 20818 -9934 20858 -9900
rect 20892 -9934 20932 -9900
rect 20966 -9934 21006 -9900
rect 21040 -9934 21080 -9900
rect 21114 -9934 21154 -9900
rect 21188 -9934 21228 -9900
rect 21262 -9934 21302 -9900
rect 21336 -9934 21376 -9900
rect 21410 -9934 21450 -9900
rect 21484 -9934 21524 -9900
rect 21558 -9934 21598 -9900
rect 21632 -9934 21672 -9900
rect 21706 -9934 21746 -9900
rect 21780 -9934 21820 -9900
rect 21854 -9934 21894 -9900
rect 21928 -9934 21968 -9900
rect 22002 -9934 22042 -9900
rect 22076 -9934 22116 -9900
rect 22150 -9934 22190 -9900
rect 22224 -9934 22264 -9900
rect 22298 -9934 22338 -9900
rect 22372 -9934 22412 -9900
rect 22446 -9934 22486 -9900
rect 22520 -9934 22560 -9900
rect 22594 -9934 22634 -9900
rect 22668 -9934 22708 -9900
rect 22742 -9934 22782 -9900
rect 22816 -9934 22856 -9900
rect 22890 -9934 22930 -9900
rect 22964 -9934 23004 -9900
rect 23038 -9934 23078 -9900
rect 23112 -9934 23152 -9900
rect 23186 -9934 23226 -9900
rect 23260 -9934 23300 -9900
rect 23334 -9934 23374 -9900
rect 23408 -9934 23448 -9900
rect 23482 -9934 23522 -9900
rect 23556 -9934 23596 -9900
rect 23630 -9934 23670 -9900
rect 23704 -9934 23744 -9900
rect 23778 -9934 23818 -9900
rect 23852 -9934 23892 -9900
rect 23926 -9934 23966 -9900
rect 24000 -9934 24040 -9900
rect 24074 -9934 24114 -9900
rect 24148 -9934 24188 -9900
rect 24222 -9934 24262 -9900
rect 24296 -9934 24336 -9900
rect 24370 -9934 24410 -9900
rect 24444 -9934 24484 -9900
rect 24518 -9934 24558 -9900
rect 24592 -9934 24632 -9900
rect 24666 -9934 24706 -9900
rect 24740 -9934 24780 -9900
rect 24814 -9934 24854 -9900
rect 24888 -9934 24928 -9900
rect 24962 -9934 25002 -9900
rect 25036 -9934 25076 -9900
rect 25110 -9934 25150 -9900
rect 25184 -9934 26250 -9900
<< viali >>
rect 4768 3118 4792 3152
rect 4792 3118 4802 3152
rect 4840 3118 4874 3152
rect 4912 3118 4946 3152
rect 4984 3118 5018 3152
rect 5056 3118 5090 3152
rect 5128 3118 5162 3152
rect 5200 3118 5234 3152
rect 5272 3118 5306 3152
rect 5344 3118 5378 3152
rect 5416 3118 5450 3152
rect 5488 3118 5522 3152
rect 5560 3118 5594 3152
rect 5632 3118 5666 3152
rect 5704 3118 5738 3152
rect 5776 3118 5810 3152
rect 5848 3118 5882 3152
rect 5920 3118 5954 3152
rect 5992 3118 6026 3152
rect 6064 3118 6098 3152
rect 6136 3118 6170 3152
rect 6208 3118 6242 3152
rect 6280 3118 6314 3152
rect 6352 3118 6386 3152
rect 6424 3118 6458 3152
rect 6496 3118 6530 3152
rect 6568 3118 6602 3152
rect 6640 3118 6674 3152
rect 6712 3118 6746 3152
rect 6784 3118 6818 3152
rect 6856 3118 6890 3152
rect 6928 3118 6962 3152
rect 7000 3118 7034 3152
rect 7072 3118 7106 3152
rect 7144 3118 7178 3152
rect 7216 3118 7250 3152
rect 7288 3118 7322 3152
rect 7360 3118 7394 3152
rect 7432 3118 7466 3152
rect 7504 3118 7538 3152
rect 7576 3118 7610 3152
rect 7648 3118 7682 3152
rect 7720 3118 7754 3152
rect 7792 3118 7826 3152
rect 7864 3118 7898 3152
rect 7936 3118 7970 3152
rect 8008 3118 8042 3152
rect 8080 3118 8114 3152
rect 8152 3118 8186 3152
rect 8224 3118 8258 3152
rect 8296 3118 8330 3152
rect 8368 3118 8402 3152
rect 8440 3118 8474 3152
rect 8512 3118 8546 3152
rect 8584 3118 8618 3152
rect 8656 3118 8690 3152
rect 8728 3118 8762 3152
rect 8800 3118 8834 3152
rect 8872 3118 8906 3152
rect 8944 3118 8978 3152
rect 9016 3118 9050 3152
rect 9088 3118 9122 3152
rect 9160 3118 9194 3152
rect 9232 3118 9266 3152
rect 9304 3118 9338 3152
rect 9376 3118 9410 3152
rect 9448 3118 9482 3152
rect 9520 3118 9554 3152
rect 9592 3118 9626 3152
rect 9664 3118 9698 3152
rect 9736 3118 9770 3152
rect 9808 3118 9842 3152
rect 9880 3118 9914 3152
rect 9952 3118 9986 3152
rect 10024 3118 10058 3152
rect 10096 3118 10130 3152
rect 10168 3118 10202 3152
rect 10240 3118 10274 3152
rect 10312 3118 10346 3152
rect 10384 3118 10418 3152
rect 10456 3118 10490 3152
rect 10528 3118 10562 3152
rect 10600 3118 10634 3152
rect 10672 3118 10706 3152
rect 10744 3118 10762 3152
rect 10762 3118 10778 3152
rect 12458 3117 12482 3151
rect 12482 3117 12492 3151
rect 12530 3117 12564 3151
rect 12602 3117 12636 3151
rect 12674 3117 12708 3151
rect 12746 3117 12780 3151
rect 12818 3117 12852 3151
rect 12890 3117 12924 3151
rect 12962 3117 12996 3151
rect 13034 3117 13068 3151
rect 13106 3117 13140 3151
rect 13178 3117 13212 3151
rect 13250 3117 13284 3151
rect 13322 3117 13356 3151
rect 13394 3117 13428 3151
rect 13466 3117 13500 3151
rect 13538 3117 13572 3151
rect 13610 3117 13644 3151
rect 13682 3117 13716 3151
rect 13754 3117 13788 3151
rect 13826 3117 13860 3151
rect 13898 3117 13932 3151
rect 13970 3117 14004 3151
rect 14042 3117 14076 3151
rect 14114 3117 14148 3151
rect 14186 3117 14220 3151
rect 14258 3117 14292 3151
rect 14330 3117 14364 3151
rect 14402 3117 14436 3151
rect 14474 3117 14508 3151
rect 14546 3117 14580 3151
rect 14618 3117 14652 3151
rect 14690 3117 14724 3151
rect 14762 3117 14796 3151
rect 14834 3117 14868 3151
rect 14906 3117 14940 3151
rect 14978 3117 15012 3151
rect 15050 3117 15084 3151
rect 15122 3117 15156 3151
rect 15194 3117 15228 3151
rect 15266 3117 15300 3151
rect 15338 3117 15372 3151
rect 15410 3117 15444 3151
rect 15482 3117 15516 3151
rect 15554 3117 15588 3151
rect 15626 3117 15660 3151
rect 15698 3117 15732 3151
rect 15770 3117 15804 3151
rect 15842 3117 15876 3151
rect 15914 3117 15948 3151
rect 15986 3117 16020 3151
rect 16058 3117 16092 3151
rect 16130 3117 16164 3151
rect 16202 3117 16236 3151
rect 16274 3117 16308 3151
rect 16346 3117 16380 3151
rect 16418 3117 16452 3151
rect 16490 3117 16524 3151
rect 16562 3117 16596 3151
rect 16634 3117 16668 3151
rect 16706 3117 16740 3151
rect 16778 3117 16812 3151
rect 16850 3117 16884 3151
rect 16922 3117 16956 3151
rect 16994 3117 17028 3151
rect 17066 3117 17100 3151
rect 17138 3117 17172 3151
rect 17210 3117 17244 3151
rect 17282 3117 17316 3151
rect 17354 3117 17388 3151
rect 17426 3117 17460 3151
rect 17498 3117 17532 3151
rect 17570 3117 17604 3151
rect 17642 3117 17676 3151
rect 17714 3117 17748 3151
rect 17786 3117 17820 3151
rect 17858 3117 17892 3151
rect 17930 3117 17964 3151
rect 18002 3117 18036 3151
rect 18074 3117 18108 3151
rect 18146 3117 18180 3151
rect 18218 3117 18252 3151
rect 18290 3117 18324 3151
rect 18362 3117 18396 3151
rect 18434 3117 18452 3151
rect 18452 3117 18468 3151
rect 18597 3117 18621 3151
rect 18621 3117 18631 3151
rect 18669 3117 18703 3151
rect 18741 3117 18775 3151
rect 18813 3117 18847 3151
rect 18885 3117 18919 3151
rect 18957 3117 18991 3151
rect 19029 3117 19063 3151
rect 19101 3117 19135 3151
rect 19173 3117 19207 3151
rect 19245 3117 19279 3151
rect 19317 3117 19351 3151
rect 19389 3117 19423 3151
rect 19461 3117 19495 3151
rect 19533 3117 19567 3151
rect 19605 3117 19639 3151
rect 19677 3117 19711 3151
rect 19749 3117 19783 3151
rect 19821 3117 19855 3151
rect 19893 3117 19927 3151
rect 19965 3117 19999 3151
rect 20037 3117 20071 3151
rect 20109 3117 20143 3151
rect 20181 3117 20215 3151
rect 20253 3117 20287 3151
rect 20325 3117 20359 3151
rect 20397 3117 20431 3151
rect 20469 3117 20503 3151
rect 20541 3117 20575 3151
rect 20613 3117 20647 3151
rect 20685 3117 20719 3151
rect 20757 3117 20791 3151
rect 20829 3117 20863 3151
rect 20901 3117 20935 3151
rect 20973 3117 21007 3151
rect 21045 3117 21079 3151
rect 21117 3117 21151 3151
rect 21189 3117 21223 3151
rect 21261 3117 21295 3151
rect 21333 3117 21367 3151
rect 21405 3117 21439 3151
rect 21477 3117 21511 3151
rect 21549 3117 21583 3151
rect 21621 3117 21655 3151
rect 21693 3117 21727 3151
rect 21765 3117 21799 3151
rect 21837 3117 21871 3151
rect 21909 3117 21943 3151
rect 21981 3117 22015 3151
rect 22053 3117 22087 3151
rect 22125 3117 22159 3151
rect 22197 3117 22231 3151
rect 22269 3117 22303 3151
rect 22341 3117 22375 3151
rect 22413 3117 22447 3151
rect 22485 3117 22519 3151
rect 22557 3117 22591 3151
rect 22629 3117 22663 3151
rect 22701 3117 22735 3151
rect 22773 3117 22807 3151
rect 22845 3117 22879 3151
rect 22917 3117 22951 3151
rect 22989 3117 23023 3151
rect 23061 3117 23095 3151
rect 23133 3117 23167 3151
rect 23205 3117 23239 3151
rect 23277 3117 23311 3151
rect 23349 3117 23383 3151
rect 23421 3117 23455 3151
rect 23493 3117 23527 3151
rect 23565 3117 23599 3151
rect 23637 3117 23671 3151
rect 23709 3117 23743 3151
rect 23781 3117 23815 3151
rect 23853 3117 23887 3151
rect 23925 3117 23959 3151
rect 23997 3117 24031 3151
rect 24069 3117 24103 3151
rect 24141 3117 24175 3151
rect 24213 3117 24247 3151
rect 24285 3117 24319 3151
rect 24357 3117 24391 3151
rect 24429 3117 24463 3151
rect 24501 3117 24535 3151
rect 24573 3117 24591 3151
rect 24591 3117 24607 3151
rect 4768 3030 4792 3064
rect 4792 3030 4802 3064
rect 4840 3030 4874 3064
rect 4912 3030 4946 3064
rect 4984 3030 5018 3064
rect 5056 3030 5090 3064
rect 5128 3030 5162 3064
rect 5200 3030 5234 3064
rect 5272 3030 5306 3064
rect 5344 3030 5378 3064
rect 5416 3030 5450 3064
rect 5488 3030 5522 3064
rect 5560 3030 5594 3064
rect 5632 3030 5666 3064
rect 5704 3030 5738 3064
rect 5776 3030 5810 3064
rect 5848 3030 5882 3064
rect 5920 3030 5954 3064
rect 5992 3030 6026 3064
rect 6064 3030 6098 3064
rect 6136 3030 6170 3064
rect 6208 3030 6242 3064
rect 6280 3030 6314 3064
rect 6352 3030 6386 3064
rect 6424 3030 6458 3064
rect 6496 3030 6530 3064
rect 6568 3030 6602 3064
rect 6640 3030 6674 3064
rect 6712 3030 6746 3064
rect 6784 3030 6818 3064
rect 6856 3030 6890 3064
rect 6928 3030 6962 3064
rect 7000 3030 7034 3064
rect 7072 3030 7106 3064
rect 7144 3030 7178 3064
rect 7216 3030 7250 3064
rect 7288 3030 7322 3064
rect 7360 3030 7394 3064
rect 7432 3030 7466 3064
rect 7504 3030 7538 3064
rect 7576 3030 7610 3064
rect 7648 3030 7682 3064
rect 7720 3030 7754 3064
rect 7792 3030 7826 3064
rect 7864 3030 7898 3064
rect 7936 3030 7970 3064
rect 8008 3030 8042 3064
rect 8080 3030 8114 3064
rect 8152 3030 8186 3064
rect 8224 3030 8258 3064
rect 8296 3030 8330 3064
rect 8368 3030 8402 3064
rect 8440 3030 8474 3064
rect 8512 3030 8546 3064
rect 8584 3030 8618 3064
rect 8656 3030 8690 3064
rect 8728 3030 8762 3064
rect 8800 3030 8834 3064
rect 8872 3030 8906 3064
rect 8944 3030 8978 3064
rect 9016 3030 9050 3064
rect 9088 3030 9122 3064
rect 9160 3030 9194 3064
rect 9232 3030 9266 3064
rect 9304 3030 9338 3064
rect 9376 3030 9410 3064
rect 9448 3030 9482 3064
rect 9520 3030 9554 3064
rect 9592 3030 9626 3064
rect 9664 3030 9698 3064
rect 9736 3030 9770 3064
rect 9808 3030 9842 3064
rect 9880 3030 9914 3064
rect 9952 3030 9986 3064
rect 10024 3030 10058 3064
rect 10096 3030 10130 3064
rect 10168 3030 10202 3064
rect 10240 3030 10274 3064
rect 10312 3030 10346 3064
rect 10384 3030 10418 3064
rect 10456 3030 10490 3064
rect 10528 3030 10562 3064
rect 10600 3030 10634 3064
rect 10672 3030 10706 3064
rect 10744 3030 10762 3064
rect 10762 3030 10778 3064
rect 12458 3029 12482 3063
rect 12482 3029 12492 3063
rect 12530 3029 12564 3063
rect 12602 3029 12636 3063
rect 12674 3029 12708 3063
rect 12746 3029 12780 3063
rect 12818 3029 12852 3063
rect 12890 3029 12924 3063
rect 12962 3029 12996 3063
rect 13034 3029 13068 3063
rect 13106 3029 13140 3063
rect 13178 3029 13212 3063
rect 13250 3029 13284 3063
rect 13322 3029 13356 3063
rect 13394 3029 13428 3063
rect 13466 3029 13500 3063
rect 13538 3029 13572 3063
rect 13610 3029 13644 3063
rect 13682 3029 13716 3063
rect 13754 3029 13788 3063
rect 13826 3029 13860 3063
rect 13898 3029 13932 3063
rect 13970 3029 14004 3063
rect 14042 3029 14076 3063
rect 14114 3029 14148 3063
rect 14186 3029 14220 3063
rect 14258 3029 14292 3063
rect 14330 3029 14364 3063
rect 14402 3029 14436 3063
rect 14474 3029 14508 3063
rect 14546 3029 14580 3063
rect 14618 3029 14652 3063
rect 14690 3029 14724 3063
rect 14762 3029 14796 3063
rect 14834 3029 14868 3063
rect 14906 3029 14940 3063
rect 14978 3029 15012 3063
rect 15050 3029 15084 3063
rect 15122 3029 15156 3063
rect 15194 3029 15228 3063
rect 15266 3029 15300 3063
rect 15338 3029 15372 3063
rect 15410 3029 15444 3063
rect 15482 3029 15516 3063
rect 15554 3029 15588 3063
rect 15626 3029 15660 3063
rect 15698 3029 15732 3063
rect 15770 3029 15804 3063
rect 15842 3029 15876 3063
rect 15914 3029 15948 3063
rect 15986 3029 16020 3063
rect 16058 3029 16092 3063
rect 16130 3029 16164 3063
rect 16202 3029 16236 3063
rect 16274 3029 16308 3063
rect 16346 3029 16380 3063
rect 16418 3029 16452 3063
rect 16490 3029 16524 3063
rect 16562 3029 16596 3063
rect 16634 3029 16668 3063
rect 16706 3029 16740 3063
rect 16778 3029 16812 3063
rect 16850 3029 16884 3063
rect 16922 3029 16956 3063
rect 16994 3029 17028 3063
rect 17066 3029 17100 3063
rect 17138 3029 17172 3063
rect 17210 3029 17244 3063
rect 17282 3029 17316 3063
rect 17354 3029 17388 3063
rect 17426 3029 17460 3063
rect 17498 3029 17532 3063
rect 17570 3029 17604 3063
rect 17642 3029 17676 3063
rect 17714 3029 17748 3063
rect 17786 3029 17820 3063
rect 17858 3029 17892 3063
rect 17930 3029 17964 3063
rect 18002 3029 18036 3063
rect 18074 3029 18108 3063
rect 18146 3029 18180 3063
rect 18218 3029 18252 3063
rect 18290 3029 18324 3063
rect 18362 3029 18396 3063
rect 18434 3029 18452 3063
rect 18452 3029 18468 3063
rect 18597 3029 18621 3063
rect 18621 3029 18631 3063
rect 18669 3029 18703 3063
rect 18741 3029 18775 3063
rect 18813 3029 18847 3063
rect 18885 3029 18919 3063
rect 18957 3029 18991 3063
rect 19029 3029 19063 3063
rect 19101 3029 19135 3063
rect 19173 3029 19207 3063
rect 19245 3029 19279 3063
rect 19317 3029 19351 3063
rect 19389 3029 19423 3063
rect 19461 3029 19495 3063
rect 19533 3029 19567 3063
rect 19605 3029 19639 3063
rect 19677 3029 19711 3063
rect 19749 3029 19783 3063
rect 19821 3029 19855 3063
rect 19893 3029 19927 3063
rect 19965 3029 19999 3063
rect 20037 3029 20071 3063
rect 20109 3029 20143 3063
rect 20181 3029 20215 3063
rect 20253 3029 20287 3063
rect 20325 3029 20359 3063
rect 20397 3029 20431 3063
rect 20469 3029 20503 3063
rect 20541 3029 20575 3063
rect 20613 3029 20647 3063
rect 20685 3029 20719 3063
rect 20757 3029 20791 3063
rect 20829 3029 20863 3063
rect 20901 3029 20935 3063
rect 20973 3029 21007 3063
rect 21045 3029 21079 3063
rect 21117 3029 21151 3063
rect 21189 3029 21223 3063
rect 21261 3029 21295 3063
rect 21333 3029 21367 3063
rect 21405 3029 21439 3063
rect 21477 3029 21511 3063
rect 21549 3029 21583 3063
rect 21621 3029 21655 3063
rect 21693 3029 21727 3063
rect 21765 3029 21799 3063
rect 21837 3029 21871 3063
rect 21909 3029 21943 3063
rect 21981 3029 22015 3063
rect 22053 3029 22087 3063
rect 22125 3029 22159 3063
rect 22197 3029 22231 3063
rect 22269 3029 22303 3063
rect 22341 3029 22375 3063
rect 22413 3029 22447 3063
rect 22485 3029 22519 3063
rect 22557 3029 22591 3063
rect 22629 3029 22663 3063
rect 22701 3029 22735 3063
rect 22773 3029 22807 3063
rect 22845 3029 22879 3063
rect 22917 3029 22951 3063
rect 22989 3029 23023 3063
rect 23061 3029 23095 3063
rect 23133 3029 23167 3063
rect 23205 3029 23239 3063
rect 23277 3029 23311 3063
rect 23349 3029 23383 3063
rect 23421 3029 23455 3063
rect 23493 3029 23527 3063
rect 23565 3029 23599 3063
rect 23637 3029 23671 3063
rect 23709 3029 23743 3063
rect 23781 3029 23815 3063
rect 23853 3029 23887 3063
rect 23925 3029 23959 3063
rect 23997 3029 24031 3063
rect 24069 3029 24103 3063
rect 24141 3029 24175 3063
rect 24213 3029 24247 3063
rect 24285 3029 24319 3063
rect 24357 3029 24391 3063
rect 24429 3029 24463 3063
rect 24501 3029 24535 3063
rect 24573 3029 24591 3063
rect 24591 3029 24607 3063
rect 4768 2942 4792 2976
rect 4792 2942 4802 2976
rect 4840 2942 4874 2976
rect 4912 2942 4946 2976
rect 4984 2942 5018 2976
rect 5056 2942 5090 2976
rect 5128 2942 5162 2976
rect 5200 2942 5234 2976
rect 5272 2942 5306 2976
rect 5344 2942 5378 2976
rect 5416 2942 5450 2976
rect 5488 2942 5522 2976
rect 5560 2942 5594 2976
rect 5632 2942 5666 2976
rect 5704 2942 5738 2976
rect 5776 2942 5810 2976
rect 5848 2942 5882 2976
rect 5920 2942 5954 2976
rect 5992 2942 6026 2976
rect 6064 2942 6098 2976
rect 6136 2942 6170 2976
rect 6208 2942 6242 2976
rect 6280 2942 6314 2976
rect 6352 2942 6386 2976
rect 6424 2942 6458 2976
rect 6496 2942 6530 2976
rect 6568 2942 6602 2976
rect 6640 2942 6674 2976
rect 6712 2942 6746 2976
rect 6784 2942 6818 2976
rect 6856 2942 6890 2976
rect 6928 2942 6962 2976
rect 7000 2942 7034 2976
rect 7072 2942 7106 2976
rect 7144 2942 7178 2976
rect 7216 2942 7250 2976
rect 7288 2942 7322 2976
rect 7360 2942 7394 2976
rect 7432 2942 7466 2976
rect 7504 2942 7538 2976
rect 7576 2942 7610 2976
rect 7648 2942 7682 2976
rect 7720 2942 7754 2976
rect 7792 2942 7826 2976
rect 7864 2942 7898 2976
rect 7936 2942 7970 2976
rect 8008 2942 8042 2976
rect 8080 2942 8114 2976
rect 8152 2942 8186 2976
rect 8224 2942 8258 2976
rect 8296 2942 8330 2976
rect 8368 2942 8402 2976
rect 8440 2942 8474 2976
rect 8512 2942 8546 2976
rect 8584 2942 8618 2976
rect 8656 2942 8690 2976
rect 8728 2942 8762 2976
rect 8800 2942 8834 2976
rect 8872 2942 8906 2976
rect 8944 2942 8978 2976
rect 9016 2942 9050 2976
rect 9088 2942 9122 2976
rect 9160 2942 9194 2976
rect 9232 2942 9266 2976
rect 9304 2942 9338 2976
rect 9376 2942 9410 2976
rect 9448 2942 9482 2976
rect 9520 2942 9554 2976
rect 9592 2942 9626 2976
rect 9664 2942 9698 2976
rect 9736 2942 9770 2976
rect 9808 2942 9842 2976
rect 9880 2942 9914 2976
rect 9952 2942 9986 2976
rect 10024 2942 10058 2976
rect 10096 2942 10130 2976
rect 10168 2942 10202 2976
rect 10240 2942 10274 2976
rect 10312 2942 10346 2976
rect 10384 2942 10418 2976
rect 10456 2942 10490 2976
rect 10528 2942 10562 2976
rect 10600 2942 10634 2976
rect 10672 2942 10706 2976
rect 10744 2942 10762 2976
rect 10762 2942 10778 2976
rect 12458 2941 12482 2975
rect 12482 2941 12492 2975
rect 12530 2941 12564 2975
rect 12602 2941 12636 2975
rect 12674 2941 12708 2975
rect 12746 2941 12780 2975
rect 12818 2941 12852 2975
rect 12890 2941 12924 2975
rect 12962 2941 12996 2975
rect 13034 2941 13068 2975
rect 13106 2941 13140 2975
rect 13178 2941 13212 2975
rect 13250 2941 13284 2975
rect 13322 2941 13356 2975
rect 13394 2941 13428 2975
rect 13466 2941 13500 2975
rect 13538 2941 13572 2975
rect 13610 2941 13644 2975
rect 13682 2941 13716 2975
rect 13754 2941 13788 2975
rect 13826 2941 13860 2975
rect 13898 2941 13932 2975
rect 13970 2941 14004 2975
rect 14042 2941 14076 2975
rect 14114 2941 14148 2975
rect 14186 2941 14220 2975
rect 14258 2941 14292 2975
rect 14330 2941 14364 2975
rect 14402 2941 14436 2975
rect 14474 2941 14508 2975
rect 14546 2941 14580 2975
rect 14618 2941 14652 2975
rect 14690 2941 14724 2975
rect 14762 2941 14796 2975
rect 14834 2941 14868 2975
rect 14906 2941 14940 2975
rect 14978 2941 15012 2975
rect 15050 2941 15084 2975
rect 15122 2941 15156 2975
rect 15194 2941 15228 2975
rect 15266 2941 15300 2975
rect 15338 2941 15372 2975
rect 15410 2941 15444 2975
rect 15482 2941 15516 2975
rect 15554 2941 15588 2975
rect 15626 2941 15660 2975
rect 15698 2941 15732 2975
rect 15770 2941 15804 2975
rect 15842 2941 15876 2975
rect 15914 2941 15948 2975
rect 15986 2941 16020 2975
rect 16058 2941 16092 2975
rect 16130 2941 16164 2975
rect 16202 2941 16236 2975
rect 16274 2941 16308 2975
rect 16346 2941 16380 2975
rect 16418 2941 16452 2975
rect 16490 2941 16524 2975
rect 16562 2941 16596 2975
rect 16634 2941 16668 2975
rect 16706 2941 16740 2975
rect 16778 2941 16812 2975
rect 16850 2941 16884 2975
rect 16922 2941 16956 2975
rect 16994 2941 17028 2975
rect 17066 2941 17100 2975
rect 17138 2941 17172 2975
rect 17210 2941 17244 2975
rect 17282 2941 17316 2975
rect 17354 2941 17388 2975
rect 17426 2941 17460 2975
rect 17498 2941 17532 2975
rect 17570 2941 17604 2975
rect 17642 2941 17676 2975
rect 17714 2941 17748 2975
rect 17786 2941 17820 2975
rect 17858 2941 17892 2975
rect 17930 2941 17964 2975
rect 18002 2941 18036 2975
rect 18074 2941 18108 2975
rect 18146 2941 18180 2975
rect 18218 2941 18252 2975
rect 18290 2941 18324 2975
rect 18362 2941 18396 2975
rect 18434 2941 18452 2975
rect 18452 2941 18468 2975
rect 18597 2941 18621 2975
rect 18621 2941 18631 2975
rect 18669 2941 18703 2975
rect 18741 2941 18775 2975
rect 18813 2941 18847 2975
rect 18885 2941 18919 2975
rect 18957 2941 18991 2975
rect 19029 2941 19063 2975
rect 19101 2941 19135 2975
rect 19173 2941 19207 2975
rect 19245 2941 19279 2975
rect 19317 2941 19351 2975
rect 19389 2941 19423 2975
rect 19461 2941 19495 2975
rect 19533 2941 19567 2975
rect 19605 2941 19639 2975
rect 19677 2941 19711 2975
rect 19749 2941 19783 2975
rect 19821 2941 19855 2975
rect 19893 2941 19927 2975
rect 19965 2941 19999 2975
rect 20037 2941 20071 2975
rect 20109 2941 20143 2975
rect 20181 2941 20215 2975
rect 20253 2941 20287 2975
rect 20325 2941 20359 2975
rect 20397 2941 20431 2975
rect 20469 2941 20503 2975
rect 20541 2941 20575 2975
rect 20613 2941 20647 2975
rect 20685 2941 20719 2975
rect 20757 2941 20791 2975
rect 20829 2941 20863 2975
rect 20901 2941 20935 2975
rect 20973 2941 21007 2975
rect 21045 2941 21079 2975
rect 21117 2941 21151 2975
rect 21189 2941 21223 2975
rect 21261 2941 21295 2975
rect 21333 2941 21367 2975
rect 21405 2941 21439 2975
rect 21477 2941 21511 2975
rect 21549 2941 21583 2975
rect 21621 2941 21655 2975
rect 21693 2941 21727 2975
rect 21765 2941 21799 2975
rect 21837 2941 21871 2975
rect 21909 2941 21943 2975
rect 21981 2941 22015 2975
rect 22053 2941 22087 2975
rect 22125 2941 22159 2975
rect 22197 2941 22231 2975
rect 22269 2941 22303 2975
rect 22341 2941 22375 2975
rect 22413 2941 22447 2975
rect 22485 2941 22519 2975
rect 22557 2941 22591 2975
rect 22629 2941 22663 2975
rect 22701 2941 22735 2975
rect 22773 2941 22807 2975
rect 22845 2941 22879 2975
rect 22917 2941 22951 2975
rect 22989 2941 23023 2975
rect 23061 2941 23095 2975
rect 23133 2941 23167 2975
rect 23205 2941 23239 2975
rect 23277 2941 23311 2975
rect 23349 2941 23383 2975
rect 23421 2941 23455 2975
rect 23493 2941 23527 2975
rect 23565 2941 23599 2975
rect 23637 2941 23671 2975
rect 23709 2941 23743 2975
rect 23781 2941 23815 2975
rect 23853 2941 23887 2975
rect 23925 2941 23959 2975
rect 23997 2941 24031 2975
rect 24069 2941 24103 2975
rect 24141 2941 24175 2975
rect 24213 2941 24247 2975
rect 24285 2941 24319 2975
rect 24357 2941 24391 2975
rect 24429 2941 24463 2975
rect 24501 2941 24535 2975
rect 24573 2941 24591 2975
rect 24591 2941 24607 2975
rect 18598 2835 18632 2869
rect 7398 2099 7432 2675
rect 12736 2098 12770 2674
rect 12854 2098 12888 2674
rect 12972 2098 13006 2674
rect 13090 2098 13124 2674
rect 13208 2098 13242 2674
rect 13326 2098 13360 2674
rect 13444 2098 13478 2674
rect 13562 2098 13596 2674
rect 13680 2098 13714 2674
rect 13798 2098 13832 2674
rect 13916 2098 13950 2674
rect 14034 2098 14068 2674
rect 14152 2098 14186 2674
rect 14270 2098 14304 2674
rect 14388 2098 14422 2674
rect 14506 2098 14540 2674
rect 14624 2098 14658 2674
rect 14742 2098 14776 2674
rect 14860 2098 14894 2674
rect 14978 2098 15012 2674
rect 15096 2098 15130 2674
rect 15214 2098 15248 2674
rect 15332 2098 15366 2674
rect 15450 2098 15484 2674
rect 15659 2653 15693 2687
rect 15731 2653 15765 2687
rect 15803 2653 15837 2687
rect 15875 2653 15909 2687
rect 15947 2653 15981 2687
rect 16019 2653 16053 2687
rect 16091 2653 16125 2687
rect 16163 2653 16197 2687
rect 16235 2653 16269 2687
rect 16307 2653 16341 2687
rect 16379 2653 16413 2687
rect 15659 2579 15693 2613
rect 15731 2579 15765 2613
rect 15803 2579 15837 2613
rect 15875 2579 15909 2613
rect 15947 2579 15981 2613
rect 16019 2579 16053 2613
rect 16091 2579 16125 2613
rect 16163 2579 16197 2613
rect 16235 2579 16269 2613
rect 16307 2579 16341 2613
rect 16379 2579 16413 2613
rect 15659 2505 15693 2539
rect 15731 2505 15765 2539
rect 15803 2505 15837 2539
rect 15875 2505 15909 2539
rect 15947 2505 15981 2539
rect 16019 2505 16053 2539
rect 16091 2505 16125 2539
rect 16163 2505 16197 2539
rect 16235 2505 16269 2539
rect 16307 2505 16341 2539
rect 16379 2505 16413 2539
rect 15659 2431 15693 2465
rect 15731 2431 15765 2465
rect 15803 2431 15837 2465
rect 15875 2431 15909 2465
rect 15947 2431 15981 2465
rect 16019 2431 16053 2465
rect 16091 2431 16125 2465
rect 16163 2431 16197 2465
rect 16235 2431 16269 2465
rect 16307 2431 16341 2465
rect 16379 2431 16413 2465
rect 15659 2357 15693 2391
rect 15731 2357 15765 2391
rect 15803 2357 15837 2391
rect 15875 2357 15909 2391
rect 15947 2357 15981 2391
rect 16019 2357 16053 2391
rect 16091 2357 16125 2391
rect 16163 2357 16197 2391
rect 16235 2357 16269 2391
rect 16307 2357 16341 2391
rect 16379 2357 16413 2391
rect 15659 2283 15693 2317
rect 15731 2283 15765 2317
rect 15803 2283 15837 2317
rect 15875 2283 15909 2317
rect 15947 2283 15981 2317
rect 16019 2283 16053 2317
rect 16091 2283 16125 2317
rect 16163 2283 16197 2317
rect 16235 2283 16269 2317
rect 16307 2283 16341 2317
rect 16379 2283 16413 2317
rect 15659 2209 15693 2243
rect 15731 2209 15765 2243
rect 15803 2209 15837 2243
rect 15875 2209 15909 2243
rect 15947 2209 15981 2243
rect 16019 2209 16053 2243
rect 16091 2209 16125 2243
rect 16163 2209 16197 2243
rect 16235 2209 16269 2243
rect 16307 2209 16341 2243
rect 16379 2209 16413 2243
rect 15659 2135 15693 2169
rect 15731 2135 15765 2169
rect 15803 2135 15837 2169
rect 15875 2135 15909 2169
rect 15947 2135 15981 2169
rect 16019 2135 16053 2169
rect 16091 2135 16125 2169
rect 16163 2135 16197 2169
rect 16235 2135 16269 2169
rect 16307 2135 16341 2169
rect 16379 2135 16413 2169
rect 16859 2098 16893 2674
rect 16977 2098 17011 2674
rect 17095 2098 17129 2674
rect 17213 2098 17247 2674
rect 17331 2098 17365 2674
rect 17449 2098 17483 2674
rect 17567 2098 17601 2674
rect 17685 2098 17719 2674
rect 17803 2098 17837 2674
rect 17921 2098 17955 2674
rect 18039 2098 18073 2674
rect 18157 2098 18191 2674
rect 18275 2098 18309 2674
rect 18393 2098 18427 2674
rect 18511 2098 18545 2674
rect 18629 2098 18663 2674
rect 18747 2098 18781 2674
rect 18865 2098 18899 2674
rect 18983 2098 19017 2674
rect 19101 2098 19135 2674
rect 19219 2098 19253 2674
rect 19337 2098 19371 2674
rect 19455 2098 19489 2674
rect 19573 2098 19607 2674
rect 19782 2653 19816 2687
rect 19854 2653 19888 2687
rect 19926 2653 19960 2687
rect 19998 2653 20032 2687
rect 20070 2653 20104 2687
rect 20142 2653 20176 2687
rect 20214 2653 20248 2687
rect 20286 2653 20320 2687
rect 20358 2653 20392 2687
rect 20430 2653 20464 2687
rect 20502 2653 20536 2687
rect 19782 2579 19816 2613
rect 19854 2579 19888 2613
rect 19926 2579 19960 2613
rect 19998 2579 20032 2613
rect 20070 2579 20104 2613
rect 20142 2579 20176 2613
rect 20214 2579 20248 2613
rect 20286 2579 20320 2613
rect 20358 2579 20392 2613
rect 20430 2579 20464 2613
rect 20502 2579 20536 2613
rect 19782 2505 19816 2539
rect 19854 2505 19888 2539
rect 19926 2505 19960 2539
rect 19998 2505 20032 2539
rect 20070 2505 20104 2539
rect 20142 2505 20176 2539
rect 20214 2505 20248 2539
rect 20286 2505 20320 2539
rect 20358 2505 20392 2539
rect 20430 2505 20464 2539
rect 20502 2505 20536 2539
rect 19782 2431 19816 2465
rect 19854 2431 19888 2465
rect 19926 2431 19960 2465
rect 19998 2431 20032 2465
rect 20070 2431 20104 2465
rect 20142 2431 20176 2465
rect 20214 2431 20248 2465
rect 20286 2431 20320 2465
rect 20358 2431 20392 2465
rect 20430 2431 20464 2465
rect 20502 2431 20536 2465
rect 19782 2357 19816 2391
rect 19854 2357 19888 2391
rect 19926 2357 19960 2391
rect 19998 2357 20032 2391
rect 20070 2357 20104 2391
rect 20142 2357 20176 2391
rect 20214 2357 20248 2391
rect 20286 2357 20320 2391
rect 20358 2357 20392 2391
rect 20430 2357 20464 2391
rect 20502 2357 20536 2391
rect 19782 2283 19816 2317
rect 19854 2283 19888 2317
rect 19926 2283 19960 2317
rect 19998 2283 20032 2317
rect 20070 2283 20104 2317
rect 20142 2283 20176 2317
rect 20214 2283 20248 2317
rect 20286 2283 20320 2317
rect 20358 2283 20392 2317
rect 20430 2283 20464 2317
rect 20502 2283 20536 2317
rect 19782 2209 19816 2243
rect 19854 2209 19888 2243
rect 19926 2209 19960 2243
rect 19998 2209 20032 2243
rect 20070 2209 20104 2243
rect 20142 2209 20176 2243
rect 20214 2209 20248 2243
rect 20286 2209 20320 2243
rect 20358 2209 20392 2243
rect 20430 2209 20464 2243
rect 20502 2209 20536 2243
rect 19782 2135 19816 2169
rect 19854 2135 19888 2169
rect 19926 2135 19960 2169
rect 19998 2135 20032 2169
rect 20070 2135 20104 2169
rect 20142 2135 20176 2169
rect 20214 2135 20248 2169
rect 20286 2135 20320 2169
rect 20358 2135 20392 2169
rect 20430 2135 20464 2169
rect 20502 2135 20536 2169
rect 20982 2098 21016 2674
rect 21100 2098 21134 2674
rect 21218 2098 21252 2674
rect 21336 2098 21370 2674
rect 21454 2098 21488 2674
rect 21572 2098 21606 2674
rect 21690 2098 21724 2674
rect 21808 2098 21842 2674
rect 21926 2098 21960 2674
rect 22044 2098 22078 2674
rect 22162 2098 22196 2674
rect 22280 2098 22314 2674
rect 22398 2098 22432 2674
rect 22516 2098 22550 2674
rect 22634 2098 22668 2674
rect 22752 2098 22786 2674
rect 22870 2098 22904 2674
rect 22988 2098 23022 2674
rect 23106 2098 23140 2674
rect 23224 2098 23258 2674
rect 23342 2098 23376 2674
rect 23460 2098 23494 2674
rect 23578 2098 23612 2674
rect 23696 2098 23730 2674
rect 23905 2653 23939 2687
rect 23977 2653 24011 2687
rect 24049 2653 24083 2687
rect 24121 2653 24155 2687
rect 24193 2653 24227 2687
rect 24265 2653 24299 2687
rect 24337 2653 24371 2687
rect 24409 2653 24443 2687
rect 24481 2653 24515 2687
rect 24553 2653 24587 2687
rect 24625 2653 24659 2687
rect 23905 2579 23939 2613
rect 23977 2579 24011 2613
rect 24049 2579 24083 2613
rect 24121 2579 24155 2613
rect 24193 2579 24227 2613
rect 24265 2579 24299 2613
rect 24337 2579 24371 2613
rect 24409 2579 24443 2613
rect 24481 2579 24515 2613
rect 24553 2579 24587 2613
rect 24625 2579 24659 2613
rect 23905 2505 23939 2539
rect 23977 2505 24011 2539
rect 24049 2505 24083 2539
rect 24121 2505 24155 2539
rect 24193 2505 24227 2539
rect 24265 2505 24299 2539
rect 24337 2505 24371 2539
rect 24409 2505 24443 2539
rect 24481 2505 24515 2539
rect 24553 2505 24587 2539
rect 24625 2505 24659 2539
rect 23905 2431 23939 2465
rect 23977 2431 24011 2465
rect 24049 2431 24083 2465
rect 24121 2431 24155 2465
rect 24193 2431 24227 2465
rect 24265 2431 24299 2465
rect 24337 2431 24371 2465
rect 24409 2431 24443 2465
rect 24481 2431 24515 2465
rect 24553 2431 24587 2465
rect 24625 2431 24659 2465
rect 23905 2357 23939 2391
rect 23977 2357 24011 2391
rect 24049 2357 24083 2391
rect 24121 2357 24155 2391
rect 24193 2357 24227 2391
rect 24265 2357 24299 2391
rect 24337 2357 24371 2391
rect 24409 2357 24443 2391
rect 24481 2357 24515 2391
rect 24553 2357 24587 2391
rect 24625 2357 24659 2391
rect 23905 2283 23939 2317
rect 23977 2283 24011 2317
rect 24049 2283 24083 2317
rect 24121 2283 24155 2317
rect 24193 2283 24227 2317
rect 24265 2283 24299 2317
rect 24337 2283 24371 2317
rect 24409 2283 24443 2317
rect 24481 2283 24515 2317
rect 24553 2283 24587 2317
rect 24625 2283 24659 2317
rect 23905 2209 23939 2243
rect 23977 2209 24011 2243
rect 24049 2209 24083 2243
rect 24121 2209 24155 2243
rect 24193 2209 24227 2243
rect 24265 2209 24299 2243
rect 24337 2209 24371 2243
rect 24409 2209 24443 2243
rect 24481 2209 24515 2243
rect 24553 2209 24587 2243
rect 24625 2209 24659 2243
rect 23905 2135 23939 2169
rect 23977 2135 24011 2169
rect 24049 2135 24083 2169
rect 24121 2135 24155 2169
rect 24193 2135 24227 2169
rect 24265 2135 24299 2169
rect 24337 2135 24371 2169
rect 24409 2135 24443 2169
rect 24481 2135 24515 2169
rect 24553 2135 24587 2169
rect 24625 2135 24659 2169
rect 15659 2061 15693 2095
rect 15731 2061 15765 2095
rect 15803 2061 15837 2095
rect 15875 2061 15909 2095
rect 15947 2061 15981 2095
rect 16019 2061 16053 2095
rect 16091 2061 16125 2095
rect 16163 2061 16197 2095
rect 16235 2061 16269 2095
rect 16307 2061 16341 2095
rect 16379 2061 16413 2095
rect 19782 2061 19816 2095
rect 19854 2061 19888 2095
rect 19926 2061 19960 2095
rect 19998 2061 20032 2095
rect 20070 2061 20104 2095
rect 20142 2061 20176 2095
rect 20214 2061 20248 2095
rect 20286 2061 20320 2095
rect 20358 2061 20392 2095
rect 20430 2061 20464 2095
rect 20502 2061 20536 2095
rect 23905 2061 23939 2095
rect 23977 2061 24011 2095
rect 24049 2061 24083 2095
rect 24121 2061 24155 2095
rect 24193 2061 24227 2095
rect 24265 2061 24299 2095
rect 24337 2061 24371 2095
rect 24409 2061 24443 2095
rect 24481 2061 24515 2095
rect 24553 2061 24587 2095
rect 24625 2061 24659 2095
rect 4869 2006 4903 2040
rect 4987 2006 5021 2040
rect 5105 2006 5139 2040
rect 5223 2006 5257 2040
rect 5341 2006 5375 2040
rect 5459 2006 5493 2040
rect 5577 2006 5611 2040
rect 5695 2006 5729 2040
rect 5813 2006 5847 2040
rect 5931 2006 5965 2040
rect 6049 2006 6083 2040
rect 6167 2006 6201 2040
rect 6285 2006 6319 2040
rect 6403 2006 6437 2040
rect 6521 2006 6555 2040
rect 7103 2006 7137 2040
rect 7221 2006 7255 2040
rect 7339 2006 7373 2040
rect 7457 2006 7491 2040
rect 7575 2006 7609 2040
rect 7693 2006 7727 2040
rect 7811 2006 7845 2040
rect 7929 2006 7963 2040
rect 8047 2006 8081 2040
rect 8165 2006 8199 2040
rect 8283 2006 8317 2040
rect 8401 2006 8435 2040
rect 8519 2006 8553 2040
rect 8865 2006 8899 2040
rect 8983 2006 9017 2040
rect 9101 2006 9135 2040
rect 9219 2006 9253 2040
rect 9337 2006 9371 2040
rect 9455 2006 9489 2040
rect 9573 2006 9607 2040
rect 9691 2006 9725 2040
rect 9809 2006 9843 2040
rect 9927 2006 9961 2040
rect 10045 2006 10079 2040
rect 10163 2006 10197 2040
rect 10281 2006 10315 2040
rect 10399 2006 10433 2040
rect 10517 2006 10551 2040
rect 12677 2005 12711 2039
rect 12795 2005 12829 2039
rect 12913 2005 12947 2039
rect 13031 2005 13065 2039
rect 13149 2005 13183 2039
rect 13267 2005 13301 2039
rect 13385 2005 13419 2039
rect 13503 2005 13537 2039
rect 13621 2005 13655 2039
rect 13739 2005 13773 2039
rect 13857 2005 13891 2039
rect 13975 2005 14009 2039
rect 14093 2005 14127 2039
rect 14211 2005 14245 2039
rect 14329 2005 14363 2039
rect 14447 2005 14481 2039
rect 14565 2005 14599 2039
rect 14683 2005 14717 2039
rect 14801 2005 14835 2039
rect 14919 2005 14953 2039
rect 15037 2005 15071 2039
rect 15155 2005 15189 2039
rect 15273 2005 15307 2039
rect 15391 2005 15425 2039
rect 15659 1987 15693 2021
rect 15731 1987 15765 2021
rect 15803 1987 15837 2021
rect 15875 1987 15909 2021
rect 15947 1987 15981 2021
rect 16019 1987 16053 2021
rect 16091 1987 16125 2021
rect 16163 1987 16197 2021
rect 16235 1987 16269 2021
rect 16307 1987 16341 2021
rect 16379 1987 16413 2021
rect 16800 2005 16834 2039
rect 16918 2005 16952 2039
rect 17036 2005 17070 2039
rect 17154 2005 17188 2039
rect 17272 2005 17306 2039
rect 17390 2005 17424 2039
rect 17508 2005 17542 2039
rect 17626 2005 17660 2039
rect 17744 2005 17778 2039
rect 17862 2005 17896 2039
rect 17980 2005 18014 2039
rect 18098 2005 18132 2039
rect 18216 2005 18250 2039
rect 18334 2005 18368 2039
rect 18452 2005 18486 2039
rect 18570 2005 18604 2039
rect 18688 2005 18722 2039
rect 18806 2005 18840 2039
rect 18924 2005 18958 2039
rect 19042 2005 19076 2039
rect 19160 2005 19194 2039
rect 19278 2005 19312 2039
rect 19396 2005 19430 2039
rect 19514 2005 19548 2039
rect 19782 1987 19816 2021
rect 19854 1987 19888 2021
rect 19926 1987 19960 2021
rect 19998 1987 20032 2021
rect 20070 1987 20104 2021
rect 20142 1987 20176 2021
rect 20214 1987 20248 2021
rect 20286 1987 20320 2021
rect 20358 1987 20392 2021
rect 20430 1987 20464 2021
rect 20502 1987 20536 2021
rect 20923 2005 20957 2039
rect 21041 2005 21075 2039
rect 21159 2005 21193 2039
rect 21277 2005 21311 2039
rect 21395 2005 21429 2039
rect 21513 2005 21547 2039
rect 21631 2005 21665 2039
rect 21749 2005 21783 2039
rect 21867 2005 21901 2039
rect 21985 2005 22019 2039
rect 22103 2005 22137 2039
rect 22221 2005 22255 2039
rect 22339 2005 22373 2039
rect 22457 2005 22491 2039
rect 22575 2005 22609 2039
rect 22693 2005 22727 2039
rect 22811 2005 22845 2039
rect 22929 2005 22963 2039
rect 23047 2005 23081 2039
rect 23165 2005 23199 2039
rect 23283 2005 23317 2039
rect 23401 2005 23435 2039
rect 23519 2005 23553 2039
rect 23637 2005 23671 2039
rect 23905 1987 23939 2021
rect 23977 1987 24011 2021
rect 24049 1987 24083 2021
rect 24121 1987 24155 2021
rect 24193 1987 24227 2021
rect 24265 1987 24299 2021
rect 24337 1987 24371 2021
rect 24409 1987 24443 2021
rect 24481 1987 24515 2021
rect 24553 1987 24587 2021
rect 24625 1987 24659 2021
rect 12677 1897 12711 1931
rect 12795 1897 12829 1931
rect 12913 1897 12947 1931
rect 13031 1897 13065 1931
rect 13149 1897 13183 1931
rect 13267 1897 13301 1931
rect 13385 1897 13419 1931
rect 13503 1897 13537 1931
rect 13621 1897 13655 1931
rect 13739 1897 13773 1931
rect 13857 1897 13891 1931
rect 13975 1897 14009 1931
rect 14093 1897 14127 1931
rect 14211 1897 14245 1931
rect 14329 1897 14363 1931
rect 14447 1897 14481 1931
rect 14565 1897 14599 1931
rect 14683 1897 14717 1931
rect 14801 1897 14835 1931
rect 14919 1897 14953 1931
rect 15037 1897 15071 1931
rect 15155 1897 15189 1931
rect 15273 1897 15307 1931
rect 15391 1897 15425 1931
rect 15659 1913 15693 1947
rect 15731 1913 15765 1947
rect 15803 1913 15837 1947
rect 15875 1913 15909 1947
rect 15947 1913 15981 1947
rect 16019 1913 16053 1947
rect 16091 1913 16125 1947
rect 16163 1913 16197 1947
rect 16235 1913 16269 1947
rect 16307 1913 16341 1947
rect 16379 1913 16413 1947
rect 16800 1897 16834 1931
rect 16918 1897 16952 1931
rect 17036 1897 17070 1931
rect 17154 1897 17188 1931
rect 17272 1897 17306 1931
rect 17390 1897 17424 1931
rect 17508 1897 17542 1931
rect 17626 1897 17660 1931
rect 17744 1897 17778 1931
rect 17862 1897 17896 1931
rect 17980 1897 18014 1931
rect 18098 1897 18132 1931
rect 18216 1897 18250 1931
rect 18334 1897 18368 1931
rect 18452 1897 18486 1931
rect 18570 1897 18604 1931
rect 18688 1897 18722 1931
rect 18806 1897 18840 1931
rect 18924 1897 18958 1931
rect 19042 1897 19076 1931
rect 19160 1897 19194 1931
rect 19278 1897 19312 1931
rect 19396 1897 19430 1931
rect 19514 1897 19548 1931
rect 19782 1913 19816 1947
rect 19854 1913 19888 1947
rect 19926 1913 19960 1947
rect 19998 1913 20032 1947
rect 20070 1913 20104 1947
rect 20142 1913 20176 1947
rect 20214 1913 20248 1947
rect 20286 1913 20320 1947
rect 20358 1913 20392 1947
rect 20430 1913 20464 1947
rect 20502 1913 20536 1947
rect 20923 1897 20957 1931
rect 21041 1897 21075 1931
rect 21159 1897 21193 1931
rect 21277 1897 21311 1931
rect 21395 1897 21429 1931
rect 21513 1897 21547 1931
rect 21631 1897 21665 1931
rect 21749 1897 21783 1931
rect 21867 1897 21901 1931
rect 21985 1897 22019 1931
rect 22103 1897 22137 1931
rect 22221 1897 22255 1931
rect 22339 1897 22373 1931
rect 22457 1897 22491 1931
rect 22575 1897 22609 1931
rect 22693 1897 22727 1931
rect 22811 1897 22845 1931
rect 22929 1897 22963 1931
rect 23047 1897 23081 1931
rect 23165 1897 23199 1931
rect 23283 1897 23317 1931
rect 23401 1897 23435 1931
rect 23519 1897 23553 1931
rect 23637 1897 23671 1931
rect 23905 1913 23939 1947
rect 23977 1913 24011 1947
rect 24049 1913 24083 1947
rect 24121 1913 24155 1947
rect 24193 1913 24227 1947
rect 24265 1913 24299 1947
rect 24337 1913 24371 1947
rect 24409 1913 24443 1947
rect 24481 1913 24515 1947
rect 24553 1913 24587 1947
rect 24625 1913 24659 1947
rect 15659 1839 15693 1873
rect 15731 1839 15765 1873
rect 15803 1839 15837 1873
rect 15875 1839 15909 1873
rect 15947 1839 15981 1873
rect 16019 1839 16053 1873
rect 16091 1839 16125 1873
rect 16163 1839 16197 1873
rect 16235 1839 16269 1873
rect 16307 1839 16341 1873
rect 16379 1839 16413 1873
rect 19782 1839 19816 1873
rect 19854 1839 19888 1873
rect 19926 1839 19960 1873
rect 19998 1839 20032 1873
rect 20070 1839 20104 1873
rect 20142 1839 20176 1873
rect 20214 1839 20248 1873
rect 20286 1839 20320 1873
rect 20358 1839 20392 1873
rect 20430 1839 20464 1873
rect 20502 1839 20536 1873
rect 23905 1839 23939 1873
rect 23977 1839 24011 1873
rect 24049 1839 24083 1873
rect 24121 1839 24155 1873
rect 24193 1839 24227 1873
rect 24265 1839 24299 1873
rect 24337 1839 24371 1873
rect 24409 1839 24443 1873
rect 24481 1839 24515 1873
rect 24553 1839 24587 1873
rect 24625 1839 24659 1873
rect 4810 602 4844 1178
rect 4928 602 4962 1178
rect 5046 602 5080 1178
rect 5164 602 5198 1178
rect 5282 602 5316 1178
rect 5400 602 5434 1178
rect 5518 602 5552 1178
rect 5636 602 5670 1178
rect 5754 602 5788 1178
rect 5872 602 5906 1178
rect 5990 602 6024 1178
rect 6108 602 6142 1178
rect 6226 602 6260 1178
rect 6344 602 6378 1178
rect 6462 602 6496 1178
rect 6580 602 6614 1178
rect 6698 602 6732 1178
rect 6816 602 6850 1178
rect 6934 602 6968 1178
rect 7052 602 7086 1178
rect 7170 602 7204 1178
rect 7288 602 7322 1178
rect 7406 602 7440 1178
rect 7524 602 7558 1178
rect 7642 602 7676 1178
rect 7760 602 7794 1178
rect 7878 602 7912 1178
rect 7996 602 8030 1178
rect 8114 602 8148 1178
rect 8232 602 8266 1178
rect 8350 602 8384 1178
rect 8468 602 8502 1178
rect 8586 602 8620 1178
rect 8704 602 8738 1178
rect 8822 602 8856 1178
rect 8940 602 8974 1178
rect 9058 602 9092 1178
rect 9176 602 9210 1178
rect 9294 602 9328 1178
rect 9412 602 9446 1178
rect 9530 602 9564 1178
rect 9648 602 9682 1178
rect 9766 602 9800 1178
rect 9884 602 9918 1178
rect 10002 602 10036 1178
rect 10120 602 10154 1178
rect 10238 602 10272 1178
rect 10356 602 10390 1178
rect 10474 602 10508 1178
rect 10592 602 10626 1178
rect 10710 602 10744 1178
rect 4869 509 4903 543
rect 4987 509 5021 543
rect 5105 509 5139 543
rect 5223 509 5257 543
rect 5341 509 5375 543
rect 5459 509 5493 543
rect 5577 509 5611 543
rect 5695 509 5729 543
rect 5813 509 5847 543
rect 5931 509 5965 543
rect 6049 509 6083 543
rect 6167 509 6201 543
rect 6285 509 6319 543
rect 6403 509 6437 543
rect 6521 509 6555 543
rect 6639 509 6673 543
rect 6757 509 6791 543
rect 6875 509 6909 543
rect 6993 509 7027 543
rect 7111 509 7145 543
rect 7229 509 7263 543
rect 7347 509 7381 543
rect 7465 509 7499 543
rect 7583 509 7617 543
rect 7701 509 7735 543
rect 7819 509 7853 543
rect 7937 509 7971 543
rect 8055 509 8089 543
rect 8173 509 8207 543
rect 8291 509 8325 543
rect 8409 509 8443 543
rect 8527 509 8561 543
rect 8645 509 8679 543
rect 8763 509 8797 543
rect 8881 509 8915 543
rect 8999 509 9033 543
rect 9117 509 9151 543
rect 9235 509 9269 543
rect 9353 509 9387 543
rect 9471 509 9505 543
rect 9589 509 9623 543
rect 9707 509 9741 543
rect 9825 509 9859 543
rect 9943 509 9977 543
rect 10061 509 10095 543
rect 10179 509 10213 543
rect 10297 509 10331 543
rect 10415 509 10449 543
rect 10533 509 10567 543
rect 10651 509 10685 543
rect 4869 401 4903 435
rect 4987 401 5021 435
rect 5105 401 5139 435
rect 5223 401 5257 435
rect 5341 401 5375 435
rect 5459 401 5493 435
rect 5577 401 5611 435
rect 5695 401 5729 435
rect 5813 401 5847 435
rect 5931 401 5965 435
rect 6049 401 6083 435
rect 6167 401 6201 435
rect 6285 401 6319 435
rect 6403 401 6437 435
rect 6521 401 6555 435
rect 6639 401 6673 435
rect 6757 401 6791 435
rect 6875 401 6909 435
rect 6993 401 7027 435
rect 7111 401 7145 435
rect 7229 401 7263 435
rect 7347 401 7381 435
rect 7465 401 7499 435
rect 7583 401 7617 435
rect 7701 401 7735 435
rect 7819 401 7853 435
rect 7937 401 7971 435
rect 8055 401 8089 435
rect 8173 401 8207 435
rect 8291 401 8325 435
rect 8409 401 8443 435
rect 8527 401 8561 435
rect 8645 401 8679 435
rect 8763 401 8797 435
rect 8881 401 8915 435
rect 8999 401 9033 435
rect 9117 401 9151 435
rect 9235 401 9269 435
rect 9353 401 9387 435
rect 9471 401 9505 435
rect 9589 401 9623 435
rect 9707 401 9741 435
rect 9825 401 9859 435
rect 9943 401 9977 435
rect 10061 401 10095 435
rect 10179 401 10213 435
rect 10297 401 10331 435
rect 10415 401 10449 435
rect 10533 401 10567 435
rect 10651 401 10685 435
rect 4810 -234 4844 342
rect 4928 -234 4962 342
rect 5046 -234 5080 342
rect 5164 -234 5198 342
rect 5282 -234 5316 342
rect 5400 -234 5434 342
rect 5518 -234 5552 342
rect 5636 -234 5670 342
rect 5754 -234 5788 342
rect 5872 -234 5906 342
rect 5990 -234 6024 342
rect 6108 -234 6142 342
rect 6226 -234 6260 342
rect 6344 -234 6378 342
rect 6462 -234 6496 342
rect 6580 -234 6614 342
rect 6698 -234 6732 342
rect 6816 -234 6850 342
rect 6934 -234 6968 342
rect 7052 -234 7086 342
rect 7170 -234 7204 342
rect 7288 -234 7322 342
rect 7406 -234 7440 342
rect 7524 -234 7558 342
rect 7642 -234 7676 342
rect 7760 -234 7794 342
rect 7878 -234 7912 342
rect 7996 -234 8030 342
rect 8114 -234 8148 342
rect 8232 -234 8266 342
rect 8350 -234 8384 342
rect 8468 -234 8502 342
rect 8586 -234 8620 342
rect 8704 -234 8738 342
rect 8822 -234 8856 342
rect 8940 -234 8974 342
rect 9058 -234 9092 342
rect 9176 -234 9210 342
rect 9294 -234 9328 342
rect 9412 -234 9446 342
rect 9530 -234 9564 342
rect 9648 -234 9682 342
rect 9766 -234 9800 342
rect 9884 -234 9918 342
rect 10002 -234 10036 342
rect 10120 -234 10154 342
rect 10238 -234 10272 342
rect 10356 -234 10390 342
rect 10474 -234 10508 342
rect 10592 -234 10626 342
rect 10710 -234 10744 342
rect 12500 1262 12534 1838
rect 12618 1262 12652 1838
rect 12736 1262 12770 1838
rect 12854 1262 12888 1838
rect 12972 1262 13006 1838
rect 13090 1262 13124 1838
rect 13208 1262 13242 1838
rect 13326 1262 13360 1838
rect 13444 1262 13478 1838
rect 13562 1262 13596 1838
rect 13680 1262 13714 1838
rect 13798 1262 13832 1838
rect 13916 1262 13950 1838
rect 14034 1262 14068 1838
rect 14152 1262 14186 1838
rect 14270 1262 14304 1838
rect 14388 1262 14422 1838
rect 14506 1262 14540 1838
rect 14624 1262 14658 1838
rect 14742 1262 14776 1838
rect 14860 1262 14894 1838
rect 14978 1262 15012 1838
rect 15096 1262 15130 1838
rect 15214 1262 15248 1838
rect 15332 1262 15366 1838
rect 15450 1262 15484 1838
rect 15659 1765 15693 1799
rect 15731 1765 15765 1799
rect 15803 1765 15837 1799
rect 15875 1765 15909 1799
rect 15947 1765 15981 1799
rect 16019 1765 16053 1799
rect 16091 1765 16125 1799
rect 16163 1765 16197 1799
rect 16235 1765 16269 1799
rect 16307 1765 16341 1799
rect 16379 1765 16413 1799
rect 15659 1691 15693 1725
rect 15731 1691 15765 1725
rect 15803 1691 15837 1725
rect 15875 1691 15909 1725
rect 15947 1691 15981 1725
rect 16019 1691 16053 1725
rect 16091 1691 16125 1725
rect 16163 1691 16197 1725
rect 16235 1691 16269 1725
rect 16307 1691 16341 1725
rect 16379 1691 16413 1725
rect 15659 1617 15693 1651
rect 15731 1617 15765 1651
rect 15803 1617 15837 1651
rect 15875 1617 15909 1651
rect 15947 1617 15981 1651
rect 16019 1617 16053 1651
rect 16091 1617 16125 1651
rect 16163 1617 16197 1651
rect 16235 1617 16269 1651
rect 16307 1617 16341 1651
rect 16379 1617 16413 1651
rect 15659 1543 15693 1577
rect 15731 1543 15765 1577
rect 15803 1543 15837 1577
rect 15875 1543 15909 1577
rect 15947 1543 15981 1577
rect 16019 1543 16053 1577
rect 16091 1543 16125 1577
rect 16163 1543 16197 1577
rect 16235 1543 16269 1577
rect 16307 1543 16341 1577
rect 16379 1543 16413 1577
rect 15659 1469 15693 1503
rect 15731 1469 15765 1503
rect 15803 1469 15837 1503
rect 15875 1469 15909 1503
rect 15947 1469 15981 1503
rect 16019 1469 16053 1503
rect 16091 1469 16125 1503
rect 16163 1469 16197 1503
rect 16235 1469 16269 1503
rect 16307 1469 16341 1503
rect 16379 1469 16413 1503
rect 15659 1395 15693 1429
rect 15731 1395 15765 1429
rect 15803 1395 15837 1429
rect 15875 1395 15909 1429
rect 15947 1395 15981 1429
rect 16019 1395 16053 1429
rect 16091 1395 16125 1429
rect 16163 1395 16197 1429
rect 16235 1395 16269 1429
rect 16307 1395 16341 1429
rect 16379 1395 16413 1429
rect 15659 1321 15693 1355
rect 15731 1321 15765 1355
rect 15803 1321 15837 1355
rect 15875 1321 15909 1355
rect 15947 1321 15981 1355
rect 16019 1321 16053 1355
rect 16091 1321 16125 1355
rect 16163 1321 16197 1355
rect 16235 1321 16269 1355
rect 16307 1321 16341 1355
rect 16379 1321 16413 1355
rect 15659 1247 15693 1281
rect 15731 1247 15765 1281
rect 15803 1247 15837 1281
rect 15875 1247 15909 1281
rect 15947 1247 15981 1281
rect 16019 1247 16053 1281
rect 16091 1247 16125 1281
rect 16163 1247 16197 1281
rect 16235 1247 16269 1281
rect 16307 1247 16341 1281
rect 16379 1247 16413 1281
rect 16623 1262 16657 1838
rect 16741 1262 16775 1838
rect 16859 1262 16893 1838
rect 16977 1262 17011 1838
rect 17095 1262 17129 1838
rect 17213 1262 17247 1838
rect 17331 1262 17365 1838
rect 17449 1262 17483 1838
rect 17567 1262 17601 1838
rect 17685 1262 17719 1838
rect 17803 1262 17837 1838
rect 17921 1262 17955 1838
rect 18039 1262 18073 1838
rect 18157 1262 18191 1838
rect 18275 1262 18309 1838
rect 18393 1262 18427 1838
rect 18511 1262 18545 1838
rect 18629 1262 18663 1838
rect 18747 1262 18781 1838
rect 18865 1262 18899 1838
rect 18983 1262 19017 1838
rect 19101 1262 19135 1838
rect 19219 1262 19253 1838
rect 19337 1262 19371 1838
rect 19455 1262 19489 1838
rect 19573 1262 19607 1838
rect 19782 1765 19816 1799
rect 19854 1765 19888 1799
rect 19926 1765 19960 1799
rect 19998 1765 20032 1799
rect 20070 1765 20104 1799
rect 20142 1765 20176 1799
rect 20214 1765 20248 1799
rect 20286 1765 20320 1799
rect 20358 1765 20392 1799
rect 20430 1765 20464 1799
rect 20502 1765 20536 1799
rect 19782 1691 19816 1725
rect 19854 1691 19888 1725
rect 19926 1691 19960 1725
rect 19998 1691 20032 1725
rect 20070 1691 20104 1725
rect 20142 1691 20176 1725
rect 20214 1691 20248 1725
rect 20286 1691 20320 1725
rect 20358 1691 20392 1725
rect 20430 1691 20464 1725
rect 20502 1691 20536 1725
rect 19782 1617 19816 1651
rect 19854 1617 19888 1651
rect 19926 1617 19960 1651
rect 19998 1617 20032 1651
rect 20070 1617 20104 1651
rect 20142 1617 20176 1651
rect 20214 1617 20248 1651
rect 20286 1617 20320 1651
rect 20358 1617 20392 1651
rect 20430 1617 20464 1651
rect 20502 1617 20536 1651
rect 19782 1543 19816 1577
rect 19854 1543 19888 1577
rect 19926 1543 19960 1577
rect 19998 1543 20032 1577
rect 20070 1543 20104 1577
rect 20142 1543 20176 1577
rect 20214 1543 20248 1577
rect 20286 1543 20320 1577
rect 20358 1543 20392 1577
rect 20430 1543 20464 1577
rect 20502 1543 20536 1577
rect 19782 1469 19816 1503
rect 19854 1469 19888 1503
rect 19926 1469 19960 1503
rect 19998 1469 20032 1503
rect 20070 1469 20104 1503
rect 20142 1469 20176 1503
rect 20214 1469 20248 1503
rect 20286 1469 20320 1503
rect 20358 1469 20392 1503
rect 20430 1469 20464 1503
rect 20502 1469 20536 1503
rect 19782 1395 19816 1429
rect 19854 1395 19888 1429
rect 19926 1395 19960 1429
rect 19998 1395 20032 1429
rect 20070 1395 20104 1429
rect 20142 1395 20176 1429
rect 20214 1395 20248 1429
rect 20286 1395 20320 1429
rect 20358 1395 20392 1429
rect 20430 1395 20464 1429
rect 20502 1395 20536 1429
rect 19782 1321 19816 1355
rect 19854 1321 19888 1355
rect 19926 1321 19960 1355
rect 19998 1321 20032 1355
rect 20070 1321 20104 1355
rect 20142 1321 20176 1355
rect 20214 1321 20248 1355
rect 20286 1321 20320 1355
rect 20358 1321 20392 1355
rect 20430 1321 20464 1355
rect 20502 1321 20536 1355
rect 19782 1247 19816 1281
rect 19854 1247 19888 1281
rect 19926 1247 19960 1281
rect 19998 1247 20032 1281
rect 20070 1247 20104 1281
rect 20142 1247 20176 1281
rect 20214 1247 20248 1281
rect 20286 1247 20320 1281
rect 20358 1247 20392 1281
rect 20430 1247 20464 1281
rect 20502 1247 20536 1281
rect 20746 1262 20780 1838
rect 20864 1262 20898 1838
rect 20982 1262 21016 1838
rect 21100 1262 21134 1838
rect 21218 1262 21252 1838
rect 21336 1262 21370 1838
rect 21454 1262 21488 1838
rect 21572 1262 21606 1838
rect 21690 1262 21724 1838
rect 21808 1262 21842 1838
rect 21926 1262 21960 1838
rect 22044 1262 22078 1838
rect 22162 1262 22196 1838
rect 22280 1262 22314 1838
rect 22398 1262 22432 1838
rect 22516 1262 22550 1838
rect 22634 1262 22668 1838
rect 22752 1262 22786 1838
rect 22870 1262 22904 1838
rect 22988 1262 23022 1838
rect 23106 1262 23140 1838
rect 23224 1262 23258 1838
rect 23342 1262 23376 1838
rect 23460 1262 23494 1838
rect 23578 1262 23612 1838
rect 23696 1262 23730 1838
rect 23905 1765 23939 1799
rect 23977 1765 24011 1799
rect 24049 1765 24083 1799
rect 24121 1765 24155 1799
rect 24193 1765 24227 1799
rect 24265 1765 24299 1799
rect 24337 1765 24371 1799
rect 24409 1765 24443 1799
rect 24481 1765 24515 1799
rect 24553 1765 24587 1799
rect 24625 1765 24659 1799
rect 23905 1691 23939 1725
rect 23977 1691 24011 1725
rect 24049 1691 24083 1725
rect 24121 1691 24155 1725
rect 24193 1691 24227 1725
rect 24265 1691 24299 1725
rect 24337 1691 24371 1725
rect 24409 1691 24443 1725
rect 24481 1691 24515 1725
rect 24553 1691 24587 1725
rect 24625 1691 24659 1725
rect 23905 1617 23939 1651
rect 23977 1617 24011 1651
rect 24049 1617 24083 1651
rect 24121 1617 24155 1651
rect 24193 1617 24227 1651
rect 24265 1617 24299 1651
rect 24337 1617 24371 1651
rect 24409 1617 24443 1651
rect 24481 1617 24515 1651
rect 24553 1617 24587 1651
rect 24625 1617 24659 1651
rect 23905 1543 23939 1577
rect 23977 1543 24011 1577
rect 24049 1543 24083 1577
rect 24121 1543 24155 1577
rect 24193 1543 24227 1577
rect 24265 1543 24299 1577
rect 24337 1543 24371 1577
rect 24409 1543 24443 1577
rect 24481 1543 24515 1577
rect 24553 1543 24587 1577
rect 24625 1543 24659 1577
rect 23905 1469 23939 1503
rect 23977 1469 24011 1503
rect 24049 1469 24083 1503
rect 24121 1469 24155 1503
rect 24193 1469 24227 1503
rect 24265 1469 24299 1503
rect 24337 1469 24371 1503
rect 24409 1469 24443 1503
rect 24481 1469 24515 1503
rect 24553 1469 24587 1503
rect 24625 1469 24659 1503
rect 23905 1395 23939 1429
rect 23977 1395 24011 1429
rect 24049 1395 24083 1429
rect 24121 1395 24155 1429
rect 24193 1395 24227 1429
rect 24265 1395 24299 1429
rect 24337 1395 24371 1429
rect 24409 1395 24443 1429
rect 24481 1395 24515 1429
rect 24553 1395 24587 1429
rect 24625 1395 24659 1429
rect 23905 1321 23939 1355
rect 23977 1321 24011 1355
rect 24049 1321 24083 1355
rect 24121 1321 24155 1355
rect 24193 1321 24227 1355
rect 24265 1321 24299 1355
rect 24337 1321 24371 1355
rect 24409 1321 24443 1355
rect 24481 1321 24515 1355
rect 24553 1321 24587 1355
rect 24625 1321 24659 1355
rect 23905 1247 23939 1281
rect 23977 1247 24011 1281
rect 24049 1247 24083 1281
rect 24121 1247 24155 1281
rect 24193 1247 24227 1281
rect 24265 1247 24299 1281
rect 24337 1247 24371 1281
rect 24409 1247 24443 1281
rect 24481 1247 24515 1281
rect 24553 1247 24587 1281
rect 24625 1247 24659 1281
rect 12479 1067 12513 1101
rect 4776 -429 4792 -395
rect 4792 -429 4810 -395
rect 4848 -429 4882 -395
rect 4920 -429 4954 -395
rect 4992 -429 5026 -395
rect 5064 -429 5098 -395
rect 5136 -429 5170 -395
rect 5208 -429 5242 -395
rect 5280 -429 5314 -395
rect 5352 -429 5386 -395
rect 5424 -429 5458 -395
rect 5496 -429 5530 -395
rect 5568 -429 5602 -395
rect 5640 -429 5674 -395
rect 5712 -429 5746 -395
rect 5784 -429 5818 -395
rect 5856 -429 5890 -395
rect 5928 -429 5962 -395
rect 6000 -429 6034 -395
rect 6072 -429 6106 -395
rect 6144 -429 6178 -395
rect 6216 -429 6250 -395
rect 6288 -429 6322 -395
rect 6360 -429 6394 -395
rect 6432 -429 6466 -395
rect 6504 -429 6538 -395
rect 6576 -429 6610 -395
rect 6648 -429 6682 -395
rect 6720 -429 6754 -395
rect 6792 -429 6826 -395
rect 6864 -429 6898 -395
rect 6936 -429 6970 -395
rect 7008 -429 7042 -395
rect 7080 -429 7114 -395
rect 7152 -429 7186 -395
rect 7224 -429 7258 -395
rect 7296 -429 7330 -395
rect 7368 -429 7402 -395
rect 7440 -429 7474 -395
rect 7512 -429 7546 -395
rect 7584 -429 7618 -395
rect 7656 -429 7690 -395
rect 7728 -429 7762 -395
rect 7800 -429 7834 -395
rect 7872 -429 7906 -395
rect 7944 -429 7978 -395
rect 8016 -429 8050 -395
rect 8088 -429 8122 -395
rect 8160 -429 8194 -395
rect 8232 -429 8266 -395
rect 8304 -429 8338 -395
rect 8376 -429 8410 -395
rect 8448 -429 8482 -395
rect 8520 -429 8554 -395
rect 8592 -429 8626 -395
rect 8664 -429 8698 -395
rect 8736 -429 8770 -395
rect 8808 -429 8842 -395
rect 8880 -429 8914 -395
rect 8952 -429 8986 -395
rect 9024 -429 9058 -395
rect 9096 -429 9130 -395
rect 9168 -429 9202 -395
rect 9240 -429 9274 -395
rect 9312 -429 9346 -395
rect 9384 -429 9418 -395
rect 9456 -429 9490 -395
rect 9528 -429 9562 -395
rect 9600 -429 9634 -395
rect 9672 -429 9706 -395
rect 9744 -429 9778 -395
rect 9816 -429 9850 -395
rect 9888 -429 9922 -395
rect 9960 -429 9994 -395
rect 10032 -429 10066 -395
rect 10104 -429 10138 -395
rect 10176 -429 10210 -395
rect 10248 -429 10282 -395
rect 10320 -429 10354 -395
rect 10392 -429 10426 -395
rect 10464 -429 10498 -395
rect 10536 -429 10570 -395
rect 10608 -429 10642 -395
rect 10680 -429 10714 -395
rect 10752 -429 10762 -395
rect 10762 -429 10786 -395
rect 4776 -517 4792 -483
rect 4792 -517 4810 -483
rect 4848 -517 4882 -483
rect 4920 -517 4954 -483
rect 4992 -517 5026 -483
rect 5064 -517 5098 -483
rect 5136 -517 5170 -483
rect 5208 -517 5242 -483
rect 5280 -517 5314 -483
rect 5352 -517 5386 -483
rect 5424 -517 5458 -483
rect 5496 -517 5530 -483
rect 5568 -517 5602 -483
rect 5640 -517 5674 -483
rect 5712 -517 5746 -483
rect 5784 -517 5818 -483
rect 5856 -517 5890 -483
rect 5928 -517 5962 -483
rect 6000 -517 6034 -483
rect 6072 -517 6106 -483
rect 6144 -517 6178 -483
rect 6216 -517 6250 -483
rect 6288 -517 6322 -483
rect 6360 -517 6394 -483
rect 6432 -517 6466 -483
rect 6504 -517 6538 -483
rect 6576 -517 6610 -483
rect 6648 -517 6682 -483
rect 6720 -517 6754 -483
rect 6792 -517 6826 -483
rect 6864 -517 6898 -483
rect 6936 -517 6970 -483
rect 7008 -517 7042 -483
rect 7080 -517 7114 -483
rect 7152 -517 7186 -483
rect 7224 -517 7258 -483
rect 7296 -517 7330 -483
rect 7368 -517 7402 -483
rect 7440 -517 7474 -483
rect 7512 -517 7546 -483
rect 7584 -517 7618 -483
rect 7656 -517 7690 -483
rect 7728 -517 7762 -483
rect 7800 -517 7834 -483
rect 7872 -517 7906 -483
rect 7944 -517 7978 -483
rect 8016 -517 8050 -483
rect 8088 -517 8122 -483
rect 8160 -517 8194 -483
rect 8232 -517 8266 -483
rect 8304 -517 8338 -483
rect 8376 -517 8410 -483
rect 8448 -517 8482 -483
rect 8520 -517 8554 -483
rect 8592 -517 8626 -483
rect 8664 -517 8698 -483
rect 8736 -517 8770 -483
rect 8808 -517 8842 -483
rect 8880 -517 8914 -483
rect 8952 -517 8986 -483
rect 9024 -517 9058 -483
rect 9096 -517 9130 -483
rect 9168 -517 9202 -483
rect 9240 -517 9274 -483
rect 9312 -517 9346 -483
rect 9384 -517 9418 -483
rect 9456 -517 9490 -483
rect 9528 -517 9562 -483
rect 9600 -517 9634 -483
rect 9672 -517 9706 -483
rect 9744 -517 9778 -483
rect 9816 -517 9850 -483
rect 9888 -517 9922 -483
rect 9960 -517 9994 -483
rect 10032 -517 10066 -483
rect 10104 -517 10138 -483
rect 10176 -517 10210 -483
rect 10248 -517 10282 -483
rect 10320 -517 10354 -483
rect 10392 -517 10426 -483
rect 10464 -517 10498 -483
rect 10536 -517 10570 -483
rect 10608 -517 10642 -483
rect 10680 -517 10714 -483
rect 10752 -517 10762 -483
rect 10762 -517 10786 -483
rect 4776 -605 4792 -571
rect 4792 -605 4810 -571
rect 4848 -605 4882 -571
rect 4920 -605 4954 -571
rect 4992 -605 5026 -571
rect 5064 -605 5098 -571
rect 5136 -605 5170 -571
rect 5208 -605 5242 -571
rect 5280 -605 5314 -571
rect 5352 -605 5386 -571
rect 5424 -605 5458 -571
rect 5496 -605 5530 -571
rect 5568 -605 5602 -571
rect 5640 -605 5674 -571
rect 5712 -605 5746 -571
rect 5784 -605 5818 -571
rect 5856 -605 5890 -571
rect 5928 -605 5962 -571
rect 6000 -605 6034 -571
rect 6072 -605 6106 -571
rect 6144 -605 6178 -571
rect 6216 -605 6250 -571
rect 6288 -605 6322 -571
rect 6360 -605 6394 -571
rect 6432 -605 6466 -571
rect 6504 -605 6538 -571
rect 6576 -605 6610 -571
rect 6648 -605 6682 -571
rect 6720 -605 6754 -571
rect 6792 -605 6826 -571
rect 6864 -605 6898 -571
rect 6936 -605 6970 -571
rect 7008 -605 7042 -571
rect 7080 -605 7114 -571
rect 7152 -605 7186 -571
rect 7224 -605 7258 -571
rect 7296 -605 7330 -571
rect 7368 -605 7402 -571
rect 7440 -605 7474 -571
rect 7512 -605 7546 -571
rect 7584 -605 7618 -571
rect 7656 -605 7690 -571
rect 7728 -605 7762 -571
rect 7800 -605 7834 -571
rect 7872 -605 7906 -571
rect 7944 -605 7978 -571
rect 8016 -605 8050 -571
rect 8088 -605 8122 -571
rect 8160 -605 8194 -571
rect 8232 -605 8266 -571
rect 8304 -605 8338 -571
rect 8376 -605 8410 -571
rect 8448 -605 8482 -571
rect 8520 -605 8554 -571
rect 8592 -605 8626 -571
rect 8664 -605 8698 -571
rect 8736 -605 8770 -571
rect 8808 -605 8842 -571
rect 8880 -605 8914 -571
rect 8952 -605 8986 -571
rect 9024 -605 9058 -571
rect 9096 -605 9130 -571
rect 9168 -605 9202 -571
rect 9240 -605 9274 -571
rect 9312 -605 9346 -571
rect 9384 -605 9418 -571
rect 9456 -605 9490 -571
rect 9528 -605 9562 -571
rect 9600 -605 9634 -571
rect 9672 -605 9706 -571
rect 9744 -605 9778 -571
rect 9816 -605 9850 -571
rect 9888 -605 9922 -571
rect 9960 -605 9994 -571
rect 10032 -605 10066 -571
rect 10104 -605 10138 -571
rect 10176 -605 10210 -571
rect 10248 -605 10282 -571
rect 10320 -605 10354 -571
rect 10392 -605 10426 -571
rect 10464 -605 10498 -571
rect 10536 -605 10570 -571
rect 10608 -605 10642 -571
rect 10680 -605 10714 -571
rect 10752 -605 10762 -571
rect 10762 -605 10786 -571
rect 4810 -1448 4844 -872
rect 4928 -1448 4962 -872
rect 5046 -1448 5080 -872
rect 5164 -1448 5198 -872
rect 5282 -1448 5316 -872
rect 5400 -1448 5434 -872
rect 5518 -1448 5552 -872
rect 5636 -1448 5670 -872
rect 5754 -1448 5788 -872
rect 5872 -1448 5906 -872
rect 5990 -1448 6024 -872
rect 6108 -1448 6142 -872
rect 6226 -1448 6260 -872
rect 6344 -1448 6378 -872
rect 6462 -1448 6496 -872
rect 6580 -1448 6614 -872
rect 6698 -1448 6732 -872
rect 6816 -1448 6850 -872
rect 6934 -1448 6968 -872
rect 7052 -1448 7086 -872
rect 7170 -1448 7204 -872
rect 7288 -1448 7322 -872
rect 7406 -1448 7440 -872
rect 7524 -1448 7558 -872
rect 7642 -1448 7676 -872
rect 7760 -1448 7794 -872
rect 7878 -1448 7912 -872
rect 7996 -1448 8030 -872
rect 8114 -1448 8148 -872
rect 8232 -1448 8266 -872
rect 8350 -1448 8384 -872
rect 8468 -1448 8502 -872
rect 8586 -1448 8620 -872
rect 8704 -1448 8738 -872
rect 8822 -1448 8856 -872
rect 8940 -1448 8974 -872
rect 9058 -1448 9092 -872
rect 9176 -1448 9210 -872
rect 9294 -1448 9328 -872
rect 9412 -1448 9446 -872
rect 9530 -1448 9564 -872
rect 9648 -1448 9682 -872
rect 9766 -1448 9800 -872
rect 9884 -1448 9918 -872
rect 10002 -1448 10036 -872
rect 10120 -1448 10154 -872
rect 10238 -1448 10272 -872
rect 10356 -1448 10390 -872
rect 10474 -1448 10508 -872
rect 10592 -1448 10626 -872
rect 10710 -1448 10744 -872
rect 4869 -1541 4903 -1507
rect 4987 -1541 5021 -1507
rect 5105 -1541 5139 -1507
rect 5223 -1541 5257 -1507
rect 5341 -1541 5375 -1507
rect 5459 -1541 5493 -1507
rect 5577 -1541 5611 -1507
rect 5695 -1541 5729 -1507
rect 5813 -1541 5847 -1507
rect 5931 -1541 5965 -1507
rect 6049 -1541 6083 -1507
rect 6167 -1541 6201 -1507
rect 6285 -1541 6319 -1507
rect 6403 -1541 6437 -1507
rect 6521 -1541 6555 -1507
rect 6639 -1541 6673 -1507
rect 6757 -1541 6791 -1507
rect 6875 -1541 6909 -1507
rect 6993 -1541 7027 -1507
rect 7111 -1541 7145 -1507
rect 7229 -1541 7263 -1507
rect 7347 -1541 7381 -1507
rect 7465 -1541 7499 -1507
rect 7583 -1541 7617 -1507
rect 7701 -1541 7735 -1507
rect 7819 -1541 7853 -1507
rect 7937 -1541 7971 -1507
rect 8055 -1541 8089 -1507
rect 8173 -1541 8207 -1507
rect 8291 -1541 8325 -1507
rect 8409 -1541 8443 -1507
rect 8527 -1541 8561 -1507
rect 8645 -1541 8679 -1507
rect 8763 -1541 8797 -1507
rect 8881 -1541 8915 -1507
rect 8999 -1541 9033 -1507
rect 9117 -1541 9151 -1507
rect 9235 -1541 9269 -1507
rect 9353 -1541 9387 -1507
rect 9471 -1541 9505 -1507
rect 9589 -1541 9623 -1507
rect 9707 -1541 9741 -1507
rect 9825 -1541 9859 -1507
rect 9943 -1541 9977 -1507
rect 10061 -1541 10095 -1507
rect 10179 -1541 10213 -1507
rect 10297 -1541 10331 -1507
rect 10415 -1541 10449 -1507
rect 10533 -1541 10567 -1507
rect 10651 -1541 10685 -1507
rect 4869 -1649 4903 -1615
rect 4987 -1649 5021 -1615
rect 5105 -1649 5139 -1615
rect 5223 -1649 5257 -1615
rect 5341 -1649 5375 -1615
rect 5459 -1649 5493 -1615
rect 5577 -1649 5611 -1615
rect 5695 -1649 5729 -1615
rect 5813 -1649 5847 -1615
rect 5931 -1649 5965 -1615
rect 6049 -1649 6083 -1615
rect 6167 -1649 6201 -1615
rect 6285 -1649 6319 -1615
rect 6403 -1649 6437 -1615
rect 6521 -1649 6555 -1615
rect 6639 -1649 6673 -1615
rect 6757 -1649 6791 -1615
rect 6875 -1649 6909 -1615
rect 6993 -1649 7027 -1615
rect 7111 -1649 7145 -1615
rect 7229 -1649 7263 -1615
rect 7347 -1649 7381 -1615
rect 7465 -1649 7499 -1615
rect 7583 -1649 7617 -1615
rect 7701 -1649 7735 -1615
rect 7819 -1649 7853 -1615
rect 7937 -1649 7971 -1615
rect 8055 -1649 8089 -1615
rect 8173 -1649 8207 -1615
rect 8291 -1649 8325 -1615
rect 8409 -1649 8443 -1615
rect 8527 -1649 8561 -1615
rect 8645 -1649 8679 -1615
rect 8763 -1649 8797 -1615
rect 8881 -1649 8915 -1615
rect 8999 -1649 9033 -1615
rect 9117 -1649 9151 -1615
rect 9235 -1649 9269 -1615
rect 9353 -1649 9387 -1615
rect 9471 -1649 9505 -1615
rect 9589 -1649 9623 -1615
rect 9707 -1649 9741 -1615
rect 9825 -1649 9859 -1615
rect 9943 -1649 9977 -1615
rect 10061 -1649 10095 -1615
rect 10179 -1649 10213 -1615
rect 10297 -1649 10331 -1615
rect 10415 -1649 10449 -1615
rect 10533 -1649 10567 -1615
rect 10651 -1649 10685 -1615
rect 4810 -2284 4844 -1708
rect 4928 -2284 4962 -1708
rect 5046 -2284 5080 -1708
rect 5164 -2284 5198 -1708
rect 5282 -2284 5316 -1708
rect 5400 -2284 5434 -1708
rect 5518 -2284 5552 -1708
rect 5636 -2284 5670 -1708
rect 5754 -2284 5788 -1708
rect 5872 -2284 5906 -1708
rect 5990 -2284 6024 -1708
rect 6108 -2284 6142 -1708
rect 6226 -2284 6260 -1708
rect 6344 -2284 6378 -1708
rect 6462 -2284 6496 -1708
rect 6580 -2284 6614 -1708
rect 6698 -2284 6732 -1708
rect 6816 -2284 6850 -1708
rect 6934 -2284 6968 -1708
rect 7052 -2284 7086 -1708
rect 7170 -2284 7204 -1708
rect 7288 -2284 7322 -1708
rect 7406 -2284 7440 -1708
rect 7524 -2284 7558 -1708
rect 7642 -2284 7676 -1708
rect 7760 -2284 7794 -1708
rect 7878 -2284 7912 -1708
rect 7996 -2284 8030 -1708
rect 8114 -2284 8148 -1708
rect 8232 -2284 8266 -1708
rect 8350 -2284 8384 -1708
rect 8468 -2284 8502 -1708
rect 8586 -2284 8620 -1708
rect 8704 -2284 8738 -1708
rect 8822 -2284 8856 -1708
rect 8940 -2284 8974 -1708
rect 9058 -2284 9092 -1708
rect 9176 -2284 9210 -1708
rect 9294 -2284 9328 -1708
rect 9412 -2284 9446 -1708
rect 9530 -2284 9564 -1708
rect 9648 -2284 9682 -1708
rect 9766 -2284 9800 -1708
rect 9884 -2284 9918 -1708
rect 10002 -2284 10036 -1708
rect 10120 -2284 10154 -1708
rect 10238 -2284 10272 -1708
rect 10356 -2284 10390 -1708
rect 10474 -2284 10508 -1708
rect 10592 -2284 10626 -1708
rect 10710 -2284 10744 -1708
rect 4776 -2479 4792 -2445
rect 4792 -2479 4810 -2445
rect 4848 -2479 4882 -2445
rect 4920 -2479 4954 -2445
rect 4992 -2479 5026 -2445
rect 5064 -2479 5098 -2445
rect 5136 -2479 5170 -2445
rect 5208 -2479 5242 -2445
rect 5280 -2479 5314 -2445
rect 5352 -2479 5386 -2445
rect 5424 -2479 5458 -2445
rect 5496 -2479 5530 -2445
rect 5568 -2479 5602 -2445
rect 5640 -2479 5674 -2445
rect 5712 -2479 5746 -2445
rect 5784 -2479 5818 -2445
rect 5856 -2479 5890 -2445
rect 5928 -2479 5962 -2445
rect 6000 -2479 6034 -2445
rect 6072 -2479 6106 -2445
rect 6144 -2479 6178 -2445
rect 6216 -2479 6250 -2445
rect 6288 -2479 6322 -2445
rect 6360 -2479 6394 -2445
rect 6432 -2479 6466 -2445
rect 6504 -2479 6538 -2445
rect 6576 -2479 6610 -2445
rect 6648 -2479 6682 -2445
rect 6720 -2479 6754 -2445
rect 6792 -2479 6826 -2445
rect 6864 -2479 6898 -2445
rect 6936 -2479 6970 -2445
rect 7008 -2479 7042 -2445
rect 7080 -2479 7114 -2445
rect 7152 -2479 7186 -2445
rect 7224 -2479 7258 -2445
rect 7296 -2479 7330 -2445
rect 7368 -2479 7402 -2445
rect 7440 -2479 7474 -2445
rect 7512 -2479 7546 -2445
rect 7584 -2479 7618 -2445
rect 7656 -2479 7690 -2445
rect 7728 -2479 7762 -2445
rect 7800 -2479 7834 -2445
rect 7872 -2479 7906 -2445
rect 7944 -2479 7978 -2445
rect 8016 -2479 8050 -2445
rect 8088 -2479 8122 -2445
rect 8160 -2479 8194 -2445
rect 8232 -2479 8266 -2445
rect 8304 -2479 8338 -2445
rect 8376 -2479 8410 -2445
rect 8448 -2479 8482 -2445
rect 8520 -2479 8554 -2445
rect 8592 -2479 8626 -2445
rect 8664 -2479 8698 -2445
rect 8736 -2479 8770 -2445
rect 8808 -2479 8842 -2445
rect 8880 -2479 8914 -2445
rect 8952 -2479 8986 -2445
rect 9024 -2479 9058 -2445
rect 9096 -2479 9130 -2445
rect 9168 -2479 9202 -2445
rect 9240 -2479 9274 -2445
rect 9312 -2479 9346 -2445
rect 9384 -2479 9418 -2445
rect 9456 -2479 9490 -2445
rect 9528 -2479 9562 -2445
rect 9600 -2479 9634 -2445
rect 9672 -2479 9706 -2445
rect 9744 -2479 9778 -2445
rect 9816 -2479 9850 -2445
rect 9888 -2479 9922 -2445
rect 9960 -2479 9994 -2445
rect 10032 -2479 10066 -2445
rect 10104 -2479 10138 -2445
rect 10176 -2479 10210 -2445
rect 10248 -2479 10282 -2445
rect 10320 -2479 10354 -2445
rect 10392 -2479 10426 -2445
rect 10464 -2479 10498 -2445
rect 10536 -2479 10570 -2445
rect 10608 -2479 10642 -2445
rect 10680 -2479 10714 -2445
rect 10752 -2479 10762 -2445
rect 10762 -2479 10786 -2445
rect 4776 -2567 4792 -2533
rect 4792 -2567 4810 -2533
rect 4848 -2567 4882 -2533
rect 4920 -2567 4954 -2533
rect 4992 -2567 5026 -2533
rect 5064 -2567 5098 -2533
rect 5136 -2567 5170 -2533
rect 5208 -2567 5242 -2533
rect 5280 -2567 5314 -2533
rect 5352 -2567 5386 -2533
rect 5424 -2567 5458 -2533
rect 5496 -2567 5530 -2533
rect 5568 -2567 5602 -2533
rect 5640 -2567 5674 -2533
rect 5712 -2567 5746 -2533
rect 5784 -2567 5818 -2533
rect 5856 -2567 5890 -2533
rect 5928 -2567 5962 -2533
rect 6000 -2567 6034 -2533
rect 6072 -2567 6106 -2533
rect 6144 -2567 6178 -2533
rect 6216 -2567 6250 -2533
rect 6288 -2567 6322 -2533
rect 6360 -2567 6394 -2533
rect 6432 -2567 6466 -2533
rect 6504 -2567 6538 -2533
rect 6576 -2567 6610 -2533
rect 6648 -2567 6682 -2533
rect 6720 -2567 6754 -2533
rect 6792 -2567 6826 -2533
rect 6864 -2567 6898 -2533
rect 6936 -2567 6970 -2533
rect 7008 -2567 7042 -2533
rect 7080 -2567 7114 -2533
rect 7152 -2567 7186 -2533
rect 7224 -2567 7258 -2533
rect 7296 -2567 7330 -2533
rect 7368 -2567 7402 -2533
rect 7440 -2567 7474 -2533
rect 7512 -2567 7546 -2533
rect 7584 -2567 7618 -2533
rect 7656 -2567 7690 -2533
rect 7728 -2567 7762 -2533
rect 7800 -2567 7834 -2533
rect 7872 -2567 7906 -2533
rect 7944 -2567 7978 -2533
rect 8016 -2567 8050 -2533
rect 8088 -2567 8122 -2533
rect 8160 -2567 8194 -2533
rect 8232 -2567 8266 -2533
rect 8304 -2567 8338 -2533
rect 8376 -2567 8410 -2533
rect 8448 -2567 8482 -2533
rect 8520 -2567 8554 -2533
rect 8592 -2567 8626 -2533
rect 8664 -2567 8698 -2533
rect 8736 -2567 8770 -2533
rect 8808 -2567 8842 -2533
rect 8880 -2567 8914 -2533
rect 8952 -2567 8986 -2533
rect 9024 -2567 9058 -2533
rect 9096 -2567 9130 -2533
rect 9168 -2567 9202 -2533
rect 9240 -2567 9274 -2533
rect 9312 -2567 9346 -2533
rect 9384 -2567 9418 -2533
rect 9456 -2567 9490 -2533
rect 9528 -2567 9562 -2533
rect 9600 -2567 9634 -2533
rect 9672 -2567 9706 -2533
rect 9744 -2567 9778 -2533
rect 9816 -2567 9850 -2533
rect 9888 -2567 9922 -2533
rect 9960 -2567 9994 -2533
rect 10032 -2567 10066 -2533
rect 10104 -2567 10138 -2533
rect 10176 -2567 10210 -2533
rect 10248 -2567 10282 -2533
rect 10320 -2567 10354 -2533
rect 10392 -2567 10426 -2533
rect 10464 -2567 10498 -2533
rect 10536 -2567 10570 -2533
rect 10608 -2567 10642 -2533
rect 10680 -2567 10714 -2533
rect 10752 -2567 10762 -2533
rect 10762 -2567 10786 -2533
rect 4776 -2655 4792 -2621
rect 4792 -2655 4810 -2621
rect 4848 -2655 4882 -2621
rect 4920 -2655 4954 -2621
rect 4992 -2655 5026 -2621
rect 5064 -2655 5098 -2621
rect 5136 -2655 5170 -2621
rect 5208 -2655 5242 -2621
rect 5280 -2655 5314 -2621
rect 5352 -2655 5386 -2621
rect 5424 -2655 5458 -2621
rect 5496 -2655 5530 -2621
rect 5568 -2655 5602 -2621
rect 5640 -2655 5674 -2621
rect 5712 -2655 5746 -2621
rect 5784 -2655 5818 -2621
rect 5856 -2655 5890 -2621
rect 5928 -2655 5962 -2621
rect 6000 -2655 6034 -2621
rect 6072 -2655 6106 -2621
rect 6144 -2655 6178 -2621
rect 6216 -2655 6250 -2621
rect 6288 -2655 6322 -2621
rect 6360 -2655 6394 -2621
rect 6432 -2655 6466 -2621
rect 6504 -2655 6538 -2621
rect 6576 -2655 6610 -2621
rect 6648 -2655 6682 -2621
rect 6720 -2655 6754 -2621
rect 6792 -2655 6826 -2621
rect 6864 -2655 6898 -2621
rect 6936 -2655 6970 -2621
rect 7008 -2655 7042 -2621
rect 7080 -2655 7114 -2621
rect 7152 -2655 7186 -2621
rect 7224 -2655 7258 -2621
rect 7296 -2655 7330 -2621
rect 7368 -2655 7402 -2621
rect 7440 -2655 7474 -2621
rect 7512 -2655 7546 -2621
rect 7584 -2655 7618 -2621
rect 7656 -2655 7690 -2621
rect 7728 -2655 7762 -2621
rect 7800 -2655 7834 -2621
rect 7872 -2655 7906 -2621
rect 7944 -2655 7978 -2621
rect 8016 -2655 8050 -2621
rect 8088 -2655 8122 -2621
rect 8160 -2655 8194 -2621
rect 8232 -2655 8266 -2621
rect 8304 -2655 8338 -2621
rect 8376 -2655 8410 -2621
rect 8448 -2655 8482 -2621
rect 8520 -2655 8554 -2621
rect 8592 -2655 8626 -2621
rect 8664 -2655 8698 -2621
rect 8736 -2655 8770 -2621
rect 8808 -2655 8842 -2621
rect 8880 -2655 8914 -2621
rect 8952 -2655 8986 -2621
rect 9024 -2655 9058 -2621
rect 9096 -2655 9130 -2621
rect 9168 -2655 9202 -2621
rect 9240 -2655 9274 -2621
rect 9312 -2655 9346 -2621
rect 9384 -2655 9418 -2621
rect 9456 -2655 9490 -2621
rect 9528 -2655 9562 -2621
rect 9600 -2655 9634 -2621
rect 9672 -2655 9706 -2621
rect 9744 -2655 9778 -2621
rect 9816 -2655 9850 -2621
rect 9888 -2655 9922 -2621
rect 9960 -2655 9994 -2621
rect 10032 -2655 10066 -2621
rect 10104 -2655 10138 -2621
rect 10176 -2655 10210 -2621
rect 10248 -2655 10282 -2621
rect 10320 -2655 10354 -2621
rect 10392 -2655 10426 -2621
rect 10464 -2655 10498 -2621
rect 10536 -2655 10570 -2621
rect 10608 -2655 10642 -2621
rect 10680 -2655 10714 -2621
rect 10752 -2655 10762 -2621
rect 10762 -2655 10786 -2621
rect 4810 -3498 4844 -2922
rect 4928 -3498 4962 -2922
rect 5046 -3498 5080 -2922
rect 5164 -3498 5198 -2922
rect 5282 -3498 5316 -2922
rect 5400 -3498 5434 -2922
rect 5518 -3498 5552 -2922
rect 5636 -3498 5670 -2922
rect 5754 -3498 5788 -2922
rect 5872 -3498 5906 -2922
rect 5990 -3498 6024 -2922
rect 6108 -3498 6142 -2922
rect 6226 -3498 6260 -2922
rect 6344 -3498 6378 -2922
rect 6462 -3498 6496 -2922
rect 6580 -3498 6614 -2922
rect 6698 -3498 6732 -2922
rect 6816 -3498 6850 -2922
rect 6934 -3498 6968 -2922
rect 7052 -3498 7086 -2922
rect 7170 -3498 7204 -2922
rect 7288 -3498 7322 -2922
rect 7406 -3498 7440 -2922
rect 7524 -3498 7558 -2922
rect 7642 -3498 7676 -2922
rect 7760 -3498 7794 -2922
rect 7878 -3498 7912 -2922
rect 7996 -3498 8030 -2922
rect 8114 -3498 8148 -2922
rect 8232 -3498 8266 -2922
rect 8350 -3498 8384 -2922
rect 8468 -3498 8502 -2922
rect 8586 -3498 8620 -2922
rect 8704 -3498 8738 -2922
rect 8822 -3498 8856 -2922
rect 8940 -3498 8974 -2922
rect 9058 -3498 9092 -2922
rect 9176 -3498 9210 -2922
rect 9294 -3498 9328 -2922
rect 9412 -3498 9446 -2922
rect 9530 -3498 9564 -2922
rect 9648 -3498 9682 -2922
rect 9766 -3498 9800 -2922
rect 9884 -3498 9918 -2922
rect 10002 -3498 10036 -2922
rect 10120 -3498 10154 -2922
rect 10238 -3498 10272 -2922
rect 10356 -3498 10390 -2922
rect 10474 -3498 10508 -2922
rect 10592 -3498 10626 -2922
rect 10710 -3498 10744 -2922
rect 4869 -3591 4903 -3557
rect 4987 -3591 5021 -3557
rect 5105 -3591 5139 -3557
rect 5223 -3591 5257 -3557
rect 5341 -3591 5375 -3557
rect 5459 -3591 5493 -3557
rect 5577 -3591 5611 -3557
rect 5695 -3591 5729 -3557
rect 5813 -3591 5847 -3557
rect 5931 -3591 5965 -3557
rect 6049 -3591 6083 -3557
rect 6167 -3591 6201 -3557
rect 6285 -3591 6319 -3557
rect 6403 -3591 6437 -3557
rect 6521 -3591 6555 -3557
rect 6639 -3591 6673 -3557
rect 6757 -3591 6791 -3557
rect 6875 -3591 6909 -3557
rect 6993 -3591 7027 -3557
rect 7111 -3591 7145 -3557
rect 7229 -3591 7263 -3557
rect 7347 -3591 7381 -3557
rect 7465 -3591 7499 -3557
rect 7583 -3591 7617 -3557
rect 7701 -3591 7735 -3557
rect 7819 -3591 7853 -3557
rect 7937 -3591 7971 -3557
rect 8055 -3591 8089 -3557
rect 8173 -3591 8207 -3557
rect 8291 -3591 8325 -3557
rect 8409 -3591 8443 -3557
rect 8527 -3591 8561 -3557
rect 8645 -3591 8679 -3557
rect 8763 -3591 8797 -3557
rect 8881 -3591 8915 -3557
rect 8999 -3591 9033 -3557
rect 9117 -3591 9151 -3557
rect 9235 -3591 9269 -3557
rect 9353 -3591 9387 -3557
rect 9471 -3591 9505 -3557
rect 9589 -3591 9623 -3557
rect 9707 -3591 9741 -3557
rect 9825 -3591 9859 -3557
rect 9943 -3591 9977 -3557
rect 10061 -3591 10095 -3557
rect 10179 -3591 10213 -3557
rect 10297 -3591 10331 -3557
rect 10415 -3591 10449 -3557
rect 10533 -3591 10567 -3557
rect 10651 -3591 10685 -3557
rect 4869 -3699 4903 -3665
rect 4987 -3699 5021 -3665
rect 5105 -3699 5139 -3665
rect 5223 -3699 5257 -3665
rect 5341 -3699 5375 -3665
rect 5459 -3699 5493 -3665
rect 5577 -3699 5611 -3665
rect 5695 -3699 5729 -3665
rect 5813 -3699 5847 -3665
rect 5931 -3699 5965 -3665
rect 6049 -3699 6083 -3665
rect 6167 -3699 6201 -3665
rect 6285 -3699 6319 -3665
rect 6403 -3699 6437 -3665
rect 6521 -3699 6555 -3665
rect 6639 -3699 6673 -3665
rect 6757 -3699 6791 -3665
rect 6875 -3699 6909 -3665
rect 6993 -3699 7027 -3665
rect 7111 -3699 7145 -3665
rect 7229 -3699 7263 -3665
rect 7347 -3699 7381 -3665
rect 7465 -3699 7499 -3665
rect 7583 -3699 7617 -3665
rect 7701 -3699 7735 -3665
rect 7819 -3699 7853 -3665
rect 7937 -3699 7971 -3665
rect 8055 -3699 8089 -3665
rect 8173 -3699 8207 -3665
rect 8291 -3699 8325 -3665
rect 8409 -3699 8443 -3665
rect 8527 -3699 8561 -3665
rect 8645 -3699 8679 -3665
rect 8763 -3699 8797 -3665
rect 8881 -3699 8915 -3665
rect 8999 -3699 9033 -3665
rect 9117 -3699 9151 -3665
rect 9235 -3699 9269 -3665
rect 9353 -3699 9387 -3665
rect 9471 -3699 9505 -3665
rect 9589 -3699 9623 -3665
rect 9707 -3699 9741 -3665
rect 9825 -3699 9859 -3665
rect 9943 -3699 9977 -3665
rect 10061 -3699 10095 -3665
rect 10179 -3699 10213 -3665
rect 10297 -3699 10331 -3665
rect 10415 -3699 10449 -3665
rect 10533 -3699 10567 -3665
rect 10651 -3699 10685 -3665
rect 4810 -4334 4844 -3758
rect 4928 -4334 4962 -3758
rect 5046 -4334 5080 -3758
rect 5164 -4334 5198 -3758
rect 5282 -4334 5316 -3758
rect 5400 -4334 5434 -3758
rect 5518 -4334 5552 -3758
rect 5636 -4334 5670 -3758
rect 5754 -4334 5788 -3758
rect 5872 -4334 5906 -3758
rect 5990 -4334 6024 -3758
rect 6108 -4334 6142 -3758
rect 6226 -4334 6260 -3758
rect 6344 -4334 6378 -3758
rect 6462 -4334 6496 -3758
rect 6580 -4334 6614 -3758
rect 6698 -4334 6732 -3758
rect 6816 -4334 6850 -3758
rect 6934 -4334 6968 -3758
rect 7052 -4334 7086 -3758
rect 7170 -4334 7204 -3758
rect 7288 -4334 7322 -3758
rect 7406 -4334 7440 -3758
rect 7524 -4334 7558 -3758
rect 7642 -4334 7676 -3758
rect 7760 -4334 7794 -3758
rect 7878 -4334 7912 -3758
rect 7996 -4334 8030 -3758
rect 8114 -4334 8148 -3758
rect 8232 -4334 8266 -3758
rect 8350 -4334 8384 -3758
rect 8468 -4334 8502 -3758
rect 8586 -4334 8620 -3758
rect 8704 -4334 8738 -3758
rect 8822 -4334 8856 -3758
rect 8940 -4334 8974 -3758
rect 9058 -4334 9092 -3758
rect 9176 -4334 9210 -3758
rect 9294 -4334 9328 -3758
rect 9412 -4334 9446 -3758
rect 9530 -4334 9564 -3758
rect 9648 -4334 9682 -3758
rect 9766 -4334 9800 -3758
rect 9884 -4334 9918 -3758
rect 10002 -4334 10036 -3758
rect 10120 -4334 10154 -3758
rect 10238 -4334 10272 -3758
rect 10356 -4334 10390 -3758
rect 10474 -4334 10508 -3758
rect 10592 -4334 10626 -3758
rect 10710 -4334 10744 -3758
rect 4768 -4529 4792 -4495
rect 4792 -4529 4802 -4495
rect 4840 -4529 4874 -4495
rect 4912 -4529 4946 -4495
rect 4984 -4529 5018 -4495
rect 5056 -4529 5090 -4495
rect 5128 -4529 5162 -4495
rect 5200 -4529 5234 -4495
rect 5272 -4529 5306 -4495
rect 5344 -4529 5378 -4495
rect 5416 -4529 5450 -4495
rect 5488 -4529 5522 -4495
rect 5560 -4529 5594 -4495
rect 5632 -4529 5666 -4495
rect 5704 -4529 5738 -4495
rect 5776 -4529 5810 -4495
rect 5848 -4529 5882 -4495
rect 5920 -4529 5954 -4495
rect 5992 -4529 6026 -4495
rect 6064 -4529 6098 -4495
rect 6136 -4529 6170 -4495
rect 6208 -4529 6242 -4495
rect 6280 -4529 6314 -4495
rect 6352 -4529 6386 -4495
rect 6424 -4529 6458 -4495
rect 6496 -4529 6530 -4495
rect 6568 -4529 6602 -4495
rect 6640 -4529 6674 -4495
rect 6712 -4529 6746 -4495
rect 6784 -4529 6818 -4495
rect 6856 -4529 6890 -4495
rect 6928 -4529 6962 -4495
rect 7000 -4529 7034 -4495
rect 7072 -4529 7106 -4495
rect 7144 -4529 7178 -4495
rect 7216 -4529 7250 -4495
rect 7288 -4529 7322 -4495
rect 7360 -4529 7394 -4495
rect 7432 -4529 7466 -4495
rect 7504 -4529 7538 -4495
rect 7576 -4529 7610 -4495
rect 7648 -4529 7682 -4495
rect 7720 -4529 7754 -4495
rect 7792 -4529 7826 -4495
rect 7864 -4529 7898 -4495
rect 7936 -4529 7970 -4495
rect 8008 -4529 8042 -4495
rect 8080 -4529 8114 -4495
rect 8152 -4529 8186 -4495
rect 8224 -4529 8258 -4495
rect 8296 -4529 8330 -4495
rect 8368 -4529 8402 -4495
rect 8440 -4529 8474 -4495
rect 8512 -4529 8546 -4495
rect 8584 -4529 8618 -4495
rect 8656 -4529 8690 -4495
rect 8728 -4529 8762 -4495
rect 8800 -4529 8834 -4495
rect 8872 -4529 8906 -4495
rect 8944 -4529 8978 -4495
rect 9016 -4529 9050 -4495
rect 9088 -4529 9122 -4495
rect 9160 -4529 9194 -4495
rect 9232 -4529 9266 -4495
rect 9304 -4529 9338 -4495
rect 9376 -4529 9410 -4495
rect 9448 -4529 9482 -4495
rect 9520 -4529 9554 -4495
rect 9592 -4529 9626 -4495
rect 9664 -4529 9698 -4495
rect 9736 -4529 9770 -4495
rect 9808 -4529 9842 -4495
rect 9880 -4529 9914 -4495
rect 9952 -4529 9986 -4495
rect 10024 -4529 10058 -4495
rect 10096 -4529 10130 -4495
rect 10168 -4529 10202 -4495
rect 10240 -4529 10274 -4495
rect 10312 -4529 10346 -4495
rect 10384 -4529 10418 -4495
rect 10456 -4529 10490 -4495
rect 10528 -4529 10562 -4495
rect 10600 -4529 10634 -4495
rect 10672 -4529 10706 -4495
rect 10744 -4529 10762 -4495
rect 10762 -4529 10778 -4495
rect 4768 -4617 4792 -4583
rect 4792 -4617 4802 -4583
rect 4840 -4617 4874 -4583
rect 4912 -4617 4946 -4583
rect 4984 -4617 5018 -4583
rect 5056 -4617 5090 -4583
rect 5128 -4617 5162 -4583
rect 5200 -4617 5234 -4583
rect 5272 -4617 5306 -4583
rect 5344 -4617 5378 -4583
rect 5416 -4617 5450 -4583
rect 5488 -4617 5522 -4583
rect 5560 -4617 5594 -4583
rect 5632 -4617 5666 -4583
rect 5704 -4617 5738 -4583
rect 5776 -4617 5810 -4583
rect 5848 -4617 5882 -4583
rect 5920 -4617 5954 -4583
rect 5992 -4617 6026 -4583
rect 6064 -4617 6098 -4583
rect 6136 -4617 6170 -4583
rect 6208 -4617 6242 -4583
rect 6280 -4617 6314 -4583
rect 6352 -4617 6386 -4583
rect 6424 -4617 6458 -4583
rect 6496 -4617 6530 -4583
rect 6568 -4617 6602 -4583
rect 6640 -4617 6674 -4583
rect 6712 -4617 6746 -4583
rect 6784 -4617 6818 -4583
rect 6856 -4617 6890 -4583
rect 6928 -4617 6962 -4583
rect 7000 -4617 7034 -4583
rect 7072 -4617 7106 -4583
rect 7144 -4617 7178 -4583
rect 7216 -4617 7250 -4583
rect 7288 -4617 7322 -4583
rect 7360 -4617 7394 -4583
rect 7432 -4617 7466 -4583
rect 7504 -4617 7538 -4583
rect 7576 -4617 7610 -4583
rect 7648 -4617 7682 -4583
rect 7720 -4617 7754 -4583
rect 7792 -4617 7826 -4583
rect 7864 -4617 7898 -4583
rect 7936 -4617 7970 -4583
rect 8008 -4617 8042 -4583
rect 8080 -4617 8114 -4583
rect 8152 -4617 8186 -4583
rect 8224 -4617 8258 -4583
rect 8296 -4617 8330 -4583
rect 8368 -4617 8402 -4583
rect 8440 -4617 8474 -4583
rect 8512 -4617 8546 -4583
rect 8584 -4617 8618 -4583
rect 8656 -4617 8690 -4583
rect 8728 -4617 8762 -4583
rect 8800 -4617 8834 -4583
rect 8872 -4617 8906 -4583
rect 8944 -4617 8978 -4583
rect 9016 -4617 9050 -4583
rect 9088 -4617 9122 -4583
rect 9160 -4617 9194 -4583
rect 9232 -4617 9266 -4583
rect 9304 -4617 9338 -4583
rect 9376 -4617 9410 -4583
rect 9448 -4617 9482 -4583
rect 9520 -4617 9554 -4583
rect 9592 -4617 9626 -4583
rect 9664 -4617 9698 -4583
rect 9736 -4617 9770 -4583
rect 9808 -4617 9842 -4583
rect 9880 -4617 9914 -4583
rect 9952 -4617 9986 -4583
rect 10024 -4617 10058 -4583
rect 10096 -4617 10130 -4583
rect 10168 -4617 10202 -4583
rect 10240 -4617 10274 -4583
rect 10312 -4617 10346 -4583
rect 10384 -4617 10418 -4583
rect 10456 -4617 10490 -4583
rect 10528 -4617 10562 -4583
rect 10600 -4617 10634 -4583
rect 10672 -4617 10706 -4583
rect 10744 -4617 10762 -4583
rect 10762 -4617 10778 -4583
rect 4768 -4705 4792 -4671
rect 4792 -4705 4802 -4671
rect 4840 -4705 4874 -4671
rect 4912 -4705 4946 -4671
rect 4984 -4705 5018 -4671
rect 5056 -4705 5090 -4671
rect 5128 -4705 5162 -4671
rect 5200 -4705 5234 -4671
rect 5272 -4705 5306 -4671
rect 5344 -4705 5378 -4671
rect 5416 -4705 5450 -4671
rect 5488 -4705 5522 -4671
rect 5560 -4705 5594 -4671
rect 5632 -4705 5666 -4671
rect 5704 -4705 5738 -4671
rect 5776 -4705 5810 -4671
rect 5848 -4705 5882 -4671
rect 5920 -4705 5954 -4671
rect 5992 -4705 6026 -4671
rect 6064 -4705 6098 -4671
rect 6136 -4705 6170 -4671
rect 6208 -4705 6242 -4671
rect 6280 -4705 6314 -4671
rect 6352 -4705 6386 -4671
rect 6424 -4705 6458 -4671
rect 6496 -4705 6530 -4671
rect 6568 -4705 6602 -4671
rect 6640 -4705 6674 -4671
rect 6712 -4705 6746 -4671
rect 6784 -4705 6818 -4671
rect 6856 -4705 6890 -4671
rect 6928 -4705 6962 -4671
rect 7000 -4705 7034 -4671
rect 7072 -4705 7106 -4671
rect 7144 -4705 7178 -4671
rect 7216 -4705 7250 -4671
rect 7288 -4705 7322 -4671
rect 7360 -4705 7394 -4671
rect 7432 -4705 7466 -4671
rect 7504 -4705 7538 -4671
rect 7576 -4705 7610 -4671
rect 7648 -4705 7682 -4671
rect 7720 -4705 7754 -4671
rect 7792 -4705 7826 -4671
rect 7864 -4705 7898 -4671
rect 7936 -4705 7970 -4671
rect 8008 -4705 8042 -4671
rect 8080 -4705 8114 -4671
rect 8152 -4705 8186 -4671
rect 8224 -4705 8258 -4671
rect 8296 -4705 8330 -4671
rect 8368 -4705 8402 -4671
rect 8440 -4705 8474 -4671
rect 8512 -4705 8546 -4671
rect 8584 -4705 8618 -4671
rect 8656 -4705 8690 -4671
rect 8728 -4705 8762 -4671
rect 8800 -4705 8834 -4671
rect 8872 -4705 8906 -4671
rect 8944 -4705 8978 -4671
rect 9016 -4705 9050 -4671
rect 9088 -4705 9122 -4671
rect 9160 -4705 9194 -4671
rect 9232 -4705 9266 -4671
rect 9304 -4705 9338 -4671
rect 9376 -4705 9410 -4671
rect 9448 -4705 9482 -4671
rect 9520 -4705 9554 -4671
rect 9592 -4705 9626 -4671
rect 9664 -4705 9698 -4671
rect 9736 -4705 9770 -4671
rect 9808 -4705 9842 -4671
rect 9880 -4705 9914 -4671
rect 9952 -4705 9986 -4671
rect 10024 -4705 10058 -4671
rect 10096 -4705 10130 -4671
rect 10168 -4705 10202 -4671
rect 10240 -4705 10274 -4671
rect 10312 -4705 10346 -4671
rect 10384 -4705 10418 -4671
rect 10456 -4705 10490 -4671
rect 10528 -4705 10562 -4671
rect 10600 -4705 10634 -4671
rect 10672 -4705 10706 -4671
rect 10744 -4705 10762 -4671
rect 10762 -4705 10778 -4671
rect 5046 -5548 5080 -4972
rect 5164 -5548 5198 -4972
rect 5282 -5548 5316 -4972
rect 5400 -5548 5434 -4972
rect 5518 -5548 5552 -4972
rect 5636 -5548 5670 -4972
rect 5754 -5548 5788 -4972
rect 5872 -5548 5906 -4972
rect 5990 -5548 6024 -4972
rect 6108 -5548 6142 -4972
rect 6226 -5548 6260 -4972
rect 6344 -5548 6378 -4972
rect 6462 -5548 6496 -4972
rect 6580 -5548 6614 -4972
rect 6698 -5548 6732 -4972
rect 6816 -5548 6850 -4972
rect 6934 -5548 6968 -4972
rect 7052 -5548 7086 -4972
rect 7170 -5548 7204 -4972
rect 7288 -5548 7322 -4972
rect 7406 -5548 7440 -4972
rect 7524 -5548 7558 -4972
rect 7642 -5548 7676 -4972
rect 7760 -5548 7794 -4972
rect 7878 -5548 7912 -4972
rect 7996 -5548 8030 -4972
rect 8114 -5548 8148 -4972
rect 8232 -5548 8266 -4972
rect 8350 -5548 8384 -4972
rect 8468 -5548 8502 -4972
rect 8586 -5548 8620 -4972
rect 8704 -5548 8738 -4972
rect 8822 -5548 8856 -4972
rect 8940 -5548 8974 -4972
rect 9058 -5548 9092 -4972
rect 9176 -5548 9210 -4972
rect 9294 -5548 9328 -4972
rect 9412 -5548 9446 -4972
rect 9530 -5548 9564 -4972
rect 9648 -5548 9682 -4972
rect 9766 -5548 9800 -4972
rect 9884 -5548 9918 -4972
rect 10002 -5548 10036 -4972
rect 10120 -5548 10154 -4972
rect 10238 -5548 10272 -4972
rect 10356 -5548 10390 -4972
rect 10474 -5548 10508 -4972
rect 10592 -5548 10626 -4972
rect 10710 -5548 10744 -4972
rect 4869 -5641 4903 -5607
rect 4987 -5641 5021 -5607
rect 5105 -5641 5139 -5607
rect 5223 -5641 5257 -5607
rect 5341 -5641 5375 -5607
rect 5459 -5641 5493 -5607
rect 5577 -5641 5611 -5607
rect 5695 -5641 5729 -5607
rect 5813 -5641 5847 -5607
rect 5931 -5641 5965 -5607
rect 6049 -5641 6083 -5607
rect 6167 -5641 6201 -5607
rect 6285 -5641 6319 -5607
rect 6403 -5641 6437 -5607
rect 6521 -5641 6555 -5607
rect 6639 -5641 6673 -5607
rect 6757 -5641 6791 -5607
rect 6875 -5641 6909 -5607
rect 6993 -5641 7027 -5607
rect 7111 -5641 7145 -5607
rect 7229 -5641 7263 -5607
rect 7347 -5641 7381 -5607
rect 7465 -5641 7499 -5607
rect 7583 -5641 7617 -5607
rect 7701 -5641 7735 -5607
rect 7819 -5641 7853 -5607
rect 7937 -5641 7971 -5607
rect 8055 -5641 8089 -5607
rect 8173 -5641 8207 -5607
rect 8291 -5641 8325 -5607
rect 8409 -5641 8443 -5607
rect 8527 -5641 8561 -5607
rect 8645 -5641 8679 -5607
rect 8763 -5641 8797 -5607
rect 8881 -5641 8915 -5607
rect 8999 -5641 9033 -5607
rect 9117 -5641 9151 -5607
rect 9235 -5641 9269 -5607
rect 9353 -5641 9387 -5607
rect 9471 -5641 9505 -5607
rect 9589 -5641 9623 -5607
rect 9707 -5641 9741 -5607
rect 9825 -5641 9859 -5607
rect 9943 -5641 9977 -5607
rect 10061 -5641 10095 -5607
rect 10179 -5641 10213 -5607
rect 10297 -5641 10331 -5607
rect 10415 -5641 10449 -5607
rect 10533 -5641 10567 -5607
rect 10651 -5641 10685 -5607
rect 4869 -5749 4903 -5715
rect 4987 -5749 5021 -5715
rect 5105 -5749 5139 -5715
rect 5223 -5749 5257 -5715
rect 5341 -5749 5375 -5715
rect 5459 -5749 5493 -5715
rect 5577 -5749 5611 -5715
rect 5695 -5749 5729 -5715
rect 5813 -5749 5847 -5715
rect 5931 -5749 5965 -5715
rect 6049 -5749 6083 -5715
rect 6167 -5749 6201 -5715
rect 6285 -5749 6319 -5715
rect 6403 -5749 6437 -5715
rect 6521 -5749 6555 -5715
rect 6639 -5749 6673 -5715
rect 6757 -5749 6791 -5715
rect 6875 -5749 6909 -5715
rect 6993 -5749 7027 -5715
rect 7111 -5749 7145 -5715
rect 7229 -5749 7263 -5715
rect 7347 -5749 7381 -5715
rect 7465 -5749 7499 -5715
rect 7583 -5749 7617 -5715
rect 7701 -5749 7735 -5715
rect 7819 -5749 7853 -5715
rect 7937 -5749 7971 -5715
rect 8055 -5749 8089 -5715
rect 8173 -5749 8207 -5715
rect 8291 -5749 8325 -5715
rect 8409 -5749 8443 -5715
rect 8527 -5749 8561 -5715
rect 8645 -5749 8679 -5715
rect 8763 -5749 8797 -5715
rect 8881 -5749 8915 -5715
rect 8999 -5749 9033 -5715
rect 9117 -5749 9151 -5715
rect 9235 -5749 9269 -5715
rect 9353 -5749 9387 -5715
rect 9471 -5749 9505 -5715
rect 9589 -5749 9623 -5715
rect 9707 -5749 9741 -5715
rect 9825 -5749 9859 -5715
rect 9943 -5749 9977 -5715
rect 10061 -5749 10095 -5715
rect 10179 -5749 10213 -5715
rect 10297 -5749 10331 -5715
rect 10415 -5749 10449 -5715
rect 10533 -5749 10567 -5715
rect 10651 -5749 10685 -5715
rect 4810 -6384 4844 -5808
rect 4928 -6384 4962 -5808
rect 5046 -6384 5080 -5808
rect 5164 -6384 5198 -5808
rect 5282 -6384 5316 -5808
rect 5400 -6384 5434 -5808
rect 5518 -6384 5552 -5808
rect 5636 -6384 5670 -5808
rect 5754 -6384 5788 -5808
rect 5872 -6384 5906 -5808
rect 5990 -6384 6024 -5808
rect 6108 -6384 6142 -5808
rect 6226 -6384 6260 -5808
rect 6344 -6384 6378 -5808
rect 6462 -6384 6496 -5808
rect 6580 -6384 6614 -5808
rect 6698 -6384 6732 -5808
rect 6816 -6384 6850 -5808
rect 6934 -6384 6968 -5808
rect 7052 -6384 7086 -5808
rect 7170 -6384 7204 -5808
rect 7288 -6384 7322 -5808
rect 7406 -6384 7440 -5808
rect 7524 -6384 7558 -5808
rect 7642 -6384 7676 -5808
rect 7760 -6384 7794 -5808
rect 7878 -6384 7912 -5808
rect 7996 -6384 8030 -5808
rect 8114 -6384 8148 -5808
rect 8232 -6384 8266 -5808
rect 8350 -6384 8384 -5808
rect 8468 -6384 8502 -5808
rect 8586 -6384 8620 -5808
rect 8704 -6384 8738 -5808
rect 8822 -6384 8856 -5808
rect 8940 -6384 8974 -5808
rect 9058 -6384 9092 -5808
rect 9176 -6384 9210 -5808
rect 9294 -6384 9328 -5808
rect 9412 -6384 9446 -5808
rect 9530 -6384 9564 -5808
rect 9648 -6384 9682 -5808
rect 9766 -6384 9800 -5808
rect 9884 -6384 9918 -5808
rect 10002 -6384 10036 -5808
rect 10120 -6384 10154 -5808
rect 10238 -6384 10272 -5808
rect 10356 -6384 10390 -5808
rect 10474 -6384 10508 -5808
rect 10592 -6384 10626 -5808
rect 10710 -6384 10744 -5808
rect 4098 -7159 4132 -7125
rect 4170 -7159 4204 -7125
rect 4242 -7159 4276 -7125
rect 4314 -7159 4348 -7125
rect 4386 -7159 4420 -7125
rect 4458 -7159 4492 -7125
rect 4530 -7159 4564 -7125
rect 4602 -7159 4636 -7125
rect 4674 -7159 4708 -7125
rect 4746 -7159 4780 -7125
rect 4818 -7159 4852 -7125
rect 4890 -7159 4924 -7125
rect 4962 -7159 4996 -7125
rect 5034 -7159 5068 -7125
rect 5106 -7159 5140 -7125
rect 5178 -7159 5212 -7125
rect 5250 -7159 5284 -7125
rect 5322 -7159 5356 -7125
rect 5394 -7159 5428 -7125
rect 5466 -7159 5500 -7125
rect 5538 -7159 5572 -7125
rect 4098 -7233 4132 -7199
rect 4170 -7233 4204 -7199
rect 4242 -7233 4276 -7199
rect 4314 -7233 4348 -7199
rect 4386 -7233 4420 -7199
rect 4458 -7233 4492 -7199
rect 4530 -7233 4564 -7199
rect 4602 -7233 4636 -7199
rect 4674 -7233 4708 -7199
rect 4746 -7233 4780 -7199
rect 4818 -7233 4852 -7199
rect 4890 -7233 4924 -7199
rect 4962 -7233 4996 -7199
rect 5034 -7233 5068 -7199
rect 5106 -7233 5140 -7199
rect 5178 -7233 5212 -7199
rect 5250 -7233 5284 -7199
rect 5322 -7233 5356 -7199
rect 5394 -7233 5428 -7199
rect 5466 -7233 5500 -7199
rect 5538 -7233 5572 -7199
rect 4098 -7307 4132 -7273
rect 4170 -7307 4204 -7273
rect 4242 -7307 4276 -7273
rect 4314 -7307 4348 -7273
rect 4386 -7307 4420 -7273
rect 4458 -7307 4492 -7273
rect 4530 -7307 4564 -7273
rect 4602 -7307 4636 -7273
rect 4674 -7307 4708 -7273
rect 4746 -7307 4780 -7273
rect 4818 -7307 4852 -7273
rect 4890 -7307 4924 -7273
rect 4962 -7307 4996 -7273
rect 5034 -7307 5068 -7273
rect 5106 -7307 5140 -7273
rect 5178 -7307 5212 -7273
rect 5250 -7307 5284 -7273
rect 5322 -7307 5356 -7273
rect 5394 -7307 5428 -7273
rect 5466 -7307 5500 -7273
rect 5538 -7307 5572 -7273
rect 4098 -7381 4132 -7347
rect 4170 -7381 4204 -7347
rect 4242 -7381 4276 -7347
rect 4314 -7381 4348 -7347
rect 4386 -7381 4420 -7347
rect 4458 -7381 4492 -7347
rect 4530 -7381 4564 -7347
rect 4602 -7381 4636 -7347
rect 4674 -7381 4708 -7347
rect 4746 -7381 4780 -7347
rect 4818 -7381 4852 -7347
rect 4890 -7381 4924 -7347
rect 4962 -7381 4996 -7347
rect 5034 -7381 5068 -7347
rect 5106 -7381 5140 -7347
rect 5178 -7381 5212 -7347
rect 5250 -7381 5284 -7347
rect 5322 -7381 5356 -7347
rect 5394 -7381 5428 -7347
rect 5466 -7381 5500 -7347
rect 5538 -7381 5572 -7347
rect 4098 -7455 4132 -7421
rect 4170 -7455 4204 -7421
rect 4242 -7455 4276 -7421
rect 4314 -7455 4348 -7421
rect 4386 -7455 4420 -7421
rect 4458 -7455 4492 -7421
rect 4530 -7455 4564 -7421
rect 4602 -7455 4636 -7421
rect 4674 -7455 4708 -7421
rect 4746 -7455 4780 -7421
rect 4818 -7455 4852 -7421
rect 4890 -7455 4924 -7421
rect 4962 -7455 4996 -7421
rect 5034 -7455 5068 -7421
rect 5106 -7455 5140 -7421
rect 5178 -7455 5212 -7421
rect 5250 -7455 5284 -7421
rect 5322 -7455 5356 -7421
rect 5394 -7455 5428 -7421
rect 5466 -7455 5500 -7421
rect 5538 -7455 5572 -7421
rect 4098 -7529 4132 -7495
rect 4170 -7529 4204 -7495
rect 4242 -7529 4276 -7495
rect 4314 -7529 4348 -7495
rect 4386 -7529 4420 -7495
rect 4458 -7529 4492 -7495
rect 4530 -7529 4564 -7495
rect 4602 -7529 4636 -7495
rect 4674 -7529 4708 -7495
rect 4746 -7529 4780 -7495
rect 4818 -7529 4852 -7495
rect 4890 -7529 4924 -7495
rect 4962 -7529 4996 -7495
rect 5034 -7529 5068 -7495
rect 5106 -7529 5140 -7495
rect 5178 -7529 5212 -7495
rect 5250 -7529 5284 -7495
rect 5322 -7529 5356 -7495
rect 5394 -7529 5428 -7495
rect 5466 -7529 5500 -7495
rect 5538 -7529 5572 -7495
rect 4098 -7603 4132 -7569
rect 4170 -7603 4204 -7569
rect 4242 -7603 4276 -7569
rect 4314 -7603 4348 -7569
rect 4386 -7603 4420 -7569
rect 4458 -7603 4492 -7569
rect 4530 -7603 4564 -7569
rect 4602 -7603 4636 -7569
rect 4674 -7603 4708 -7569
rect 4746 -7603 4780 -7569
rect 4818 -7603 4852 -7569
rect 4890 -7603 4924 -7569
rect 4962 -7603 4996 -7569
rect 5034 -7603 5068 -7569
rect 5106 -7603 5140 -7569
rect 5178 -7603 5212 -7569
rect 5250 -7603 5284 -7569
rect 5322 -7603 5356 -7569
rect 5394 -7603 5428 -7569
rect 5466 -7603 5500 -7569
rect 5538 -7603 5572 -7569
rect 4098 -7677 4132 -7643
rect 4170 -7677 4204 -7643
rect 4242 -7677 4276 -7643
rect 4314 -7677 4348 -7643
rect 4386 -7677 4420 -7643
rect 4458 -7677 4492 -7643
rect 4530 -7677 4564 -7643
rect 4602 -7677 4636 -7643
rect 4674 -7677 4708 -7643
rect 4746 -7677 4780 -7643
rect 4818 -7677 4852 -7643
rect 4890 -7677 4924 -7643
rect 4962 -7677 4996 -7643
rect 5034 -7677 5068 -7643
rect 5106 -7677 5140 -7643
rect 5178 -7677 5212 -7643
rect 5250 -7677 5284 -7643
rect 5322 -7677 5356 -7643
rect 5394 -7677 5428 -7643
rect 5466 -7677 5500 -7643
rect 5538 -7677 5572 -7643
rect 4098 -7751 4132 -7717
rect 4170 -7751 4204 -7717
rect 4242 -7751 4276 -7717
rect 4314 -7751 4348 -7717
rect 4386 -7751 4420 -7717
rect 4458 -7751 4492 -7717
rect 4530 -7751 4564 -7717
rect 4602 -7751 4636 -7717
rect 4674 -7751 4708 -7717
rect 4746 -7751 4780 -7717
rect 4818 -7751 4852 -7717
rect 4890 -7751 4924 -7717
rect 4962 -7751 4996 -7717
rect 5034 -7751 5068 -7717
rect 5106 -7751 5140 -7717
rect 5178 -7751 5212 -7717
rect 5250 -7751 5284 -7717
rect 5322 -7751 5356 -7717
rect 5394 -7751 5428 -7717
rect 5466 -7751 5500 -7717
rect 5538 -7751 5572 -7717
rect 6112 -7791 6146 -7215
rect 6230 -7791 6264 -7215
rect 6348 -7791 6382 -7215
rect 6466 -7791 6500 -7215
rect 6584 -7791 6618 -7215
rect 6702 -7791 6736 -7215
rect 6820 -7791 6854 -7215
rect 6938 -7791 6972 -7215
rect 7056 -7791 7090 -7215
rect 7174 -7791 7208 -7215
rect 7292 -7791 7326 -7215
rect 7410 -7791 7444 -7215
rect 7528 -7791 7562 -7215
rect 7646 -7791 7680 -7215
rect 7874 -7791 7908 -7215
rect 7992 -7791 8026 -7215
rect 8110 -7791 8144 -7215
rect 8228 -7791 8262 -7215
rect 8346 -7791 8380 -7215
rect 8464 -7791 8498 -7215
rect 8582 -7791 8616 -7215
rect 8700 -7791 8734 -7215
rect 8818 -7791 8852 -7215
rect 8936 -7791 8970 -7215
rect 9054 -7791 9088 -7215
rect 9172 -7791 9206 -7215
rect 9290 -7791 9324 -7215
rect 9408 -7791 9442 -7215
rect 9526 -7791 9560 -7215
rect 9644 -7791 9678 -7215
rect 9834 -7223 9868 -7189
rect 9906 -7223 9940 -7189
rect 9978 -7223 10012 -7189
rect 10050 -7223 10084 -7189
rect 10122 -7223 10156 -7189
rect 10194 -7223 10228 -7189
rect 10266 -7223 10300 -7189
rect 10421 -7225 10455 -7191
rect 10737 -7225 10771 -7191
rect 11053 -7225 11087 -7191
rect 11369 -7225 11403 -7191
rect 11685 -7225 11719 -7191
rect 12001 -7225 12035 -7191
rect 12317 -7225 12351 -7191
rect 9834 -7297 9868 -7263
rect 9906 -7297 9940 -7263
rect 9978 -7297 10012 -7263
rect 10050 -7297 10084 -7263
rect 10122 -7297 10156 -7263
rect 10194 -7297 10228 -7263
rect 10266 -7297 10300 -7263
rect 10421 -7298 10455 -7264
rect 9834 -7371 9868 -7337
rect 9906 -7371 9940 -7337
rect 9978 -7371 10012 -7337
rect 10050 -7371 10084 -7337
rect 10122 -7371 10156 -7337
rect 10194 -7371 10228 -7337
rect 10266 -7371 10300 -7337
rect 10421 -7371 10455 -7337
rect 9834 -7445 9868 -7411
rect 9906 -7445 9940 -7411
rect 9978 -7445 10012 -7411
rect 10050 -7445 10084 -7411
rect 10122 -7445 10156 -7411
rect 10194 -7445 10228 -7411
rect 10266 -7445 10300 -7411
rect 10421 -7444 10455 -7410
rect 9834 -7519 9868 -7485
rect 9906 -7519 9940 -7485
rect 9978 -7519 10012 -7485
rect 10050 -7519 10084 -7485
rect 10122 -7519 10156 -7485
rect 10194 -7519 10228 -7485
rect 10266 -7519 10300 -7485
rect 10421 -7517 10455 -7483
rect 9834 -7593 9868 -7559
rect 9906 -7593 9940 -7559
rect 9978 -7593 10012 -7559
rect 10050 -7593 10084 -7559
rect 10122 -7593 10156 -7559
rect 10194 -7593 10228 -7559
rect 10266 -7593 10300 -7559
rect 10421 -7590 10455 -7556
rect 9834 -7667 9868 -7633
rect 9906 -7667 9940 -7633
rect 9978 -7667 10012 -7633
rect 10050 -7667 10084 -7633
rect 10122 -7667 10156 -7633
rect 10194 -7667 10228 -7633
rect 10266 -7667 10300 -7633
rect 10737 -7287 10771 -7264
rect 10737 -7298 10771 -7287
rect 10737 -7371 10771 -7337
rect 11053 -7287 11087 -7264
rect 11053 -7298 11087 -7287
rect 10737 -7444 10771 -7410
rect 10737 -7517 10771 -7483
rect 10851 -7503 10885 -7377
rect 10939 -7503 10973 -7377
rect 11053 -7371 11087 -7337
rect 11369 -7287 11403 -7264
rect 11369 -7298 11403 -7287
rect 11053 -7444 11087 -7410
rect 11053 -7517 11087 -7483
rect 10737 -7590 10771 -7556
rect 11167 -7503 11201 -7377
rect 11255 -7503 11289 -7377
rect 11369 -7371 11403 -7337
rect 11685 -7287 11719 -7264
rect 11685 -7298 11719 -7287
rect 11369 -7444 11403 -7410
rect 11369 -7517 11403 -7483
rect 11053 -7590 11087 -7556
rect 11483 -7503 11517 -7377
rect 11571 -7503 11605 -7377
rect 11685 -7371 11719 -7337
rect 12001 -7287 12035 -7264
rect 12001 -7298 12035 -7287
rect 11685 -7444 11719 -7410
rect 11685 -7517 11719 -7483
rect 11369 -7590 11403 -7556
rect 11799 -7503 11833 -7377
rect 11887 -7503 11921 -7377
rect 12001 -7371 12035 -7337
rect 12317 -7287 12351 -7264
rect 12317 -7298 12351 -7287
rect 12001 -7444 12035 -7410
rect 12001 -7517 12035 -7483
rect 11685 -7590 11719 -7556
rect 12115 -7503 12149 -7377
rect 12203 -7503 12237 -7377
rect 12317 -7371 12351 -7337
rect 12317 -7444 12351 -7410
rect 12317 -7517 12351 -7483
rect 12001 -7590 12035 -7556
rect 12317 -7590 12351 -7556
rect 10421 -7689 10455 -7655
rect 10494 -7689 10528 -7655
rect 10567 -7689 10601 -7655
rect 10640 -7689 10674 -7655
rect 10713 -7689 10747 -7655
rect 10786 -7689 10820 -7655
rect 10859 -7689 10893 -7655
rect 10932 -7689 10966 -7655
rect 11005 -7689 11039 -7655
rect 11078 -7689 11112 -7655
rect 11151 -7689 11185 -7655
rect 11224 -7689 11258 -7655
rect 11297 -7689 11331 -7655
rect 11370 -7689 11404 -7655
rect 11443 -7689 11477 -7655
rect 11516 -7689 11550 -7655
rect 11589 -7689 11623 -7655
rect 11662 -7689 11696 -7655
rect 11735 -7689 11769 -7655
rect 11808 -7689 11842 -7655
rect 11881 -7689 11915 -7655
rect 11954 -7689 11988 -7655
rect 12027 -7689 12061 -7655
rect 12100 -7689 12134 -7655
rect 12173 -7689 12207 -7655
rect 12246 -7689 12280 -7655
rect 12319 -7689 12353 -7655
rect 9834 -7741 9868 -7707
rect 9906 -7741 9940 -7707
rect 9978 -7741 10012 -7707
rect 10050 -7741 10084 -7707
rect 10122 -7741 10156 -7707
rect 10194 -7741 10228 -7707
rect 10266 -7741 10300 -7707
rect 4098 -7825 4132 -7791
rect 4170 -7825 4204 -7791
rect 4242 -7825 4276 -7791
rect 4314 -7825 4348 -7791
rect 4386 -7825 4420 -7791
rect 4458 -7825 4492 -7791
rect 4530 -7825 4564 -7791
rect 4602 -7825 4636 -7791
rect 4674 -7825 4708 -7791
rect 4746 -7825 4780 -7791
rect 4818 -7825 4852 -7791
rect 4890 -7825 4924 -7791
rect 4962 -7825 4996 -7791
rect 5034 -7825 5068 -7791
rect 5106 -7825 5140 -7791
rect 5178 -7825 5212 -7791
rect 5250 -7825 5284 -7791
rect 5322 -7825 5356 -7791
rect 5394 -7825 5428 -7791
rect 5466 -7825 5500 -7791
rect 5538 -7825 5572 -7791
rect 9834 -7815 9868 -7781
rect 9906 -7815 9940 -7781
rect 9978 -7815 10012 -7781
rect 10050 -7815 10084 -7781
rect 10122 -7815 10156 -7781
rect 10194 -7815 10228 -7781
rect 10266 -7815 10300 -7781
rect 10338 -7815 10372 -7781
rect 10410 -7815 10444 -7781
rect 10482 -7815 10516 -7781
rect 10554 -7815 10588 -7781
rect 4098 -7899 4132 -7865
rect 4170 -7899 4204 -7865
rect 4242 -7899 4276 -7865
rect 4314 -7899 4348 -7865
rect 4386 -7899 4420 -7865
rect 4458 -7899 4492 -7865
rect 4530 -7899 4564 -7865
rect 4602 -7899 4636 -7865
rect 4674 -7899 4708 -7865
rect 4746 -7899 4780 -7865
rect 4818 -7899 4852 -7865
rect 4890 -7899 4924 -7865
rect 4962 -7899 4996 -7865
rect 5034 -7899 5068 -7865
rect 5106 -7899 5140 -7865
rect 5178 -7899 5212 -7865
rect 5250 -7899 5284 -7865
rect 5322 -7899 5356 -7865
rect 5394 -7899 5428 -7865
rect 5466 -7899 5500 -7865
rect 5538 -7899 5572 -7865
rect 5935 -7875 5969 -7841
rect 6053 -7875 6087 -7841
rect 6171 -7875 6205 -7841
rect 6289 -7875 6323 -7841
rect 6407 -7875 6441 -7841
rect 6525 -7875 6559 -7841
rect 6643 -7875 6677 -7841
rect 6761 -7875 6795 -7841
rect 6879 -7875 6913 -7841
rect 6997 -7875 7031 -7841
rect 7115 -7875 7149 -7841
rect 7233 -7875 7267 -7841
rect 7351 -7875 7385 -7841
rect 7469 -7875 7503 -7841
rect 7587 -7875 7621 -7841
rect 7933 -7875 7967 -7841
rect 8051 -7875 8085 -7841
rect 8169 -7875 8203 -7841
rect 8287 -7875 8321 -7841
rect 8405 -7875 8439 -7841
rect 8523 -7875 8557 -7841
rect 8641 -7875 8675 -7841
rect 8759 -7875 8793 -7841
rect 8877 -7875 8911 -7841
rect 8995 -7875 9029 -7841
rect 9113 -7875 9147 -7841
rect 9231 -7875 9265 -7841
rect 9349 -7875 9383 -7841
rect 9467 -7875 9501 -7841
rect 9585 -7875 9619 -7841
rect 9834 -7889 9868 -7855
rect 9906 -7889 9940 -7855
rect 9978 -7889 10012 -7855
rect 10050 -7889 10084 -7855
rect 10122 -7889 10156 -7855
rect 10194 -7889 10228 -7855
rect 10266 -7889 10300 -7855
rect 10338 -7889 10372 -7855
rect 10410 -7889 10444 -7855
rect 10482 -7889 10516 -7855
rect 10554 -7889 10588 -7855
rect 4098 -7973 4132 -7939
rect 4170 -7973 4204 -7939
rect 4242 -7973 4276 -7939
rect 4314 -7973 4348 -7939
rect 4386 -7973 4420 -7939
rect 4458 -7973 4492 -7939
rect 4530 -7973 4564 -7939
rect 4602 -7973 4636 -7939
rect 4674 -7973 4708 -7939
rect 4746 -7973 4780 -7939
rect 4818 -7973 4852 -7939
rect 4890 -7973 4924 -7939
rect 4962 -7973 4996 -7939
rect 5034 -7973 5068 -7939
rect 5106 -7973 5140 -7939
rect 5178 -7973 5212 -7939
rect 5250 -7973 5284 -7939
rect 5322 -7973 5356 -7939
rect 5394 -7973 5428 -7939
rect 5466 -7973 5500 -7939
rect 5538 -7973 5572 -7939
rect 5935 -7983 5969 -7949
rect 6053 -7983 6087 -7949
rect 6171 -7983 6205 -7949
rect 6289 -7983 6323 -7949
rect 6407 -7983 6441 -7949
rect 6525 -7983 6559 -7949
rect 6643 -7983 6677 -7949
rect 6761 -7983 6795 -7949
rect 6879 -7983 6913 -7949
rect 6997 -7983 7031 -7949
rect 7115 -7983 7149 -7949
rect 7233 -7983 7267 -7949
rect 7351 -7983 7385 -7949
rect 7469 -7983 7503 -7949
rect 7587 -7983 7621 -7949
rect 7933 -7983 7967 -7949
rect 8051 -7983 8085 -7949
rect 8169 -7983 8203 -7949
rect 8287 -7983 8321 -7949
rect 8405 -7983 8439 -7949
rect 8523 -7983 8557 -7949
rect 8641 -7983 8675 -7949
rect 8759 -7983 8793 -7949
rect 8877 -7983 8911 -7949
rect 8995 -7983 9029 -7949
rect 9113 -7983 9147 -7949
rect 9231 -7983 9265 -7949
rect 9349 -7983 9383 -7949
rect 9467 -7983 9501 -7949
rect 9585 -7983 9619 -7949
rect 9834 -7963 9868 -7929
rect 9906 -7963 9940 -7929
rect 9978 -7963 10012 -7929
rect 10050 -7963 10084 -7929
rect 10122 -7963 10156 -7929
rect 10194 -7963 10228 -7929
rect 10266 -7963 10300 -7929
rect 10338 -7963 10372 -7929
rect 10410 -7963 10444 -7929
rect 4098 -8047 4132 -8013
rect 4170 -8047 4204 -8013
rect 4242 -8047 4276 -8013
rect 4314 -8047 4348 -8013
rect 4386 -8047 4420 -8013
rect 4458 -8047 4492 -8013
rect 4530 -8047 4564 -8013
rect 4602 -8047 4636 -8013
rect 4674 -8047 4708 -8013
rect 4746 -8047 4780 -8013
rect 4818 -8047 4852 -8013
rect 4890 -8047 4924 -8013
rect 4962 -8047 4996 -8013
rect 5034 -8047 5068 -8013
rect 5106 -8047 5140 -8013
rect 5178 -8047 5212 -8013
rect 5250 -8047 5284 -8013
rect 5322 -8047 5356 -8013
rect 5394 -8047 5428 -8013
rect 5466 -8047 5500 -8013
rect 5538 -8047 5572 -8013
rect 4098 -8121 4132 -8087
rect 4170 -8121 4204 -8087
rect 4242 -8121 4276 -8087
rect 4314 -8121 4348 -8087
rect 4386 -8121 4420 -8087
rect 4458 -8121 4492 -8087
rect 4530 -8121 4564 -8087
rect 4602 -8121 4636 -8087
rect 4674 -8121 4708 -8087
rect 4746 -8121 4780 -8087
rect 4818 -8121 4852 -8087
rect 4890 -8121 4924 -8087
rect 4962 -8121 4996 -8087
rect 5034 -8121 5068 -8087
rect 5106 -8121 5140 -8087
rect 5178 -8121 5212 -8087
rect 5250 -8121 5284 -8087
rect 5322 -8121 5356 -8087
rect 5394 -8121 5428 -8087
rect 5466 -8121 5500 -8087
rect 5538 -8121 5572 -8087
rect 4098 -8195 4132 -8161
rect 4170 -8195 4204 -8161
rect 4242 -8195 4276 -8161
rect 4314 -8195 4348 -8161
rect 4386 -8195 4420 -8161
rect 4458 -8195 4492 -8161
rect 4530 -8195 4564 -8161
rect 4602 -8195 4636 -8161
rect 4674 -8195 4708 -8161
rect 4746 -8195 4780 -8161
rect 4818 -8195 4852 -8161
rect 4890 -8195 4924 -8161
rect 4962 -8195 4996 -8161
rect 5034 -8195 5068 -8161
rect 5106 -8195 5140 -8161
rect 5178 -8195 5212 -8161
rect 5250 -8195 5284 -8161
rect 5322 -8195 5356 -8161
rect 5394 -8195 5428 -8161
rect 5466 -8195 5500 -8161
rect 5538 -8195 5572 -8161
rect 4098 -8269 4132 -8235
rect 4170 -8269 4204 -8235
rect 4242 -8269 4276 -8235
rect 4314 -8269 4348 -8235
rect 4386 -8269 4420 -8235
rect 4458 -8269 4492 -8235
rect 4530 -8269 4564 -8235
rect 4602 -8269 4636 -8235
rect 4674 -8269 4708 -8235
rect 4746 -8269 4780 -8235
rect 4818 -8269 4852 -8235
rect 4890 -8269 4924 -8235
rect 4962 -8269 4996 -8235
rect 5034 -8269 5068 -8235
rect 5106 -8269 5140 -8235
rect 5178 -8269 5212 -8235
rect 5250 -8269 5284 -8235
rect 5322 -8269 5356 -8235
rect 5394 -8269 5428 -8235
rect 5466 -8269 5500 -8235
rect 5538 -8269 5572 -8235
rect 4098 -8343 4132 -8309
rect 4170 -8343 4204 -8309
rect 4242 -8343 4276 -8309
rect 4314 -8343 4348 -8309
rect 4386 -8343 4420 -8309
rect 4458 -8343 4492 -8309
rect 4530 -8343 4564 -8309
rect 4602 -8343 4636 -8309
rect 4674 -8343 4708 -8309
rect 4746 -8343 4780 -8309
rect 4818 -8343 4852 -8309
rect 4890 -8343 4924 -8309
rect 4962 -8343 4996 -8309
rect 5034 -8343 5068 -8309
rect 5106 -8343 5140 -8309
rect 5178 -8343 5212 -8309
rect 5250 -8343 5284 -8309
rect 5322 -8343 5356 -8309
rect 5394 -8343 5428 -8309
rect 5466 -8343 5500 -8309
rect 5538 -8343 5572 -8309
rect 4098 -8417 4132 -8383
rect 4170 -8417 4204 -8383
rect 4242 -8417 4276 -8383
rect 4314 -8417 4348 -8383
rect 4386 -8417 4420 -8383
rect 4458 -8417 4492 -8383
rect 4530 -8417 4564 -8383
rect 4602 -8417 4636 -8383
rect 4674 -8417 4708 -8383
rect 4746 -8417 4780 -8383
rect 4818 -8417 4852 -8383
rect 4890 -8417 4924 -8383
rect 4962 -8417 4996 -8383
rect 5034 -8417 5068 -8383
rect 5106 -8417 5140 -8383
rect 5178 -8417 5212 -8383
rect 5250 -8417 5284 -8383
rect 5322 -8417 5356 -8383
rect 5394 -8417 5428 -8383
rect 5466 -8417 5500 -8383
rect 5538 -8417 5572 -8383
rect 4098 -8491 4132 -8457
rect 4170 -8491 4204 -8457
rect 4242 -8491 4276 -8457
rect 4314 -8491 4348 -8457
rect 4386 -8491 4420 -8457
rect 4458 -8491 4492 -8457
rect 4530 -8491 4564 -8457
rect 4602 -8491 4636 -8457
rect 4674 -8491 4708 -8457
rect 4746 -8491 4780 -8457
rect 4818 -8491 4852 -8457
rect 4890 -8491 4924 -8457
rect 4962 -8491 4996 -8457
rect 5034 -8491 5068 -8457
rect 5106 -8491 5140 -8457
rect 5178 -8491 5212 -8457
rect 5250 -8491 5284 -8457
rect 5322 -8491 5356 -8457
rect 5394 -8491 5428 -8457
rect 5466 -8491 5500 -8457
rect 5538 -8491 5572 -8457
rect 4098 -8565 4132 -8531
rect 4170 -8565 4204 -8531
rect 4242 -8565 4276 -8531
rect 4314 -8565 4348 -8531
rect 4386 -8565 4420 -8531
rect 4458 -8565 4492 -8531
rect 4530 -8565 4564 -8531
rect 4602 -8565 4636 -8531
rect 4674 -8565 4708 -8531
rect 4746 -8565 4780 -8531
rect 4818 -8565 4852 -8531
rect 4890 -8565 4924 -8531
rect 4962 -8565 4996 -8531
rect 5034 -8565 5068 -8531
rect 5106 -8565 5140 -8531
rect 5178 -8565 5212 -8531
rect 5250 -8565 5284 -8531
rect 5322 -8565 5356 -8531
rect 5394 -8565 5428 -8531
rect 5466 -8565 5500 -8531
rect 5538 -8565 5572 -8531
rect 5876 -8609 5910 -8033
rect 5994 -8609 6028 -8033
rect 6112 -8609 6146 -8033
rect 6230 -8609 6264 -8033
rect 6348 -8609 6382 -8033
rect 6466 -8609 6500 -8033
rect 6584 -8609 6618 -8033
rect 6702 -8609 6736 -8033
rect 6820 -8609 6854 -8033
rect 6938 -8609 6972 -8033
rect 7056 -8609 7090 -8033
rect 7174 -8609 7208 -8033
rect 7292 -8609 7326 -8033
rect 7410 -8609 7444 -8033
rect 7528 -8609 7562 -8033
rect 7646 -8609 7680 -8033
rect 7874 -8609 7908 -8033
rect 7992 -8609 8026 -8033
rect 8110 -8609 8144 -8033
rect 8228 -8609 8262 -8033
rect 8346 -8609 8380 -8033
rect 8464 -8609 8498 -8033
rect 8582 -8609 8616 -8033
rect 8700 -8609 8734 -8033
rect 8818 -8609 8852 -8033
rect 8936 -8609 8970 -8033
rect 9054 -8609 9088 -8033
rect 9172 -8609 9206 -8033
rect 9290 -8609 9324 -8033
rect 9408 -8609 9442 -8033
rect 9526 -8609 9560 -8033
rect 9644 -8609 9678 -8033
rect 9834 -8037 9868 -8003
rect 9906 -8037 9940 -8003
rect 9978 -8037 10012 -8003
rect 10050 -8037 10084 -8003
rect 10122 -8037 10156 -8003
rect 10194 -8037 10228 -8003
rect 10266 -8037 10300 -8003
rect 10338 -8037 10372 -8003
rect 10410 -8037 10444 -8003
rect 9834 -8111 9868 -8077
rect 9906 -8111 9940 -8077
rect 9978 -8111 10012 -8077
rect 10050 -8111 10084 -8077
rect 10122 -8111 10156 -8077
rect 10194 -8111 10228 -8077
rect 10266 -8111 10300 -8077
rect 10338 -8111 10372 -8077
rect 10410 -8111 10444 -8077
rect 12534 -8091 12568 -7215
rect 12682 -8091 12716 -7215
rect 12830 -8091 12864 -7215
rect 12978 -8091 13012 -7215
rect 13126 -8091 13160 -7215
rect 13274 -8091 13308 -7215
rect 13422 -8091 13456 -7215
rect 13570 -8091 13604 -7215
rect 13718 -8091 13752 -7215
rect 13866 -8091 13900 -7215
rect 14014 -8091 14048 -7215
rect 14162 -8091 14196 -7215
rect 14310 -8091 14344 -7215
rect 14458 -8091 14492 -7215
rect 14606 -8091 14640 -7215
rect 14754 -8091 14788 -7215
rect 14902 -8091 14936 -7215
rect 15050 -8091 15084 -7215
rect 15198 -8091 15232 -7215
rect 15346 -8091 15380 -7215
rect 15494 -8091 15528 -7215
rect 15642 -8091 15676 -7215
rect 15790 -8091 15824 -7215
rect 15938 -8091 15972 -7215
rect 16086 -8091 16120 -7215
rect 16234 -8091 16268 -7215
rect 16382 -8091 16416 -7215
rect 16530 -8091 16564 -7215
rect 16678 -8091 16712 -7215
rect 16826 -8091 16860 -7215
rect 16974 -8091 17008 -7215
rect 17122 -8091 17156 -7215
rect 17270 -8091 17304 -7215
rect 17418 -8091 17452 -7215
rect 17566 -8091 17600 -7215
rect 17714 -8091 17748 -7215
rect 17862 -8091 17896 -7215
rect 18010 -8091 18044 -7215
rect 18158 -8091 18192 -7215
rect 18306 -8091 18340 -7215
rect 18454 -8091 18488 -7215
rect 18602 -8091 18636 -7215
rect 18750 -8091 18784 -7215
rect 18898 -8091 18932 -7215
rect 19046 -8091 19080 -7215
rect 19194 -8091 19228 -7215
rect 19342 -8091 19376 -7215
rect 19490 -8091 19524 -7215
rect 19638 -8091 19672 -7215
rect 19786 -8091 19820 -7215
rect 19934 -8091 19968 -7215
rect 20082 -8091 20116 -7215
rect 20230 -8091 20264 -7215
rect 20378 -8091 20412 -7215
rect 20526 -8091 20560 -7215
rect 20674 -8091 20708 -7215
rect 20822 -8091 20856 -7215
rect 20970 -8091 21004 -7215
rect 21118 -8091 21152 -7215
rect 21266 -8091 21300 -7215
rect 21414 -8091 21448 -7215
rect 21562 -8091 21596 -7215
rect 21710 -8091 21744 -7215
rect 21858 -8091 21892 -7215
rect 22006 -8091 22040 -7215
rect 22154 -8091 22188 -7215
rect 22302 -8091 22336 -7215
rect 22450 -8091 22484 -7215
rect 22598 -8091 22632 -7215
rect 22746 -8091 22780 -7215
rect 22894 -8091 22928 -7215
rect 23042 -8091 23076 -7215
rect 23190 -8091 23224 -7215
rect 23338 -8091 23372 -7215
rect 23634 -8091 23668 -7215
rect 9834 -8185 9868 -8151
rect 9906 -8185 9940 -8151
rect 9978 -8185 10012 -8151
rect 10050 -8185 10084 -8151
rect 10122 -8185 10156 -8151
rect 10194 -8185 10228 -8151
rect 10266 -8185 10300 -8151
rect 10338 -8185 10372 -8151
rect 10410 -8185 10444 -8151
rect 12744 -8175 12802 -8141
rect 12892 -8175 12950 -8141
rect 13040 -8175 13098 -8141
rect 13188 -8175 13246 -8141
rect 13336 -8175 13394 -8141
rect 13484 -8175 13542 -8141
rect 13632 -8175 13690 -8141
rect 13780 -8175 13838 -8141
rect 13928 -8175 13986 -8141
rect 14076 -8175 14134 -8141
rect 14224 -8175 14282 -8141
rect 14372 -8175 14430 -8141
rect 14520 -8175 14578 -8141
rect 14668 -8175 14726 -8141
rect 14816 -8175 14874 -8141
rect 14964 -8175 15022 -8141
rect 15112 -8175 15170 -8141
rect 15260 -8175 15318 -8141
rect 15408 -8175 15466 -8141
rect 15556 -8175 15614 -8141
rect 15704 -8175 15762 -8141
rect 15852 -8175 15910 -8141
rect 16000 -8175 16058 -8141
rect 16148 -8175 16206 -8141
rect 16296 -8175 16354 -8141
rect 16444 -8175 16502 -8141
rect 16592 -8175 16650 -8141
rect 16740 -8175 16798 -8141
rect 16888 -8175 16946 -8141
rect 17036 -8175 17094 -8141
rect 17184 -8175 17242 -8141
rect 17332 -8175 17390 -8141
rect 17480 -8175 17538 -8141
rect 17628 -8175 17686 -8141
rect 17776 -8175 17834 -8141
rect 17924 -8175 17982 -8141
rect 18072 -8175 18130 -8141
rect 18220 -8175 18278 -8141
rect 18368 -8175 18426 -8141
rect 18516 -8175 18574 -8141
rect 18664 -8175 18722 -8141
rect 18812 -8175 18870 -8141
rect 18960 -8175 19018 -8141
rect 19108 -8175 19166 -8141
rect 19256 -8175 19314 -8141
rect 19404 -8175 19462 -8141
rect 19552 -8175 19610 -8141
rect 19700 -8175 19758 -8141
rect 19848 -8175 19906 -8141
rect 19996 -8175 20054 -8141
rect 20144 -8175 20202 -8141
rect 20292 -8175 20350 -8141
rect 20440 -8175 20498 -8141
rect 20588 -8175 20646 -8141
rect 20736 -8175 20794 -8141
rect 20884 -8175 20942 -8141
rect 21032 -8175 21090 -8141
rect 21180 -8175 21238 -8141
rect 21328 -8175 21386 -8141
rect 21476 -8175 21534 -8141
rect 21624 -8175 21682 -8141
rect 21772 -8175 21830 -8141
rect 21920 -8175 21978 -8141
rect 22068 -8175 22126 -8141
rect 22216 -8175 22274 -8141
rect 22364 -8175 22422 -8141
rect 22512 -8175 22570 -8141
rect 22660 -8175 22718 -8141
rect 22808 -8175 22866 -8141
rect 22956 -8175 23014 -8141
rect 23104 -8175 23162 -8141
rect 23252 -8175 23310 -8141
rect 23400 -8175 23458 -8141
rect 23548 -8175 23606 -8141
rect 9834 -8259 9868 -8225
rect 9906 -8259 9940 -8225
rect 9978 -8259 10012 -8225
rect 10050 -8259 10084 -8225
rect 10122 -8259 10156 -8225
rect 10194 -8259 10228 -8225
rect 10266 -8259 10300 -8225
rect 10338 -8259 10372 -8225
rect 10410 -8259 10444 -8225
rect 12744 -8283 12802 -8249
rect 12892 -8283 12950 -8249
rect 13040 -8283 13098 -8249
rect 13188 -8283 13246 -8249
rect 13336 -8283 13394 -8249
rect 13484 -8283 13542 -8249
rect 13632 -8283 13690 -8249
rect 13780 -8283 13838 -8249
rect 13928 -8283 13986 -8249
rect 14076 -8283 14134 -8249
rect 14224 -8283 14282 -8249
rect 14372 -8283 14430 -8249
rect 14520 -8283 14578 -8249
rect 14668 -8283 14726 -8249
rect 14816 -8283 14874 -8249
rect 14964 -8283 15022 -8249
rect 15112 -8283 15170 -8249
rect 15260 -8283 15318 -8249
rect 15408 -8283 15466 -8249
rect 15556 -8283 15614 -8249
rect 15704 -8283 15762 -8249
rect 15852 -8283 15910 -8249
rect 16000 -8283 16058 -8249
rect 16148 -8283 16206 -8249
rect 16296 -8283 16354 -8249
rect 16444 -8283 16502 -8249
rect 16592 -8283 16650 -8249
rect 16740 -8283 16798 -8249
rect 16888 -8283 16946 -8249
rect 17036 -8283 17094 -8249
rect 17184 -8283 17242 -8249
rect 17332 -8283 17390 -8249
rect 17480 -8283 17538 -8249
rect 17628 -8283 17686 -8249
rect 17776 -8283 17834 -8249
rect 17924 -8283 17982 -8249
rect 18072 -8283 18130 -8249
rect 18220 -8283 18278 -8249
rect 18368 -8283 18426 -8249
rect 18516 -8283 18574 -8249
rect 18664 -8283 18722 -8249
rect 18812 -8283 18870 -8249
rect 18960 -8283 19018 -8249
rect 19108 -8283 19166 -8249
rect 19256 -8283 19314 -8249
rect 19404 -8283 19462 -8249
rect 19552 -8283 19610 -8249
rect 19700 -8283 19758 -8249
rect 19848 -8283 19906 -8249
rect 19996 -8283 20054 -8249
rect 20144 -8283 20202 -8249
rect 20292 -8283 20350 -8249
rect 20440 -8283 20498 -8249
rect 20588 -8283 20646 -8249
rect 20736 -8283 20794 -8249
rect 20884 -8283 20942 -8249
rect 21032 -8283 21090 -8249
rect 21180 -8283 21238 -8249
rect 21328 -8283 21386 -8249
rect 21476 -8283 21534 -8249
rect 21624 -8283 21682 -8249
rect 21772 -8283 21830 -8249
rect 21920 -8283 21978 -8249
rect 22068 -8283 22126 -8249
rect 22216 -8283 22274 -8249
rect 22364 -8283 22422 -8249
rect 22512 -8283 22570 -8249
rect 22660 -8283 22718 -8249
rect 22808 -8283 22866 -8249
rect 22956 -8283 23014 -8249
rect 23104 -8283 23162 -8249
rect 23252 -8283 23310 -8249
rect 23400 -8283 23458 -8249
rect 23548 -8283 23606 -8249
rect 9834 -8333 9868 -8299
rect 9906 -8333 9940 -8299
rect 9978 -8333 10012 -8299
rect 10050 -8333 10084 -8299
rect 10122 -8333 10156 -8299
rect 10194 -8333 10228 -8299
rect 10266 -8333 10300 -8299
rect 10338 -8333 10372 -8299
rect 10410 -8333 10444 -8299
rect 10482 -8333 10516 -8299
rect 10554 -8333 10588 -8299
rect 9834 -8407 9868 -8373
rect 9906 -8407 9940 -8373
rect 9978 -8407 10012 -8373
rect 10050 -8407 10084 -8373
rect 10122 -8407 10156 -8373
rect 10194 -8407 10228 -8373
rect 10266 -8407 10300 -8373
rect 10338 -8407 10372 -8373
rect 10410 -8407 10444 -8373
rect 10482 -8407 10516 -8373
rect 10554 -8407 10588 -8373
rect 9834 -8481 9868 -8447
rect 9906 -8481 9940 -8447
rect 9978 -8481 10012 -8447
rect 10050 -8481 10084 -8447
rect 10122 -8481 10156 -8447
rect 10194 -8481 10228 -8447
rect 10266 -8481 10300 -8447
rect 10338 -8481 10372 -8447
rect 10410 -8481 10444 -8447
rect 10482 -8481 10516 -8447
rect 10554 -8481 10588 -8447
rect 9834 -8555 9868 -8521
rect 9906 -8555 9940 -8521
rect 9978 -8555 10012 -8521
rect 10050 -8555 10084 -8521
rect 10122 -8555 10156 -8521
rect 10194 -8555 10228 -8521
rect 10266 -8555 10300 -8521
rect 10338 -8555 10372 -8521
rect 10410 -8555 10444 -8521
rect 10482 -8555 10516 -8521
rect 10554 -8555 10588 -8521
rect 9834 -8629 9868 -8595
rect 9906 -8629 9940 -8595
rect 9978 -8629 10012 -8595
rect 10050 -8629 10084 -8595
rect 10122 -8629 10156 -8595
rect 10194 -8629 10228 -8595
rect 10266 -8629 10300 -8595
rect 10338 -8629 10372 -8595
rect 10410 -8629 10444 -8595
rect 10482 -8629 10516 -8595
rect 10554 -8629 10588 -8595
rect 9834 -8703 9868 -8669
rect 9906 -8703 9940 -8669
rect 9978 -8703 10012 -8669
rect 10050 -8703 10084 -8669
rect 10122 -8703 10156 -8669
rect 10194 -8703 10228 -8669
rect 10266 -8703 10300 -8669
rect 10338 -8703 10372 -8669
rect 10410 -8703 10444 -8669
rect 10482 -8703 10516 -8669
rect 10554 -8703 10588 -8669
rect 4080 -8905 4114 -8871
rect 4152 -8905 4186 -8871
rect 4234 -8905 4268 -8871
rect 4306 -8905 4340 -8871
rect 4388 -8905 4422 -8871
rect 4460 -8905 4494 -8871
rect 4542 -8905 4576 -8871
rect 4614 -8905 4648 -8871
rect 4696 -8905 4730 -8871
rect 4768 -8905 4802 -8871
rect 4850 -8905 4884 -8871
rect 4922 -8905 4956 -8871
rect 5004 -8905 5038 -8871
rect 5076 -8905 5110 -8871
rect 5158 -8905 5192 -8871
rect 5230 -8905 5264 -8871
rect 5312 -8905 5346 -8871
rect 5384 -8905 5418 -8871
rect 5466 -8905 5500 -8871
rect 5538 -8905 5572 -8871
rect 5620 -8905 5654 -8871
rect 5692 -8905 5726 -8871
rect 4080 -8979 4114 -8945
rect 4152 -8979 4186 -8945
rect 4234 -8979 4268 -8945
rect 4306 -8979 4340 -8945
rect 4388 -8979 4422 -8945
rect 4460 -8979 4494 -8945
rect 4542 -8979 4576 -8945
rect 4614 -8979 4648 -8945
rect 4696 -8979 4730 -8945
rect 4768 -8979 4802 -8945
rect 4850 -8979 4884 -8945
rect 4922 -8979 4956 -8945
rect 5004 -8979 5038 -8945
rect 5076 -8979 5110 -8945
rect 5158 -8979 5192 -8945
rect 5230 -8979 5264 -8945
rect 5312 -8979 5346 -8945
rect 5384 -8979 5418 -8945
rect 5466 -8979 5500 -8945
rect 5538 -8979 5572 -8945
rect 5620 -8979 5654 -8945
rect 5692 -8979 5726 -8945
rect 5774 -8979 5808 -8945
rect 5846 -8979 5880 -8945
rect 5928 -8979 5962 -8945
rect 6000 -8979 6034 -8945
rect 6082 -8979 6116 -8945
rect 6154 -8979 6188 -8945
rect 6236 -8979 6270 -8945
rect 6308 -8979 6342 -8945
rect 6390 -8979 6424 -8945
rect 6462 -8979 6496 -8945
rect 6544 -8979 6578 -8945
rect 6616 -8979 6650 -8945
rect 6698 -8979 6732 -8945
rect 6770 -8979 6804 -8945
rect 6852 -8979 6886 -8945
rect 6924 -8979 6958 -8945
rect 7006 -8979 7040 -8945
rect 7078 -8979 7112 -8945
rect 7160 -8979 7194 -8945
rect 7232 -8979 7266 -8945
rect 7314 -8979 7348 -8945
rect 7386 -8979 7420 -8945
rect 7468 -8979 7502 -8945
rect 7540 -8979 7574 -8945
rect 7622 -8979 7656 -8945
rect 7694 -8979 7728 -8945
rect 7776 -8979 7810 -8945
rect 7848 -8979 7882 -8945
rect 7930 -8979 7964 -8945
rect 8002 -8979 8036 -8945
rect 8084 -8979 8118 -8945
rect 8156 -8979 8190 -8945
rect 8238 -8979 8272 -8945
rect 8310 -8979 8344 -8945
rect 8392 -8979 8426 -8945
rect 8464 -8979 8498 -8945
rect 8546 -8979 8580 -8945
rect 8618 -8979 8652 -8945
rect 8700 -8979 8734 -8945
rect 8772 -8979 8806 -8945
rect 8854 -8979 8888 -8945
rect 8926 -8979 8960 -8945
rect 9008 -8979 9042 -8945
rect 9080 -8979 9114 -8945
rect 9162 -8979 9196 -8945
rect 9234 -8979 9268 -8945
rect 9316 -8979 9350 -8945
rect 9388 -8979 9422 -8945
rect 9470 -8979 9504 -8945
rect 9542 -8979 9576 -8945
rect 9624 -8979 9658 -8945
rect 9696 -8979 9730 -8945
rect 9778 -8979 9812 -8945
rect 9850 -8979 9884 -8945
rect 9932 -8979 9966 -8945
rect 10004 -8979 10038 -8945
rect 10086 -8979 10120 -8945
rect 10158 -8979 10192 -8945
rect 10240 -8979 10274 -8945
rect 10312 -8979 10346 -8945
rect 10394 -8979 10428 -8945
rect 10466 -8979 10500 -8945
rect 10548 -8979 10582 -8945
rect 10620 -8979 10654 -8945
rect 10702 -8979 10736 -8945
rect 10774 -8979 10808 -8945
rect 10856 -8979 10890 -8945
rect 10928 -8979 10962 -8945
rect 11010 -8979 11044 -8945
rect 11082 -8979 11116 -8945
rect 11164 -8979 11198 -8945
rect 11236 -8979 11270 -8945
rect 11318 -8979 11352 -8945
rect 11390 -8979 11424 -8945
rect 11472 -8979 11506 -8945
rect 11544 -8979 11578 -8945
rect 11626 -8979 11660 -8945
rect 11698 -8979 11732 -8945
rect 11780 -8979 11814 -8945
rect 11852 -8979 11886 -8945
rect 11934 -8979 11968 -8945
rect 12006 -8979 12040 -8945
rect 4080 -9053 4114 -9019
rect 4152 -9053 4186 -9019
rect 4234 -9053 4268 -9019
rect 4306 -9053 4340 -9019
rect 4388 -9053 4422 -9019
rect 4460 -9053 4494 -9019
rect 4542 -9053 4576 -9019
rect 4614 -9053 4648 -9019
rect 4696 -9053 4730 -9019
rect 4768 -9053 4802 -9019
rect 4850 -9053 4884 -9019
rect 4922 -9053 4956 -9019
rect 5004 -9053 5038 -9019
rect 5076 -9053 5110 -9019
rect 5158 -9053 5192 -9019
rect 5230 -9053 5264 -9019
rect 5312 -9053 5346 -9019
rect 5384 -9053 5418 -9019
rect 5466 -9053 5500 -9019
rect 5538 -9053 5572 -9019
rect 5620 -9053 5654 -9019
rect 5692 -9053 5726 -9019
rect 5774 -9053 5808 -9019
rect 5846 -9053 5880 -9019
rect 5928 -9053 5962 -9019
rect 6000 -9053 6034 -9019
rect 6082 -9053 6116 -9019
rect 6154 -9053 6188 -9019
rect 6236 -9053 6270 -9019
rect 6308 -9053 6342 -9019
rect 6390 -9053 6424 -9019
rect 6462 -9053 6496 -9019
rect 6544 -9053 6578 -9019
rect 6616 -9053 6650 -9019
rect 6698 -9053 6732 -9019
rect 6770 -9053 6804 -9019
rect 6852 -9053 6886 -9019
rect 6924 -9053 6958 -9019
rect 7006 -9053 7040 -9019
rect 7078 -9053 7112 -9019
rect 7160 -9053 7194 -9019
rect 7232 -9053 7266 -9019
rect 7314 -9053 7348 -9019
rect 7386 -9053 7420 -9019
rect 7468 -9053 7502 -9019
rect 7540 -9053 7574 -9019
rect 7622 -9053 7656 -9019
rect 7694 -9053 7728 -9019
rect 7776 -9053 7810 -9019
rect 7848 -9053 7882 -9019
rect 7930 -9053 7964 -9019
rect 8002 -9053 8036 -9019
rect 8084 -9053 8118 -9019
rect 8156 -9053 8190 -9019
rect 8238 -9053 8272 -9019
rect 8310 -9053 8344 -9019
rect 8392 -9053 8426 -9019
rect 8464 -9053 8498 -9019
rect 8546 -9053 8580 -9019
rect 8618 -9053 8652 -9019
rect 8700 -9053 8734 -9019
rect 8772 -9053 8806 -9019
rect 8854 -9053 8888 -9019
rect 8926 -9053 8960 -9019
rect 9008 -9053 9042 -9019
rect 9080 -9053 9114 -9019
rect 9162 -9053 9196 -9019
rect 9234 -9053 9268 -9019
rect 9316 -9053 9350 -9019
rect 9388 -9053 9422 -9019
rect 9470 -9053 9504 -9019
rect 9542 -9053 9576 -9019
rect 9624 -9053 9658 -9019
rect 9696 -9053 9730 -9019
rect 9778 -9053 9812 -9019
rect 9850 -9053 9884 -9019
rect 9932 -9053 9966 -9019
rect 10004 -9053 10038 -9019
rect 10086 -9053 10120 -9019
rect 10158 -9053 10192 -9019
rect 10240 -9053 10274 -9019
rect 10312 -9053 10346 -9019
rect 10394 -9053 10428 -9019
rect 10466 -9053 10500 -9019
rect 10548 -9053 10582 -9019
rect 10620 -9053 10654 -9019
rect 10702 -9053 10736 -9019
rect 10774 -9053 10808 -9019
rect 10856 -9053 10890 -9019
rect 10928 -9053 10962 -9019
rect 11010 -9053 11044 -9019
rect 11082 -9053 11116 -9019
rect 11164 -9053 11198 -9019
rect 11236 -9053 11270 -9019
rect 11318 -9053 11352 -9019
rect 11390 -9053 11424 -9019
rect 11472 -9053 11506 -9019
rect 11544 -9053 11578 -9019
rect 11626 -9053 11660 -9019
rect 11698 -9053 11732 -9019
rect 11780 -9053 11814 -9019
rect 11852 -9053 11886 -9019
rect 11934 -9053 11968 -9019
rect 12006 -9053 12040 -9019
rect 4080 -9127 4114 -9093
rect 4152 -9127 4186 -9093
rect 4234 -9127 4268 -9093
rect 4306 -9127 4340 -9093
rect 4388 -9127 4422 -9093
rect 4460 -9127 4494 -9093
rect 4542 -9127 4576 -9093
rect 4614 -9127 4648 -9093
rect 4696 -9127 4730 -9093
rect 4768 -9127 4802 -9093
rect 4850 -9127 4884 -9093
rect 4922 -9127 4956 -9093
rect 5004 -9127 5038 -9093
rect 5076 -9127 5110 -9093
rect 5158 -9127 5192 -9093
rect 5230 -9127 5264 -9093
rect 5312 -9127 5346 -9093
rect 5384 -9127 5418 -9093
rect 5466 -9127 5500 -9093
rect 5538 -9127 5572 -9093
rect 5620 -9127 5654 -9093
rect 5692 -9127 5726 -9093
rect 5774 -9127 5808 -9093
rect 5846 -9127 5880 -9093
rect 5928 -9127 5962 -9093
rect 6000 -9127 6034 -9093
rect 6082 -9127 6116 -9093
rect 6154 -9127 6188 -9093
rect 6236 -9127 6270 -9093
rect 6308 -9127 6342 -9093
rect 6390 -9127 6424 -9093
rect 6462 -9127 6496 -9093
rect 6544 -9127 6578 -9093
rect 6616 -9127 6650 -9093
rect 6698 -9127 6732 -9093
rect 6770 -9127 6804 -9093
rect 6852 -9127 6886 -9093
rect 6924 -9127 6958 -9093
rect 7006 -9127 7040 -9093
rect 7078 -9127 7112 -9093
rect 7160 -9127 7194 -9093
rect 7232 -9127 7266 -9093
rect 7314 -9127 7348 -9093
rect 7386 -9127 7420 -9093
rect 7468 -9127 7502 -9093
rect 7540 -9127 7574 -9093
rect 7622 -9127 7656 -9093
rect 7694 -9127 7728 -9093
rect 7776 -9127 7810 -9093
rect 7848 -9127 7882 -9093
rect 7930 -9127 7964 -9093
rect 8002 -9127 8036 -9093
rect 8084 -9127 8118 -9093
rect 8156 -9127 8190 -9093
rect 8238 -9127 8272 -9093
rect 8310 -9127 8344 -9093
rect 8392 -9127 8426 -9093
rect 8464 -9127 8498 -9093
rect 8546 -9127 8580 -9093
rect 8618 -9127 8652 -9093
rect 8700 -9127 8734 -9093
rect 8772 -9127 8806 -9093
rect 8854 -9127 8888 -9093
rect 8926 -9127 8960 -9093
rect 9008 -9127 9042 -9093
rect 9080 -9127 9114 -9093
rect 9162 -9127 9196 -9093
rect 9234 -9127 9268 -9093
rect 9316 -9127 9350 -9093
rect 9388 -9127 9422 -9093
rect 9470 -9127 9504 -9093
rect 9542 -9127 9576 -9093
rect 9624 -9127 9658 -9093
rect 9696 -9127 9730 -9093
rect 9778 -9127 9812 -9093
rect 9850 -9127 9884 -9093
rect 9932 -9127 9966 -9093
rect 10004 -9127 10038 -9093
rect 10086 -9127 10120 -9093
rect 10158 -9127 10192 -9093
rect 10240 -9127 10274 -9093
rect 10312 -9127 10346 -9093
rect 10394 -9127 10428 -9093
rect 10466 -9127 10500 -9093
rect 10548 -9127 10582 -9093
rect 10620 -9127 10654 -9093
rect 10702 -9127 10736 -9093
rect 10774 -9127 10808 -9093
rect 10856 -9127 10890 -9093
rect 10928 -9127 10962 -9093
rect 11010 -9127 11044 -9093
rect 11082 -9127 11116 -9093
rect 11164 -9127 11198 -9093
rect 11236 -9127 11270 -9093
rect 11318 -9127 11352 -9093
rect 11390 -9127 11424 -9093
rect 11472 -9127 11506 -9093
rect 11544 -9127 11578 -9093
rect 11626 -9127 11660 -9093
rect 11698 -9127 11732 -9093
rect 11780 -9127 11814 -9093
rect 11852 -9127 11886 -9093
rect 11934 -9127 11968 -9093
rect 12006 -9127 12040 -9093
rect 4080 -9201 4114 -9167
rect 4152 -9201 4186 -9167
rect 4234 -9201 4268 -9167
rect 4306 -9201 4340 -9167
rect 4388 -9201 4422 -9167
rect 4460 -9201 4494 -9167
rect 4542 -9201 4576 -9167
rect 4614 -9201 4648 -9167
rect 4696 -9201 4730 -9167
rect 4768 -9201 4802 -9167
rect 4850 -9201 4884 -9167
rect 4922 -9201 4956 -9167
rect 5004 -9201 5038 -9167
rect 5076 -9201 5110 -9167
rect 5158 -9201 5192 -9167
rect 5230 -9201 5264 -9167
rect 5312 -9201 5346 -9167
rect 5384 -9201 5418 -9167
rect 5466 -9201 5500 -9167
rect 5538 -9201 5572 -9167
rect 5620 -9201 5654 -9167
rect 5692 -9201 5726 -9167
rect 5774 -9201 5808 -9167
rect 5846 -9201 5880 -9167
rect 5928 -9201 5962 -9167
rect 6000 -9201 6034 -9167
rect 6082 -9201 6116 -9167
rect 6154 -9201 6188 -9167
rect 6236 -9201 6270 -9167
rect 6308 -9201 6342 -9167
rect 6390 -9201 6424 -9167
rect 6462 -9201 6496 -9167
rect 6544 -9201 6578 -9167
rect 6616 -9201 6650 -9167
rect 6698 -9201 6732 -9167
rect 6770 -9201 6804 -9167
rect 6852 -9201 6886 -9167
rect 6924 -9201 6958 -9167
rect 7006 -9201 7040 -9167
rect 7078 -9201 7112 -9167
rect 7160 -9201 7194 -9167
rect 7232 -9201 7266 -9167
rect 7314 -9201 7348 -9167
rect 7386 -9201 7420 -9167
rect 7468 -9201 7502 -9167
rect 7540 -9201 7574 -9167
rect 7622 -9201 7656 -9167
rect 7694 -9201 7728 -9167
rect 7776 -9201 7810 -9167
rect 7848 -9201 7882 -9167
rect 7930 -9201 7964 -9167
rect 8002 -9201 8036 -9167
rect 8084 -9201 8118 -9167
rect 8156 -9201 8190 -9167
rect 8238 -9201 8272 -9167
rect 8310 -9201 8344 -9167
rect 8392 -9201 8426 -9167
rect 8464 -9201 8498 -9167
rect 8546 -9201 8580 -9167
rect 8618 -9201 8652 -9167
rect 8700 -9201 8734 -9167
rect 8772 -9201 8806 -9167
rect 8854 -9201 8888 -9167
rect 8926 -9201 8960 -9167
rect 9008 -9201 9042 -9167
rect 9080 -9201 9114 -9167
rect 9162 -9201 9196 -9167
rect 9234 -9201 9268 -9167
rect 9316 -9201 9350 -9167
rect 9388 -9201 9422 -9167
rect 9470 -9201 9504 -9167
rect 9542 -9201 9576 -9167
rect 9624 -9201 9658 -9167
rect 9696 -9201 9730 -9167
rect 9778 -9201 9812 -9167
rect 9850 -9201 9884 -9167
rect 9932 -9201 9966 -9167
rect 10004 -9201 10038 -9167
rect 10086 -9201 10120 -9167
rect 10158 -9201 10192 -9167
rect 10240 -9201 10274 -9167
rect 10312 -9201 10346 -9167
rect 10394 -9201 10428 -9167
rect 10466 -9201 10500 -9167
rect 10548 -9201 10582 -9167
rect 10620 -9201 10654 -9167
rect 10702 -9201 10736 -9167
rect 10774 -9201 10808 -9167
rect 10856 -9201 10890 -9167
rect 10928 -9201 10962 -9167
rect 11010 -9201 11044 -9167
rect 11082 -9201 11116 -9167
rect 11164 -9201 11198 -9167
rect 11236 -9201 11270 -9167
rect 11318 -9201 11352 -9167
rect 11390 -9201 11424 -9167
rect 11472 -9201 11506 -9167
rect 11544 -9201 11578 -9167
rect 11626 -9201 11660 -9167
rect 11698 -9201 11732 -9167
rect 11780 -9201 11814 -9167
rect 11852 -9201 11886 -9167
rect 11934 -9201 11968 -9167
rect 12006 -9201 12040 -9167
rect 12534 -9209 12568 -8333
rect 12682 -9209 12716 -8333
rect 12830 -9209 12864 -8333
rect 12978 -9209 13012 -8333
rect 13126 -9209 13160 -8333
rect 13274 -9209 13308 -8333
rect 13422 -9209 13456 -8333
rect 13570 -9209 13604 -8333
rect 13718 -9209 13752 -8333
rect 13866 -9209 13900 -8333
rect 14014 -9209 14048 -8333
rect 14162 -9209 14196 -8333
rect 14310 -9209 14344 -8333
rect 14458 -9209 14492 -8333
rect 14606 -9209 14640 -8333
rect 14754 -9209 14788 -8333
rect 14902 -9209 14936 -8333
rect 15050 -9209 15084 -8333
rect 15198 -9209 15232 -8333
rect 15346 -9209 15380 -8333
rect 15494 -9209 15528 -8333
rect 15642 -9209 15676 -8333
rect 15790 -9209 15824 -8333
rect 15938 -9209 15972 -8333
rect 16086 -9209 16120 -8333
rect 16234 -9209 16268 -8333
rect 16382 -9209 16416 -8333
rect 16530 -9209 16564 -8333
rect 16678 -9209 16712 -8333
rect 16826 -9209 16860 -8333
rect 16974 -9209 17008 -8333
rect 17122 -9209 17156 -8333
rect 17270 -9209 17304 -8333
rect 17418 -9209 17452 -8333
rect 17566 -9209 17600 -8333
rect 17714 -9209 17748 -8333
rect 17862 -9209 17896 -8333
rect 18010 -9209 18044 -8333
rect 18158 -9209 18192 -8333
rect 18306 -9209 18340 -8333
rect 18454 -9209 18488 -8333
rect 18602 -9209 18636 -8333
rect 18750 -9209 18784 -8333
rect 18898 -9209 18932 -8333
rect 19046 -9209 19080 -8333
rect 19194 -9209 19228 -8333
rect 19342 -9209 19376 -8333
rect 19490 -9209 19524 -8333
rect 19638 -9209 19672 -8333
rect 19786 -9209 19820 -8333
rect 19934 -9209 19968 -8333
rect 20082 -9209 20116 -8333
rect 20230 -9209 20264 -8333
rect 20378 -9209 20412 -8333
rect 20526 -9209 20560 -8333
rect 20674 -9209 20708 -8333
rect 20822 -9209 20856 -8333
rect 20970 -9209 21004 -8333
rect 21118 -9209 21152 -8333
rect 21266 -9209 21300 -8333
rect 21414 -9209 21448 -8333
rect 21562 -9209 21596 -8333
rect 21710 -9209 21744 -8333
rect 21858 -9209 21892 -8333
rect 22006 -9209 22040 -8333
rect 22154 -9209 22188 -8333
rect 22302 -9209 22336 -8333
rect 22450 -9209 22484 -8333
rect 22598 -9209 22632 -8333
rect 22746 -9209 22780 -8333
rect 22894 -9209 22928 -8333
rect 23042 -9209 23076 -8333
rect 23190 -9209 23224 -8333
rect 23338 -9209 23372 -8333
rect 4080 -9275 4114 -9241
rect 4152 -9275 4186 -9241
rect 4234 -9275 4268 -9241
rect 4306 -9275 4340 -9241
rect 4388 -9275 4422 -9241
rect 4460 -9275 4494 -9241
rect 4542 -9275 4576 -9241
rect 4614 -9275 4648 -9241
rect 4696 -9275 4730 -9241
rect 4768 -9275 4802 -9241
rect 4850 -9275 4884 -9241
rect 4922 -9275 4956 -9241
rect 5004 -9275 5038 -9241
rect 5076 -9275 5110 -9241
rect 5158 -9275 5192 -9241
rect 5230 -9275 5264 -9241
rect 5312 -9275 5346 -9241
rect 5384 -9275 5418 -9241
rect 5466 -9275 5500 -9241
rect 5538 -9275 5572 -9241
rect 5620 -9275 5654 -9241
rect 5692 -9275 5726 -9241
rect 5774 -9275 5808 -9241
rect 5846 -9275 5880 -9241
rect 5928 -9275 5962 -9241
rect 6000 -9275 6034 -9241
rect 6082 -9275 6116 -9241
rect 6154 -9275 6188 -9241
rect 6236 -9275 6270 -9241
rect 6308 -9275 6342 -9241
rect 6390 -9275 6424 -9241
rect 6462 -9275 6496 -9241
rect 6544 -9275 6578 -9241
rect 6616 -9275 6650 -9241
rect 6698 -9275 6732 -9241
rect 6770 -9275 6804 -9241
rect 6852 -9275 6886 -9241
rect 6924 -9275 6958 -9241
rect 7006 -9275 7040 -9241
rect 7078 -9275 7112 -9241
rect 7160 -9275 7194 -9241
rect 7232 -9275 7266 -9241
rect 7314 -9275 7348 -9241
rect 7386 -9275 7420 -9241
rect 7468 -9275 7502 -9241
rect 7540 -9275 7574 -9241
rect 7622 -9275 7656 -9241
rect 7694 -9275 7728 -9241
rect 7776 -9275 7810 -9241
rect 7848 -9275 7882 -9241
rect 7930 -9275 7964 -9241
rect 8002 -9275 8036 -9241
rect 8084 -9275 8118 -9241
rect 8156 -9275 8190 -9241
rect 8238 -9275 8272 -9241
rect 8310 -9275 8344 -9241
rect 8392 -9275 8426 -9241
rect 8464 -9275 8498 -9241
rect 8546 -9275 8580 -9241
rect 8618 -9275 8652 -9241
rect 8700 -9275 8734 -9241
rect 8772 -9275 8806 -9241
rect 8854 -9275 8888 -9241
rect 8926 -9275 8960 -9241
rect 9008 -9275 9042 -9241
rect 9080 -9275 9114 -9241
rect 9162 -9275 9196 -9241
rect 9234 -9275 9268 -9241
rect 9316 -9275 9350 -9241
rect 9388 -9275 9422 -9241
rect 9470 -9275 9504 -9241
rect 9542 -9275 9576 -9241
rect 9624 -9275 9658 -9241
rect 9696 -9275 9730 -9241
rect 9778 -9275 9812 -9241
rect 9850 -9275 9884 -9241
rect 9932 -9275 9966 -9241
rect 10004 -9275 10038 -9241
rect 10086 -9275 10120 -9241
rect 10158 -9275 10192 -9241
rect 10240 -9275 10274 -9241
rect 10312 -9275 10346 -9241
rect 10394 -9275 10428 -9241
rect 10466 -9275 10500 -9241
rect 10548 -9275 10582 -9241
rect 10620 -9275 10654 -9241
rect 10702 -9275 10736 -9241
rect 10774 -9275 10808 -9241
rect 10856 -9275 10890 -9241
rect 10928 -9275 10962 -9241
rect 11010 -9275 11044 -9241
rect 11082 -9275 11116 -9241
rect 11164 -9275 11198 -9241
rect 11236 -9275 11270 -9241
rect 11318 -9275 11352 -9241
rect 11390 -9275 11424 -9241
rect 11472 -9275 11506 -9241
rect 11544 -9275 11578 -9241
rect 11626 -9275 11660 -9241
rect 11698 -9275 11732 -9241
rect 11780 -9275 11814 -9241
rect 11852 -9275 11886 -9241
rect 11934 -9275 11968 -9241
rect 12006 -9275 12040 -9241
rect 4080 -9349 4114 -9315
rect 4152 -9349 4186 -9315
rect 4234 -9349 4268 -9315
rect 4306 -9349 4340 -9315
rect 4388 -9349 4422 -9315
rect 4460 -9349 4494 -9315
rect 4542 -9349 4576 -9315
rect 4614 -9349 4648 -9315
rect 4696 -9349 4730 -9315
rect 4768 -9349 4802 -9315
rect 4850 -9349 4884 -9315
rect 4922 -9349 4956 -9315
rect 5004 -9349 5038 -9315
rect 5076 -9349 5110 -9315
rect 5158 -9349 5192 -9315
rect 5230 -9349 5264 -9315
rect 5312 -9349 5346 -9315
rect 5384 -9349 5418 -9315
rect 5466 -9349 5500 -9315
rect 5538 -9349 5572 -9315
rect 5620 -9349 5654 -9315
rect 5692 -9349 5726 -9315
rect 5774 -9349 5808 -9315
rect 5846 -9349 5880 -9315
rect 5928 -9349 5962 -9315
rect 6000 -9349 6034 -9315
rect 6082 -9349 6116 -9315
rect 6154 -9349 6188 -9315
rect 6236 -9349 6270 -9315
rect 6308 -9349 6342 -9315
rect 6390 -9349 6424 -9315
rect 6462 -9349 6496 -9315
rect 6544 -9349 6578 -9315
rect 6616 -9349 6650 -9315
rect 6698 -9349 6732 -9315
rect 6770 -9349 6804 -9315
rect 6852 -9349 6886 -9315
rect 6924 -9349 6958 -9315
rect 7006 -9349 7040 -9315
rect 7078 -9349 7112 -9315
rect 7160 -9349 7194 -9315
rect 7232 -9349 7266 -9315
rect 7314 -9349 7348 -9315
rect 7386 -9349 7420 -9315
rect 7468 -9349 7502 -9315
rect 7540 -9349 7574 -9315
rect 7622 -9349 7656 -9315
rect 7694 -9349 7728 -9315
rect 7776 -9349 7810 -9315
rect 7848 -9349 7882 -9315
rect 7930 -9349 7964 -9315
rect 8002 -9349 8036 -9315
rect 8084 -9349 8118 -9315
rect 8156 -9349 8190 -9315
rect 8238 -9349 8272 -9315
rect 8310 -9349 8344 -9315
rect 8392 -9349 8426 -9315
rect 8464 -9349 8498 -9315
rect 8546 -9349 8580 -9315
rect 8618 -9349 8652 -9315
rect 8700 -9349 8734 -9315
rect 8772 -9349 8806 -9315
rect 8854 -9349 8888 -9315
rect 8926 -9349 8960 -9315
rect 9008 -9349 9042 -9315
rect 9080 -9349 9114 -9315
rect 9162 -9349 9196 -9315
rect 9234 -9349 9268 -9315
rect 9316 -9349 9350 -9315
rect 9388 -9349 9422 -9315
rect 9470 -9349 9504 -9315
rect 9542 -9349 9576 -9315
rect 9624 -9349 9658 -9315
rect 9696 -9349 9730 -9315
rect 9778 -9349 9812 -9315
rect 9850 -9349 9884 -9315
rect 9932 -9349 9966 -9315
rect 10004 -9349 10038 -9315
rect 10086 -9349 10120 -9315
rect 10158 -9349 10192 -9315
rect 10240 -9349 10274 -9315
rect 10312 -9349 10346 -9315
rect 10394 -9349 10428 -9315
rect 10466 -9349 10500 -9315
rect 10548 -9349 10582 -9315
rect 10620 -9349 10654 -9315
rect 10702 -9349 10736 -9315
rect 10774 -9349 10808 -9315
rect 10856 -9349 10890 -9315
rect 10928 -9349 10962 -9315
rect 11010 -9349 11044 -9315
rect 11082 -9349 11116 -9315
rect 11164 -9349 11198 -9315
rect 11236 -9349 11270 -9315
rect 11318 -9349 11352 -9315
rect 11390 -9349 11424 -9315
rect 11472 -9349 11506 -9315
rect 11544 -9349 11578 -9315
rect 11626 -9349 11660 -9315
rect 11698 -9349 11732 -9315
rect 11780 -9349 11814 -9315
rect 11852 -9349 11886 -9315
rect 11934 -9349 11968 -9315
rect 12006 -9349 12040 -9315
rect 4080 -9423 4114 -9389
rect 4152 -9423 4186 -9389
rect 4234 -9423 4268 -9389
rect 4306 -9423 4340 -9389
rect 4388 -9423 4422 -9389
rect 4460 -9423 4494 -9389
rect 4542 -9423 4576 -9389
rect 4614 -9423 4648 -9389
rect 4696 -9423 4730 -9389
rect 4768 -9423 4802 -9389
rect 4850 -9423 4884 -9389
rect 4922 -9423 4956 -9389
rect 5004 -9423 5038 -9389
rect 5076 -9423 5110 -9389
rect 5158 -9423 5192 -9389
rect 5230 -9423 5264 -9389
rect 5312 -9423 5346 -9389
rect 5384 -9423 5418 -9389
rect 5466 -9423 5500 -9389
rect 5538 -9423 5572 -9389
rect 5620 -9423 5654 -9389
rect 5692 -9423 5726 -9389
rect 5774 -9423 5808 -9389
rect 5846 -9423 5880 -9389
rect 5928 -9423 5962 -9389
rect 6000 -9423 6034 -9389
rect 6082 -9423 6116 -9389
rect 6154 -9423 6188 -9389
rect 6236 -9423 6270 -9389
rect 6308 -9423 6342 -9389
rect 6390 -9423 6424 -9389
rect 6462 -9423 6496 -9389
rect 6544 -9423 6578 -9389
rect 6616 -9423 6650 -9389
rect 6698 -9423 6732 -9389
rect 6770 -9423 6804 -9389
rect 6852 -9423 6886 -9389
rect 6924 -9423 6958 -9389
rect 7006 -9423 7040 -9389
rect 7078 -9423 7112 -9389
rect 7160 -9423 7194 -9389
rect 7232 -9423 7266 -9389
rect 7314 -9423 7348 -9389
rect 7386 -9423 7420 -9389
rect 7468 -9423 7502 -9389
rect 7540 -9423 7574 -9389
rect 7622 -9423 7656 -9389
rect 7694 -9423 7728 -9389
rect 7776 -9423 7810 -9389
rect 7848 -9423 7882 -9389
rect 7930 -9423 7964 -9389
rect 8002 -9423 8036 -9389
rect 8084 -9423 8118 -9389
rect 8156 -9423 8190 -9389
rect 8238 -9423 8272 -9389
rect 8310 -9423 8344 -9389
rect 8392 -9423 8426 -9389
rect 8464 -9423 8498 -9389
rect 8546 -9423 8580 -9389
rect 8618 -9423 8652 -9389
rect 8700 -9423 8734 -9389
rect 8772 -9423 8806 -9389
rect 8854 -9423 8888 -9389
rect 8926 -9423 8960 -9389
rect 9008 -9423 9042 -9389
rect 9080 -9423 9114 -9389
rect 9162 -9423 9196 -9389
rect 9234 -9423 9268 -9389
rect 9316 -9423 9350 -9389
rect 9388 -9423 9422 -9389
rect 9470 -9423 9504 -9389
rect 9542 -9423 9576 -9389
rect 9624 -9423 9658 -9389
rect 9696 -9423 9730 -9389
rect 9778 -9423 9812 -9389
rect 9850 -9423 9884 -9389
rect 9932 -9423 9966 -9389
rect 10004 -9423 10038 -9389
rect 10086 -9423 10120 -9389
rect 10158 -9423 10192 -9389
rect 10240 -9423 10274 -9389
rect 10312 -9423 10346 -9389
rect 10394 -9423 10428 -9389
rect 10466 -9423 10500 -9389
rect 10548 -9423 10582 -9389
rect 10620 -9423 10654 -9389
rect 10702 -9423 10736 -9389
rect 10774 -9423 10808 -9389
rect 10856 -9423 10890 -9389
rect 10928 -9423 10962 -9389
rect 11010 -9423 11044 -9389
rect 11082 -9423 11116 -9389
rect 11164 -9423 11198 -9389
rect 11236 -9423 11270 -9389
rect 11318 -9423 11352 -9389
rect 11390 -9423 11424 -9389
rect 11472 -9423 11506 -9389
rect 11544 -9423 11578 -9389
rect 11626 -9423 11660 -9389
rect 11698 -9423 11732 -9389
rect 11780 -9423 11814 -9389
rect 11852 -9423 11886 -9389
rect 11934 -9423 11968 -9389
rect 12006 -9423 12040 -9389
<< metal1 >>
rect 18489 3182 25078 3188
rect 3012 3181 25078 3182
rect 3012 3172 25079 3181
rect 3012 3120 3038 3172
rect 3090 3120 3120 3172
rect 3172 3120 3201 3172
rect 3253 3120 3282 3172
rect 3334 3120 3363 3172
rect 3415 3120 3444 3172
rect 3496 3120 3525 3172
rect 3577 3120 3606 3172
rect 3658 3120 3688 3172
rect 3740 3120 3769 3172
rect 3821 3120 3850 3172
rect 3902 3120 3931 3172
rect 3983 3120 4012 3172
rect 4064 3120 4093 3172
rect 4145 3120 4174 3172
rect 4226 3120 4256 3172
rect 4308 3120 4337 3172
rect 4389 3120 4418 3172
rect 4470 3120 4499 3172
rect 4551 3120 4580 3172
rect 4632 3120 4661 3172
rect 4713 3120 4742 3172
rect 4794 3152 4824 3172
rect 4802 3120 4824 3152
rect 4876 3120 4905 3172
rect 4957 3152 4986 3172
rect 5038 3152 5067 3172
rect 5119 3152 5148 3172
rect 5200 3152 5229 3172
rect 5281 3152 5310 3172
rect 5362 3152 5392 3172
rect 5444 3152 5473 3172
rect 4957 3120 4984 3152
rect 5038 3120 5056 3152
rect 5119 3120 5128 3152
rect 5306 3120 5310 3152
rect 5378 3120 5392 3152
rect 5450 3120 5473 3152
rect 5525 3120 5554 3172
rect 5606 3152 5635 3172
rect 5687 3152 5716 3172
rect 5768 3152 5797 3172
rect 5849 3152 5878 3172
rect 5930 3152 5960 3172
rect 6012 3152 6041 3172
rect 6093 3152 6122 3172
rect 5606 3120 5632 3152
rect 5687 3120 5704 3152
rect 5768 3120 5776 3152
rect 5954 3120 5960 3152
rect 6026 3120 6041 3152
rect 6098 3120 6122 3152
rect 6174 3120 6203 3172
rect 6255 3152 6284 3172
rect 6336 3152 6365 3172
rect 6417 3152 6446 3172
rect 6498 3152 6528 3172
rect 6580 3152 6609 3172
rect 6661 3152 6690 3172
rect 6742 3152 6771 3172
rect 6255 3120 6280 3152
rect 6336 3120 6352 3152
rect 6417 3120 6424 3152
rect 6602 3120 6609 3152
rect 6674 3120 6690 3152
rect 6746 3120 6771 3152
rect 6823 3120 6852 3172
rect 6904 3152 6933 3172
rect 6985 3152 7014 3172
rect 7066 3152 7096 3172
rect 7148 3152 7177 3172
rect 7229 3152 7258 3172
rect 7310 3152 7339 3172
rect 7391 3152 7420 3172
rect 6904 3120 6928 3152
rect 6985 3120 7000 3152
rect 7066 3120 7072 3152
rect 7250 3120 7258 3152
rect 7322 3120 7339 3152
rect 7394 3120 7420 3152
rect 7472 3120 7501 3172
rect 7553 3152 7582 3172
rect 7634 3152 7664 3172
rect 7716 3152 7745 3172
rect 7797 3152 7826 3172
rect 7878 3152 7907 3172
rect 7959 3152 7988 3172
rect 8040 3152 8069 3172
rect 7553 3120 7576 3152
rect 7634 3120 7648 3152
rect 7716 3120 7720 3152
rect 7898 3120 7907 3152
rect 7970 3120 7988 3152
rect 8042 3120 8069 3152
rect 8121 3120 8150 3172
rect 8202 3152 8232 3172
rect 8284 3152 8313 3172
rect 8365 3152 8394 3172
rect 8446 3152 8475 3172
rect 8527 3152 8556 3172
rect 8608 3152 8637 3172
rect 8689 3152 8718 3172
rect 8202 3120 8224 3152
rect 8284 3120 8296 3152
rect 8365 3120 8368 3152
rect 8474 3120 8475 3152
rect 8546 3120 8556 3152
rect 8618 3120 8637 3152
rect 8690 3120 8718 3152
rect 8770 3120 8800 3172
rect 8852 3152 8881 3172
rect 8933 3152 8962 3172
rect 9014 3152 9043 3172
rect 9095 3152 9124 3172
rect 9176 3152 9205 3172
rect 9257 3152 9286 3172
rect 8852 3120 8872 3152
rect 8933 3120 8944 3152
rect 9014 3120 9016 3152
rect 9122 3120 9124 3152
rect 9194 3120 9205 3152
rect 9266 3120 9286 3152
rect 9338 3120 9368 3172
rect 9420 3152 9449 3172
rect 9501 3152 9530 3172
rect 9582 3152 9611 3172
rect 9663 3152 9692 3172
rect 9744 3152 9773 3172
rect 9825 3152 9854 3172
rect 9906 3152 9936 3172
rect 9420 3120 9448 3152
rect 9501 3120 9520 3152
rect 9582 3120 9592 3152
rect 9663 3120 9664 3152
rect 9770 3120 9773 3152
rect 9842 3120 9854 3152
rect 9914 3120 9936 3152
rect 9988 3120 10017 3172
rect 10069 3152 10098 3172
rect 10150 3152 10179 3172
rect 10231 3152 10260 3172
rect 10312 3152 10341 3172
rect 10393 3152 10422 3172
rect 10474 3152 10504 3172
rect 10556 3152 10585 3172
rect 10069 3120 10096 3152
rect 10150 3120 10168 3152
rect 10231 3120 10240 3152
rect 10418 3120 10422 3152
rect 10490 3120 10504 3152
rect 10562 3120 10585 3152
rect 10637 3120 10666 3172
rect 10718 3152 10747 3172
rect 10718 3120 10744 3152
rect 10799 3120 10828 3172
rect 10880 3120 10909 3172
rect 10961 3120 10990 3172
rect 11042 3120 11118 3172
rect 11170 3120 11199 3172
rect 11251 3120 11280 3172
rect 11332 3120 11361 3172
rect 11413 3120 11442 3172
rect 11494 3120 11523 3172
rect 11575 3120 11604 3172
rect 11656 3120 11686 3172
rect 11738 3120 11767 3172
rect 11819 3120 11848 3172
rect 11900 3120 11929 3172
rect 11981 3120 12010 3172
rect 12062 3120 12091 3172
rect 12143 3120 12172 3172
rect 12224 3120 12254 3172
rect 12306 3120 12335 3172
rect 12387 3120 12416 3172
rect 12468 3151 12497 3172
rect 12549 3151 12578 3172
rect 12630 3151 12659 3172
rect 12492 3120 12497 3151
rect 12564 3120 12578 3151
rect 12636 3120 12659 3151
rect 12711 3120 12740 3172
rect 12792 3151 12822 3172
rect 12874 3151 12903 3172
rect 12955 3151 12984 3172
rect 13036 3151 13065 3172
rect 13117 3151 13146 3172
rect 13198 3151 13227 3172
rect 13279 3151 13308 3172
rect 12792 3120 12818 3151
rect 12874 3120 12890 3151
rect 12955 3120 12962 3151
rect 13140 3120 13146 3151
rect 13212 3120 13227 3151
rect 13284 3120 13308 3151
rect 13360 3120 13390 3172
rect 13442 3151 13471 3172
rect 13523 3151 13552 3172
rect 13604 3151 13633 3172
rect 13685 3151 13714 3172
rect 13766 3151 13795 3172
rect 13847 3151 13876 3172
rect 13928 3151 13958 3172
rect 13442 3120 13466 3151
rect 13523 3120 13538 3151
rect 13604 3120 13610 3151
rect 13788 3120 13795 3151
rect 13860 3120 13876 3151
rect 13932 3120 13958 3151
rect 14010 3120 14039 3172
rect 14091 3151 14120 3172
rect 14172 3151 14201 3172
rect 14253 3151 14282 3172
rect 14334 3151 14363 3172
rect 14415 3151 14444 3172
rect 14496 3151 14526 3172
rect 14578 3151 14607 3172
rect 14091 3120 14114 3151
rect 14172 3120 14186 3151
rect 14253 3120 14258 3151
rect 14436 3120 14444 3151
rect 14508 3120 14526 3151
rect 14580 3120 14607 3151
rect 14659 3120 14688 3172
rect 14740 3151 14769 3172
rect 14821 3151 14850 3172
rect 14902 3151 14931 3172
rect 14983 3151 15012 3172
rect 15064 3151 15094 3172
rect 15146 3151 15175 3172
rect 15227 3151 15256 3172
rect 14740 3120 14762 3151
rect 14821 3120 14834 3151
rect 14902 3120 14906 3151
rect 15084 3120 15094 3151
rect 15156 3120 15175 3151
rect 15228 3120 15256 3151
rect 15308 3120 15337 3172
rect 15389 3151 15418 3172
rect 15470 3151 15499 3172
rect 15551 3151 15580 3172
rect 15632 3151 15662 3172
rect 15714 3151 15743 3172
rect 15795 3151 15824 3172
rect 15389 3120 15410 3151
rect 15470 3120 15482 3151
rect 15551 3120 15554 3151
rect 15660 3120 15662 3151
rect 15732 3120 15743 3151
rect 15804 3120 15824 3151
rect 15876 3120 15905 3172
rect 15957 3120 15986 3172
rect 16038 3151 16067 3172
rect 16119 3151 16148 3172
rect 16200 3151 16230 3172
rect 16282 3151 16311 3172
rect 16363 3151 16392 3172
rect 16444 3151 16473 3172
rect 16038 3120 16058 3151
rect 16119 3120 16130 3151
rect 16200 3120 16202 3151
rect 16308 3120 16311 3151
rect 16380 3120 16392 3151
rect 16452 3120 16473 3151
rect 16525 3120 16554 3172
rect 16606 3151 16635 3172
rect 16687 3151 16716 3172
rect 16768 3151 16798 3172
rect 16850 3151 16879 3172
rect 16931 3151 16960 3172
rect 17012 3151 17041 3172
rect 17093 3151 17122 3172
rect 16606 3120 16634 3151
rect 16687 3120 16706 3151
rect 16768 3120 16778 3151
rect 16956 3120 16960 3151
rect 17028 3120 17041 3151
rect 17100 3120 17122 3151
rect 17174 3120 17203 3172
rect 17255 3151 17284 3172
rect 17336 3151 17366 3172
rect 17418 3151 17447 3172
rect 17499 3151 17528 3172
rect 17580 3151 17609 3172
rect 17661 3151 17690 3172
rect 17742 3151 17771 3172
rect 17255 3120 17282 3151
rect 17336 3120 17354 3151
rect 17418 3120 17426 3151
rect 17604 3120 17609 3151
rect 17676 3120 17690 3151
rect 17748 3120 17771 3151
rect 17823 3120 17852 3172
rect 17904 3151 17934 3172
rect 17986 3151 18015 3172
rect 18067 3151 18096 3172
rect 18148 3151 18177 3172
rect 18229 3151 18258 3172
rect 18310 3151 18339 3172
rect 18391 3151 18420 3172
rect 17904 3120 17930 3151
rect 17986 3120 18002 3151
rect 18067 3120 18074 3151
rect 18252 3120 18258 3151
rect 18324 3120 18339 3151
rect 18396 3120 18420 3151
rect 18472 3120 18502 3172
rect 18554 3120 18583 3172
rect 18635 3120 18664 3172
rect 18716 3151 18745 3172
rect 18797 3151 18826 3172
rect 18878 3151 18907 3172
rect 18959 3151 18988 3172
rect 19040 3151 19070 3172
rect 19122 3151 19151 3172
rect 19203 3151 19232 3172
rect 18716 3120 18741 3151
rect 18797 3120 18813 3151
rect 18878 3120 18885 3151
rect 19063 3120 19070 3151
rect 19135 3120 19151 3151
rect 19207 3120 19232 3151
rect 19284 3120 19313 3172
rect 19365 3151 19394 3172
rect 19446 3151 19475 3172
rect 19527 3151 19556 3172
rect 19608 3151 19638 3172
rect 19690 3151 19719 3172
rect 19771 3151 19800 3172
rect 19852 3151 19881 3172
rect 19365 3120 19389 3151
rect 19446 3120 19461 3151
rect 19527 3120 19533 3151
rect 19711 3120 19719 3151
rect 19783 3120 19800 3151
rect 19855 3120 19881 3151
rect 19933 3120 19962 3172
rect 20014 3151 20043 3172
rect 20095 3151 20124 3172
rect 20176 3151 20206 3172
rect 20258 3151 20287 3172
rect 20339 3151 20368 3172
rect 20420 3151 20449 3172
rect 20501 3151 20530 3172
rect 20014 3120 20037 3151
rect 20095 3120 20109 3151
rect 20176 3120 20181 3151
rect 20359 3120 20368 3151
rect 20431 3120 20449 3151
rect 20503 3120 20530 3151
rect 20582 3120 20611 3172
rect 20663 3151 20692 3172
rect 20744 3151 20774 3172
rect 20826 3151 20855 3172
rect 20907 3151 20936 3172
rect 20988 3151 21017 3172
rect 21069 3151 21098 3172
rect 21150 3151 21179 3172
rect 20663 3120 20685 3151
rect 20744 3120 20757 3151
rect 20826 3120 20829 3151
rect 20935 3120 20936 3151
rect 21007 3120 21017 3151
rect 21079 3120 21098 3151
rect 21151 3120 21179 3151
rect 21231 3120 21260 3172
rect 21312 3151 21342 3172
rect 21394 3151 21423 3172
rect 21475 3151 21504 3172
rect 21556 3151 21585 3172
rect 21637 3151 21666 3172
rect 21718 3151 21747 3172
rect 21312 3120 21333 3151
rect 21394 3120 21405 3151
rect 21475 3120 21477 3151
rect 21583 3120 21585 3151
rect 21655 3120 21666 3151
rect 21727 3120 21747 3151
rect 21799 3120 21828 3172
rect 21880 3151 21910 3172
rect 21962 3151 21991 3172
rect 22043 3151 22072 3172
rect 22124 3151 22153 3172
rect 22205 3151 22234 3172
rect 22286 3151 22315 3172
rect 22367 3151 22396 3172
rect 21880 3120 21909 3151
rect 21962 3120 21981 3151
rect 22043 3120 22053 3151
rect 22124 3120 22125 3151
rect 22231 3120 22234 3151
rect 22303 3120 22315 3151
rect 22375 3120 22396 3151
rect 22448 3120 22478 3172
rect 22530 3151 22559 3172
rect 22611 3151 22640 3172
rect 22692 3151 22721 3172
rect 22773 3151 22802 3172
rect 22854 3151 22883 3172
rect 22935 3151 22964 3172
rect 23016 3151 23046 3172
rect 22530 3120 22557 3151
rect 22611 3120 22629 3151
rect 22692 3120 22701 3151
rect 22879 3120 22883 3151
rect 22951 3120 22964 3151
rect 23023 3120 23046 3151
rect 23098 3120 23127 3172
rect 23179 3151 23208 3172
rect 23260 3151 23289 3172
rect 23341 3151 23370 3172
rect 23422 3151 23451 3172
rect 23503 3151 23532 3172
rect 23584 3151 23614 3172
rect 23666 3151 23695 3172
rect 23179 3120 23205 3151
rect 23260 3120 23277 3151
rect 23341 3120 23349 3151
rect 23527 3120 23532 3151
rect 23599 3120 23614 3151
rect 23671 3120 23695 3151
rect 23747 3120 23776 3172
rect 23828 3151 23857 3172
rect 23909 3151 23938 3172
rect 23990 3151 24019 3172
rect 24071 3151 24100 3172
rect 24152 3151 24182 3172
rect 24234 3151 24263 3172
rect 24315 3151 24344 3172
rect 23828 3120 23853 3151
rect 23909 3120 23925 3151
rect 23990 3120 23997 3151
rect 24175 3120 24182 3151
rect 24247 3120 24263 3151
rect 24319 3120 24344 3151
rect 24396 3120 24425 3172
rect 24477 3151 24506 3172
rect 24558 3151 24587 3172
rect 24477 3120 24501 3151
rect 24558 3120 24573 3151
rect 24639 3120 24668 3172
rect 24720 3120 25079 3172
rect 3012 3118 4768 3120
rect 4802 3118 4840 3120
rect 4874 3118 4912 3120
rect 4946 3118 4984 3120
rect 5018 3118 5056 3120
rect 5090 3118 5128 3120
rect 5162 3118 5200 3120
rect 5234 3118 5272 3120
rect 5306 3118 5344 3120
rect 5378 3118 5416 3120
rect 5450 3118 5488 3120
rect 5522 3118 5560 3120
rect 5594 3118 5632 3120
rect 5666 3118 5704 3120
rect 5738 3118 5776 3120
rect 5810 3118 5848 3120
rect 5882 3118 5920 3120
rect 5954 3118 5992 3120
rect 6026 3118 6064 3120
rect 6098 3118 6136 3120
rect 6170 3118 6208 3120
rect 6242 3118 6280 3120
rect 6314 3118 6352 3120
rect 6386 3118 6424 3120
rect 6458 3118 6496 3120
rect 6530 3118 6568 3120
rect 6602 3118 6640 3120
rect 6674 3118 6712 3120
rect 6746 3118 6784 3120
rect 6818 3118 6856 3120
rect 6890 3118 6928 3120
rect 6962 3118 7000 3120
rect 7034 3118 7072 3120
rect 7106 3118 7144 3120
rect 7178 3118 7216 3120
rect 7250 3118 7288 3120
rect 7322 3118 7360 3120
rect 7394 3118 7432 3120
rect 7466 3118 7504 3120
rect 7538 3118 7576 3120
rect 7610 3118 7648 3120
rect 7682 3118 7720 3120
rect 7754 3118 7792 3120
rect 7826 3118 7864 3120
rect 7898 3118 7936 3120
rect 7970 3118 8008 3120
rect 8042 3118 8080 3120
rect 8114 3118 8152 3120
rect 8186 3118 8224 3120
rect 8258 3118 8296 3120
rect 8330 3118 8368 3120
rect 8402 3118 8440 3120
rect 8474 3118 8512 3120
rect 8546 3118 8584 3120
rect 8618 3118 8656 3120
rect 8690 3118 8728 3120
rect 8762 3118 8800 3120
rect 8834 3118 8872 3120
rect 8906 3118 8944 3120
rect 8978 3118 9016 3120
rect 9050 3118 9088 3120
rect 9122 3118 9160 3120
rect 9194 3118 9232 3120
rect 9266 3118 9304 3120
rect 9338 3118 9376 3120
rect 9410 3118 9448 3120
rect 9482 3118 9520 3120
rect 9554 3118 9592 3120
rect 9626 3118 9664 3120
rect 9698 3118 9736 3120
rect 9770 3118 9808 3120
rect 9842 3118 9880 3120
rect 9914 3118 9952 3120
rect 9986 3118 10024 3120
rect 10058 3118 10096 3120
rect 10130 3118 10168 3120
rect 10202 3118 10240 3120
rect 10274 3118 10312 3120
rect 10346 3118 10384 3120
rect 10418 3118 10456 3120
rect 10490 3118 10528 3120
rect 10562 3118 10600 3120
rect 10634 3118 10672 3120
rect 10706 3118 10744 3120
rect 10778 3118 12458 3120
rect 3012 3117 12458 3118
rect 12492 3117 12530 3120
rect 12564 3117 12602 3120
rect 12636 3117 12674 3120
rect 12708 3117 12746 3120
rect 12780 3117 12818 3120
rect 12852 3117 12890 3120
rect 12924 3117 12962 3120
rect 12996 3117 13034 3120
rect 13068 3117 13106 3120
rect 13140 3117 13178 3120
rect 13212 3117 13250 3120
rect 13284 3117 13322 3120
rect 13356 3117 13394 3120
rect 13428 3117 13466 3120
rect 13500 3117 13538 3120
rect 13572 3117 13610 3120
rect 13644 3117 13682 3120
rect 13716 3117 13754 3120
rect 13788 3117 13826 3120
rect 13860 3117 13898 3120
rect 13932 3117 13970 3120
rect 14004 3117 14042 3120
rect 14076 3117 14114 3120
rect 14148 3117 14186 3120
rect 14220 3117 14258 3120
rect 14292 3117 14330 3120
rect 14364 3117 14402 3120
rect 14436 3117 14474 3120
rect 14508 3117 14546 3120
rect 14580 3117 14618 3120
rect 14652 3117 14690 3120
rect 14724 3117 14762 3120
rect 14796 3117 14834 3120
rect 14868 3117 14906 3120
rect 14940 3117 14978 3120
rect 15012 3117 15050 3120
rect 15084 3117 15122 3120
rect 15156 3117 15194 3120
rect 15228 3117 15266 3120
rect 15300 3117 15338 3120
rect 15372 3117 15410 3120
rect 15444 3117 15482 3120
rect 15516 3117 15554 3120
rect 15588 3117 15626 3120
rect 15660 3117 15698 3120
rect 15732 3117 15770 3120
rect 15804 3117 15842 3120
rect 15876 3117 15914 3120
rect 15948 3117 15986 3120
rect 16020 3117 16058 3120
rect 16092 3117 16130 3120
rect 16164 3117 16202 3120
rect 16236 3117 16274 3120
rect 16308 3117 16346 3120
rect 16380 3117 16418 3120
rect 16452 3117 16490 3120
rect 16524 3117 16562 3120
rect 16596 3117 16634 3120
rect 16668 3117 16706 3120
rect 16740 3117 16778 3120
rect 16812 3117 16850 3120
rect 16884 3117 16922 3120
rect 16956 3117 16994 3120
rect 17028 3117 17066 3120
rect 17100 3117 17138 3120
rect 17172 3117 17210 3120
rect 17244 3117 17282 3120
rect 17316 3117 17354 3120
rect 17388 3117 17426 3120
rect 17460 3117 17498 3120
rect 17532 3117 17570 3120
rect 17604 3117 17642 3120
rect 17676 3117 17714 3120
rect 17748 3117 17786 3120
rect 17820 3117 17858 3120
rect 17892 3117 17930 3120
rect 17964 3117 18002 3120
rect 18036 3117 18074 3120
rect 18108 3117 18146 3120
rect 18180 3117 18218 3120
rect 18252 3117 18290 3120
rect 18324 3117 18362 3120
rect 18396 3117 18434 3120
rect 18468 3117 18597 3120
rect 18631 3117 18669 3120
rect 18703 3117 18741 3120
rect 18775 3117 18813 3120
rect 18847 3117 18885 3120
rect 18919 3117 18957 3120
rect 18991 3117 19029 3120
rect 19063 3117 19101 3120
rect 19135 3117 19173 3120
rect 19207 3117 19245 3120
rect 19279 3117 19317 3120
rect 19351 3117 19389 3120
rect 19423 3117 19461 3120
rect 19495 3117 19533 3120
rect 19567 3117 19605 3120
rect 19639 3117 19677 3120
rect 19711 3117 19749 3120
rect 19783 3117 19821 3120
rect 19855 3117 19893 3120
rect 19927 3117 19965 3120
rect 19999 3117 20037 3120
rect 20071 3117 20109 3120
rect 20143 3117 20181 3120
rect 20215 3117 20253 3120
rect 20287 3117 20325 3120
rect 20359 3117 20397 3120
rect 20431 3117 20469 3120
rect 20503 3117 20541 3120
rect 20575 3117 20613 3120
rect 20647 3117 20685 3120
rect 20719 3117 20757 3120
rect 20791 3117 20829 3120
rect 20863 3117 20901 3120
rect 20935 3117 20973 3120
rect 21007 3117 21045 3120
rect 21079 3117 21117 3120
rect 21151 3117 21189 3120
rect 21223 3117 21261 3120
rect 21295 3117 21333 3120
rect 21367 3117 21405 3120
rect 21439 3117 21477 3120
rect 21511 3117 21549 3120
rect 21583 3117 21621 3120
rect 21655 3117 21693 3120
rect 21727 3117 21765 3120
rect 21799 3117 21837 3120
rect 21871 3117 21909 3120
rect 21943 3117 21981 3120
rect 22015 3117 22053 3120
rect 22087 3117 22125 3120
rect 22159 3117 22197 3120
rect 22231 3117 22269 3120
rect 22303 3117 22341 3120
rect 22375 3117 22413 3120
rect 22447 3117 22485 3120
rect 22519 3117 22557 3120
rect 22591 3117 22629 3120
rect 22663 3117 22701 3120
rect 22735 3117 22773 3120
rect 22807 3117 22845 3120
rect 22879 3117 22917 3120
rect 22951 3117 22989 3120
rect 23023 3117 23061 3120
rect 23095 3117 23133 3120
rect 23167 3117 23205 3120
rect 23239 3117 23277 3120
rect 23311 3117 23349 3120
rect 23383 3117 23421 3120
rect 23455 3117 23493 3120
rect 23527 3117 23565 3120
rect 23599 3117 23637 3120
rect 23671 3117 23709 3120
rect 23743 3117 23781 3120
rect 23815 3117 23853 3120
rect 23887 3117 23925 3120
rect 23959 3117 23997 3120
rect 24031 3117 24069 3120
rect 24103 3117 24141 3120
rect 24175 3117 24213 3120
rect 24247 3117 24285 3120
rect 24319 3117 24357 3120
rect 24391 3117 24429 3120
rect 24463 3117 24501 3120
rect 24535 3117 24573 3120
rect 24607 3117 25079 3120
rect 3012 3068 25079 3117
rect 3012 3016 3038 3068
rect 3090 3016 3120 3068
rect 3172 3016 3201 3068
rect 3253 3016 3282 3068
rect 3334 3016 3363 3068
rect 3415 3016 3444 3068
rect 3496 3016 3525 3068
rect 3577 3016 3606 3068
rect 3658 3016 3688 3068
rect 3740 3016 3769 3068
rect 3821 3016 3850 3068
rect 3902 3016 3931 3068
rect 3983 3016 4012 3068
rect 4064 3016 4093 3068
rect 4145 3016 4174 3068
rect 4226 3016 4256 3068
rect 4308 3016 4337 3068
rect 4389 3016 4418 3068
rect 4470 3016 4499 3068
rect 4551 3016 4580 3068
rect 4632 3016 4661 3068
rect 4713 3016 4742 3068
rect 4794 3064 4824 3068
rect 4802 3030 4824 3064
rect 4794 3016 4824 3030
rect 4876 3016 4905 3068
rect 4957 3064 4986 3068
rect 5038 3064 5067 3068
rect 5119 3064 5148 3068
rect 5200 3064 5229 3068
rect 5281 3064 5310 3068
rect 5362 3064 5392 3068
rect 5444 3064 5473 3068
rect 4957 3030 4984 3064
rect 5038 3030 5056 3064
rect 5119 3030 5128 3064
rect 5306 3030 5310 3064
rect 5378 3030 5392 3064
rect 5450 3030 5473 3064
rect 4957 3016 4986 3030
rect 5038 3016 5067 3030
rect 5119 3016 5148 3030
rect 5200 3016 5229 3030
rect 5281 3016 5310 3030
rect 5362 3016 5392 3030
rect 5444 3016 5473 3030
rect 5525 3016 5554 3068
rect 5606 3064 5635 3068
rect 5687 3064 5716 3068
rect 5768 3064 5797 3068
rect 5849 3064 5878 3068
rect 5930 3064 5960 3068
rect 6012 3064 6041 3068
rect 6093 3064 6122 3068
rect 5606 3030 5632 3064
rect 5687 3030 5704 3064
rect 5768 3030 5776 3064
rect 5954 3030 5960 3064
rect 6026 3030 6041 3064
rect 6098 3030 6122 3064
rect 5606 3016 5635 3030
rect 5687 3016 5716 3030
rect 5768 3016 5797 3030
rect 5849 3016 5878 3030
rect 5930 3016 5960 3030
rect 6012 3016 6041 3030
rect 6093 3016 6122 3030
rect 6174 3016 6203 3068
rect 6255 3064 6284 3068
rect 6336 3064 6365 3068
rect 6417 3064 6446 3068
rect 6498 3064 6528 3068
rect 6580 3064 6609 3068
rect 6661 3064 6690 3068
rect 6742 3064 6771 3068
rect 6255 3030 6280 3064
rect 6336 3030 6352 3064
rect 6417 3030 6424 3064
rect 6602 3030 6609 3064
rect 6674 3030 6690 3064
rect 6746 3030 6771 3064
rect 6255 3016 6284 3030
rect 6336 3016 6365 3030
rect 6417 3016 6446 3030
rect 6498 3016 6528 3030
rect 6580 3016 6609 3030
rect 6661 3016 6690 3030
rect 6742 3016 6771 3030
rect 6823 3016 6852 3068
rect 6904 3064 6933 3068
rect 6985 3064 7014 3068
rect 7066 3064 7096 3068
rect 7148 3064 7177 3068
rect 7229 3064 7258 3068
rect 7310 3064 7339 3068
rect 7391 3064 7420 3068
rect 6904 3030 6928 3064
rect 6985 3030 7000 3064
rect 7066 3030 7072 3064
rect 7250 3030 7258 3064
rect 7322 3030 7339 3064
rect 7394 3030 7420 3064
rect 6904 3016 6933 3030
rect 6985 3016 7014 3030
rect 7066 3016 7096 3030
rect 7148 3016 7177 3030
rect 7229 3016 7258 3030
rect 7310 3016 7339 3030
rect 7391 3016 7420 3030
rect 7472 3016 7501 3068
rect 7553 3064 7582 3068
rect 7634 3064 7664 3068
rect 7716 3064 7745 3068
rect 7797 3064 7826 3068
rect 7878 3064 7907 3068
rect 7959 3064 7988 3068
rect 8040 3064 8069 3068
rect 7553 3030 7576 3064
rect 7634 3030 7648 3064
rect 7716 3030 7720 3064
rect 7898 3030 7907 3064
rect 7970 3030 7988 3064
rect 8042 3030 8069 3064
rect 7553 3016 7582 3030
rect 7634 3016 7664 3030
rect 7716 3016 7745 3030
rect 7797 3016 7826 3030
rect 7878 3016 7907 3030
rect 7959 3016 7988 3030
rect 8040 3016 8069 3030
rect 8121 3016 8150 3068
rect 8202 3064 8232 3068
rect 8284 3064 8313 3068
rect 8365 3064 8394 3068
rect 8446 3064 8475 3068
rect 8527 3064 8556 3068
rect 8608 3064 8637 3068
rect 8689 3064 8718 3068
rect 8202 3030 8224 3064
rect 8284 3030 8296 3064
rect 8365 3030 8368 3064
rect 8474 3030 8475 3064
rect 8546 3030 8556 3064
rect 8618 3030 8637 3064
rect 8690 3030 8718 3064
rect 8202 3016 8232 3030
rect 8284 3016 8313 3030
rect 8365 3016 8394 3030
rect 8446 3016 8475 3030
rect 8527 3016 8556 3030
rect 8608 3016 8637 3030
rect 8689 3016 8718 3030
rect 8770 3016 8800 3068
rect 8852 3064 8881 3068
rect 8933 3064 8962 3068
rect 9014 3064 9043 3068
rect 9095 3064 9124 3068
rect 9176 3064 9205 3068
rect 9257 3064 9286 3068
rect 8852 3030 8872 3064
rect 8933 3030 8944 3064
rect 9014 3030 9016 3064
rect 9122 3030 9124 3064
rect 9194 3030 9205 3064
rect 9266 3030 9286 3064
rect 8852 3016 8881 3030
rect 8933 3016 8962 3030
rect 9014 3016 9043 3030
rect 9095 3016 9124 3030
rect 9176 3016 9205 3030
rect 9257 3016 9286 3030
rect 9338 3016 9368 3068
rect 9420 3064 9449 3068
rect 9501 3064 9530 3068
rect 9582 3064 9611 3068
rect 9663 3064 9692 3068
rect 9744 3064 9773 3068
rect 9825 3064 9854 3068
rect 9906 3064 9936 3068
rect 9420 3030 9448 3064
rect 9501 3030 9520 3064
rect 9582 3030 9592 3064
rect 9663 3030 9664 3064
rect 9770 3030 9773 3064
rect 9842 3030 9854 3064
rect 9914 3030 9936 3064
rect 9420 3016 9449 3030
rect 9501 3016 9530 3030
rect 9582 3016 9611 3030
rect 9663 3016 9692 3030
rect 9744 3016 9773 3030
rect 9825 3016 9854 3030
rect 9906 3016 9936 3030
rect 9988 3016 10017 3068
rect 10069 3064 10098 3068
rect 10150 3064 10179 3068
rect 10231 3064 10260 3068
rect 10312 3064 10341 3068
rect 10393 3064 10422 3068
rect 10474 3064 10504 3068
rect 10556 3064 10585 3068
rect 10069 3030 10096 3064
rect 10150 3030 10168 3064
rect 10231 3030 10240 3064
rect 10418 3030 10422 3064
rect 10490 3030 10504 3064
rect 10562 3030 10585 3064
rect 10069 3016 10098 3030
rect 10150 3016 10179 3030
rect 10231 3016 10260 3030
rect 10312 3016 10341 3030
rect 10393 3016 10422 3030
rect 10474 3016 10504 3030
rect 10556 3016 10585 3030
rect 10637 3016 10666 3068
rect 10718 3064 10747 3068
rect 10718 3030 10744 3064
rect 10718 3016 10747 3030
rect 10799 3016 10828 3068
rect 10880 3016 10909 3068
rect 10961 3016 10990 3068
rect 11042 3016 11118 3068
rect 11170 3016 11199 3068
rect 11251 3016 11280 3068
rect 11332 3016 11361 3068
rect 11413 3016 11442 3068
rect 11494 3016 11523 3068
rect 11575 3016 11604 3068
rect 11656 3016 11686 3068
rect 11738 3016 11767 3068
rect 11819 3016 11848 3068
rect 11900 3016 11929 3068
rect 11981 3016 12010 3068
rect 12062 3016 12091 3068
rect 12143 3016 12172 3068
rect 12224 3016 12254 3068
rect 12306 3016 12335 3068
rect 12387 3016 12416 3068
rect 12468 3063 12497 3068
rect 12549 3063 12578 3068
rect 12630 3063 12659 3068
rect 12492 3029 12497 3063
rect 12564 3029 12578 3063
rect 12636 3029 12659 3063
rect 12468 3016 12497 3029
rect 12549 3016 12578 3029
rect 12630 3016 12659 3029
rect 12711 3016 12740 3068
rect 12792 3063 12822 3068
rect 12874 3063 12903 3068
rect 12955 3063 12984 3068
rect 13036 3063 13065 3068
rect 13117 3063 13146 3068
rect 13198 3063 13227 3068
rect 13279 3063 13308 3068
rect 12792 3029 12818 3063
rect 12874 3029 12890 3063
rect 12955 3029 12962 3063
rect 13140 3029 13146 3063
rect 13212 3029 13227 3063
rect 13284 3029 13308 3063
rect 12792 3016 12822 3029
rect 12874 3016 12903 3029
rect 12955 3016 12984 3029
rect 13036 3016 13065 3029
rect 13117 3016 13146 3029
rect 13198 3016 13227 3029
rect 13279 3016 13308 3029
rect 13360 3016 13390 3068
rect 13442 3063 13471 3068
rect 13523 3063 13552 3068
rect 13604 3063 13633 3068
rect 13685 3063 13714 3068
rect 13766 3063 13795 3068
rect 13847 3063 13876 3068
rect 13928 3063 13958 3068
rect 13442 3029 13466 3063
rect 13523 3029 13538 3063
rect 13604 3029 13610 3063
rect 13788 3029 13795 3063
rect 13860 3029 13876 3063
rect 13932 3029 13958 3063
rect 13442 3016 13471 3029
rect 13523 3016 13552 3029
rect 13604 3016 13633 3029
rect 13685 3016 13714 3029
rect 13766 3016 13795 3029
rect 13847 3016 13876 3029
rect 13928 3016 13958 3029
rect 14010 3016 14039 3068
rect 14091 3063 14120 3068
rect 14172 3063 14201 3068
rect 14253 3063 14282 3068
rect 14334 3063 14363 3068
rect 14415 3063 14444 3068
rect 14496 3063 14526 3068
rect 14578 3063 14607 3068
rect 14091 3029 14114 3063
rect 14172 3029 14186 3063
rect 14253 3029 14258 3063
rect 14436 3029 14444 3063
rect 14508 3029 14526 3063
rect 14580 3029 14607 3063
rect 14091 3016 14120 3029
rect 14172 3016 14201 3029
rect 14253 3016 14282 3029
rect 14334 3016 14363 3029
rect 14415 3016 14444 3029
rect 14496 3016 14526 3029
rect 14578 3016 14607 3029
rect 14659 3016 14688 3068
rect 14740 3063 14769 3068
rect 14821 3063 14850 3068
rect 14902 3063 14931 3068
rect 14983 3063 15012 3068
rect 15064 3063 15094 3068
rect 15146 3063 15175 3068
rect 15227 3063 15256 3068
rect 14740 3029 14762 3063
rect 14821 3029 14834 3063
rect 14902 3029 14906 3063
rect 15084 3029 15094 3063
rect 15156 3029 15175 3063
rect 15228 3029 15256 3063
rect 14740 3016 14769 3029
rect 14821 3016 14850 3029
rect 14902 3016 14931 3029
rect 14983 3016 15012 3029
rect 15064 3016 15094 3029
rect 15146 3016 15175 3029
rect 15227 3016 15256 3029
rect 15308 3016 15337 3068
rect 15389 3063 15418 3068
rect 15470 3063 15499 3068
rect 15551 3063 15580 3068
rect 15632 3063 15662 3068
rect 15714 3063 15743 3068
rect 15795 3063 15824 3068
rect 15389 3029 15410 3063
rect 15470 3029 15482 3063
rect 15551 3029 15554 3063
rect 15660 3029 15662 3063
rect 15732 3029 15743 3063
rect 15804 3029 15824 3063
rect 15389 3016 15418 3029
rect 15470 3016 15499 3029
rect 15551 3016 15580 3029
rect 15632 3016 15662 3029
rect 15714 3016 15743 3029
rect 15795 3016 15824 3029
rect 15876 3016 15905 3068
rect 15957 3016 15986 3068
rect 16038 3063 16067 3068
rect 16119 3063 16148 3068
rect 16200 3063 16230 3068
rect 16282 3063 16311 3068
rect 16363 3063 16392 3068
rect 16444 3063 16473 3068
rect 16038 3029 16058 3063
rect 16119 3029 16130 3063
rect 16200 3029 16202 3063
rect 16308 3029 16311 3063
rect 16380 3029 16392 3063
rect 16452 3029 16473 3063
rect 16038 3016 16067 3029
rect 16119 3016 16148 3029
rect 16200 3016 16230 3029
rect 16282 3016 16311 3029
rect 16363 3016 16392 3029
rect 16444 3016 16473 3029
rect 16525 3016 16554 3068
rect 16606 3063 16635 3068
rect 16687 3063 16716 3068
rect 16768 3063 16798 3068
rect 16850 3063 16879 3068
rect 16931 3063 16960 3068
rect 17012 3063 17041 3068
rect 17093 3063 17122 3068
rect 16606 3029 16634 3063
rect 16687 3029 16706 3063
rect 16768 3029 16778 3063
rect 16956 3029 16960 3063
rect 17028 3029 17041 3063
rect 17100 3029 17122 3063
rect 16606 3016 16635 3029
rect 16687 3016 16716 3029
rect 16768 3016 16798 3029
rect 16850 3016 16879 3029
rect 16931 3016 16960 3029
rect 17012 3016 17041 3029
rect 17093 3016 17122 3029
rect 17174 3016 17203 3068
rect 17255 3063 17284 3068
rect 17336 3063 17366 3068
rect 17418 3063 17447 3068
rect 17499 3063 17528 3068
rect 17580 3063 17609 3068
rect 17661 3063 17690 3068
rect 17742 3063 17771 3068
rect 17255 3029 17282 3063
rect 17336 3029 17354 3063
rect 17418 3029 17426 3063
rect 17604 3029 17609 3063
rect 17676 3029 17690 3063
rect 17748 3029 17771 3063
rect 17255 3016 17284 3029
rect 17336 3016 17366 3029
rect 17418 3016 17447 3029
rect 17499 3016 17528 3029
rect 17580 3016 17609 3029
rect 17661 3016 17690 3029
rect 17742 3016 17771 3029
rect 17823 3016 17852 3068
rect 17904 3063 17934 3068
rect 17986 3063 18015 3068
rect 18067 3063 18096 3068
rect 18148 3063 18177 3068
rect 18229 3063 18258 3068
rect 18310 3063 18339 3068
rect 18391 3063 18420 3068
rect 17904 3029 17930 3063
rect 17986 3029 18002 3063
rect 18067 3029 18074 3063
rect 18252 3029 18258 3063
rect 18324 3029 18339 3063
rect 18396 3029 18420 3063
rect 17904 3016 17934 3029
rect 17986 3016 18015 3029
rect 18067 3016 18096 3029
rect 18148 3016 18177 3029
rect 18229 3016 18258 3029
rect 18310 3016 18339 3029
rect 18391 3016 18420 3029
rect 18472 3016 18502 3068
rect 18554 3016 18583 3068
rect 18635 3016 18664 3068
rect 18716 3063 18745 3068
rect 18797 3063 18826 3068
rect 18878 3063 18907 3068
rect 18959 3063 18988 3068
rect 19040 3063 19070 3068
rect 19122 3063 19151 3068
rect 19203 3063 19232 3068
rect 18716 3029 18741 3063
rect 18797 3029 18813 3063
rect 18878 3029 18885 3063
rect 19063 3029 19070 3063
rect 19135 3029 19151 3063
rect 19207 3029 19232 3063
rect 18716 3016 18745 3029
rect 18797 3016 18826 3029
rect 18878 3016 18907 3029
rect 18959 3016 18988 3029
rect 19040 3016 19070 3029
rect 19122 3016 19151 3029
rect 19203 3016 19232 3029
rect 19284 3016 19313 3068
rect 19365 3063 19394 3068
rect 19446 3063 19475 3068
rect 19527 3063 19556 3068
rect 19608 3063 19638 3068
rect 19690 3063 19719 3068
rect 19771 3063 19800 3068
rect 19852 3063 19881 3068
rect 19365 3029 19389 3063
rect 19446 3029 19461 3063
rect 19527 3029 19533 3063
rect 19711 3029 19719 3063
rect 19783 3029 19800 3063
rect 19855 3029 19881 3063
rect 19365 3016 19394 3029
rect 19446 3016 19475 3029
rect 19527 3016 19556 3029
rect 19608 3016 19638 3029
rect 19690 3016 19719 3029
rect 19771 3016 19800 3029
rect 19852 3016 19881 3029
rect 19933 3016 19962 3068
rect 20014 3063 20043 3068
rect 20095 3063 20124 3068
rect 20176 3063 20206 3068
rect 20258 3063 20287 3068
rect 20339 3063 20368 3068
rect 20420 3063 20449 3068
rect 20501 3063 20530 3068
rect 20014 3029 20037 3063
rect 20095 3029 20109 3063
rect 20176 3029 20181 3063
rect 20359 3029 20368 3063
rect 20431 3029 20449 3063
rect 20503 3029 20530 3063
rect 20014 3016 20043 3029
rect 20095 3016 20124 3029
rect 20176 3016 20206 3029
rect 20258 3016 20287 3029
rect 20339 3016 20368 3029
rect 20420 3016 20449 3029
rect 20501 3016 20530 3029
rect 20582 3016 20611 3068
rect 20663 3063 20692 3068
rect 20744 3063 20774 3068
rect 20826 3063 20855 3068
rect 20907 3063 20936 3068
rect 20988 3063 21017 3068
rect 21069 3063 21098 3068
rect 21150 3063 21179 3068
rect 20663 3029 20685 3063
rect 20744 3029 20757 3063
rect 20826 3029 20829 3063
rect 20935 3029 20936 3063
rect 21007 3029 21017 3063
rect 21079 3029 21098 3063
rect 21151 3029 21179 3063
rect 20663 3016 20692 3029
rect 20744 3016 20774 3029
rect 20826 3016 20855 3029
rect 20907 3016 20936 3029
rect 20988 3016 21017 3029
rect 21069 3016 21098 3029
rect 21150 3016 21179 3029
rect 21231 3016 21260 3068
rect 21312 3063 21342 3068
rect 21394 3063 21423 3068
rect 21475 3063 21504 3068
rect 21556 3063 21585 3068
rect 21637 3063 21666 3068
rect 21718 3063 21747 3068
rect 21312 3029 21333 3063
rect 21394 3029 21405 3063
rect 21475 3029 21477 3063
rect 21583 3029 21585 3063
rect 21655 3029 21666 3063
rect 21727 3029 21747 3063
rect 21312 3016 21342 3029
rect 21394 3016 21423 3029
rect 21475 3016 21504 3029
rect 21556 3016 21585 3029
rect 21637 3016 21666 3029
rect 21718 3016 21747 3029
rect 21799 3016 21828 3068
rect 21880 3063 21910 3068
rect 21962 3063 21991 3068
rect 22043 3063 22072 3068
rect 22124 3063 22153 3068
rect 22205 3063 22234 3068
rect 22286 3063 22315 3068
rect 22367 3063 22396 3068
rect 21880 3029 21909 3063
rect 21962 3029 21981 3063
rect 22043 3029 22053 3063
rect 22124 3029 22125 3063
rect 22231 3029 22234 3063
rect 22303 3029 22315 3063
rect 22375 3029 22396 3063
rect 21880 3016 21910 3029
rect 21962 3016 21991 3029
rect 22043 3016 22072 3029
rect 22124 3016 22153 3029
rect 22205 3016 22234 3029
rect 22286 3016 22315 3029
rect 22367 3016 22396 3029
rect 22448 3016 22478 3068
rect 22530 3063 22559 3068
rect 22611 3063 22640 3068
rect 22692 3063 22721 3068
rect 22773 3063 22802 3068
rect 22854 3063 22883 3068
rect 22935 3063 22964 3068
rect 23016 3063 23046 3068
rect 22530 3029 22557 3063
rect 22611 3029 22629 3063
rect 22692 3029 22701 3063
rect 22879 3029 22883 3063
rect 22951 3029 22964 3063
rect 23023 3029 23046 3063
rect 22530 3016 22559 3029
rect 22611 3016 22640 3029
rect 22692 3016 22721 3029
rect 22773 3016 22802 3029
rect 22854 3016 22883 3029
rect 22935 3016 22964 3029
rect 23016 3016 23046 3029
rect 23098 3016 23127 3068
rect 23179 3063 23208 3068
rect 23260 3063 23289 3068
rect 23341 3063 23370 3068
rect 23422 3063 23451 3068
rect 23503 3063 23532 3068
rect 23584 3063 23614 3068
rect 23666 3063 23695 3068
rect 23179 3029 23205 3063
rect 23260 3029 23277 3063
rect 23341 3029 23349 3063
rect 23527 3029 23532 3063
rect 23599 3029 23614 3063
rect 23671 3029 23695 3063
rect 23179 3016 23208 3029
rect 23260 3016 23289 3029
rect 23341 3016 23370 3029
rect 23422 3016 23451 3029
rect 23503 3016 23532 3029
rect 23584 3016 23614 3029
rect 23666 3016 23695 3029
rect 23747 3016 23776 3068
rect 23828 3063 23857 3068
rect 23909 3063 23938 3068
rect 23990 3063 24019 3068
rect 24071 3063 24100 3068
rect 24152 3063 24182 3068
rect 24234 3063 24263 3068
rect 24315 3063 24344 3068
rect 23828 3029 23853 3063
rect 23909 3029 23925 3063
rect 23990 3029 23997 3063
rect 24175 3029 24182 3063
rect 24247 3029 24263 3063
rect 24319 3029 24344 3063
rect 23828 3016 23857 3029
rect 23909 3016 23938 3029
rect 23990 3016 24019 3029
rect 24071 3016 24100 3029
rect 24152 3016 24182 3029
rect 24234 3016 24263 3029
rect 24315 3016 24344 3029
rect 24396 3016 24425 3068
rect 24477 3063 24506 3068
rect 24558 3063 24587 3068
rect 24477 3029 24501 3063
rect 24558 3029 24573 3063
rect 24477 3016 24506 3029
rect 24558 3016 24587 3029
rect 24639 3016 24668 3068
rect 24720 3016 25079 3068
rect 3012 2976 25079 3016
rect 3012 2964 4768 2976
rect 4802 2964 4840 2976
rect 4874 2964 4912 2976
rect 4946 2964 4984 2976
rect 5018 2964 5056 2976
rect 5090 2964 5128 2976
rect 5162 2964 5200 2976
rect 5234 2964 5272 2976
rect 5306 2964 5344 2976
rect 5378 2964 5416 2976
rect 5450 2964 5488 2976
rect 5522 2964 5560 2976
rect 5594 2964 5632 2976
rect 5666 2964 5704 2976
rect 5738 2964 5776 2976
rect 5810 2964 5848 2976
rect 5882 2964 5920 2976
rect 5954 2964 5992 2976
rect 6026 2964 6064 2976
rect 6098 2964 6136 2976
rect 6170 2964 6208 2976
rect 6242 2964 6280 2976
rect 6314 2964 6352 2976
rect 6386 2964 6424 2976
rect 6458 2964 6496 2976
rect 6530 2964 6568 2976
rect 6602 2964 6640 2976
rect 6674 2964 6712 2976
rect 6746 2964 6784 2976
rect 6818 2964 6856 2976
rect 6890 2964 6928 2976
rect 6962 2964 7000 2976
rect 7034 2964 7072 2976
rect 7106 2964 7144 2976
rect 7178 2964 7216 2976
rect 7250 2964 7288 2976
rect 7322 2964 7360 2976
rect 7394 2964 7432 2976
rect 7466 2964 7504 2976
rect 7538 2964 7576 2976
rect 7610 2964 7648 2976
rect 7682 2964 7720 2976
rect 7754 2964 7792 2976
rect 7826 2964 7864 2976
rect 7898 2964 7936 2976
rect 7970 2964 8008 2976
rect 8042 2964 8080 2976
rect 8114 2964 8152 2976
rect 8186 2964 8224 2976
rect 8258 2964 8296 2976
rect 8330 2964 8368 2976
rect 8402 2964 8440 2976
rect 8474 2964 8512 2976
rect 8546 2964 8584 2976
rect 8618 2964 8656 2976
rect 8690 2964 8728 2976
rect 8762 2964 8800 2976
rect 8834 2964 8872 2976
rect 8906 2964 8944 2976
rect 8978 2964 9016 2976
rect 9050 2964 9088 2976
rect 9122 2964 9160 2976
rect 9194 2964 9232 2976
rect 9266 2964 9304 2976
rect 9338 2964 9376 2976
rect 9410 2964 9448 2976
rect 9482 2964 9520 2976
rect 9554 2964 9592 2976
rect 9626 2964 9664 2976
rect 9698 2964 9736 2976
rect 9770 2964 9808 2976
rect 9842 2964 9880 2976
rect 9914 2964 9952 2976
rect 9986 2964 10024 2976
rect 10058 2964 10096 2976
rect 10130 2964 10168 2976
rect 10202 2964 10240 2976
rect 10274 2964 10312 2976
rect 10346 2964 10384 2976
rect 10418 2964 10456 2976
rect 10490 2964 10528 2976
rect 10562 2964 10600 2976
rect 10634 2964 10672 2976
rect 10706 2964 10744 2976
rect 10778 2975 25079 2976
rect 10778 2964 12458 2975
rect 12492 2964 12530 2975
rect 12564 2964 12602 2975
rect 12636 2964 12674 2975
rect 12708 2964 12746 2975
rect 12780 2964 12818 2975
rect 12852 2964 12890 2975
rect 12924 2964 12962 2975
rect 12996 2964 13034 2975
rect 13068 2964 13106 2975
rect 13140 2964 13178 2975
rect 13212 2964 13250 2975
rect 13284 2964 13322 2975
rect 13356 2964 13394 2975
rect 13428 2964 13466 2975
rect 13500 2964 13538 2975
rect 13572 2964 13610 2975
rect 13644 2964 13682 2975
rect 13716 2964 13754 2975
rect 13788 2964 13826 2975
rect 13860 2964 13898 2975
rect 13932 2964 13970 2975
rect 14004 2964 14042 2975
rect 14076 2964 14114 2975
rect 14148 2964 14186 2975
rect 14220 2964 14258 2975
rect 14292 2964 14330 2975
rect 14364 2964 14402 2975
rect 14436 2964 14474 2975
rect 14508 2964 14546 2975
rect 14580 2964 14618 2975
rect 14652 2964 14690 2975
rect 14724 2964 14762 2975
rect 14796 2964 14834 2975
rect 14868 2964 14906 2975
rect 14940 2964 14978 2975
rect 15012 2964 15050 2975
rect 15084 2964 15122 2975
rect 15156 2964 15194 2975
rect 15228 2964 15266 2975
rect 15300 2964 15338 2975
rect 15372 2964 15410 2975
rect 15444 2964 15482 2975
rect 15516 2964 15554 2975
rect 15588 2964 15626 2975
rect 15660 2964 15698 2975
rect 15732 2964 15770 2975
rect 15804 2964 15842 2975
rect 15876 2964 15914 2975
rect 15948 2964 15986 2975
rect 16020 2964 16058 2975
rect 16092 2964 16130 2975
rect 16164 2964 16202 2975
rect 16236 2964 16274 2975
rect 16308 2964 16346 2975
rect 16380 2964 16418 2975
rect 16452 2964 16490 2975
rect 16524 2964 16562 2975
rect 16596 2964 16634 2975
rect 16668 2964 16706 2975
rect 16740 2964 16778 2975
rect 16812 2964 16850 2975
rect 16884 2964 16922 2975
rect 16956 2964 16994 2975
rect 17028 2964 17066 2975
rect 17100 2964 17138 2975
rect 17172 2964 17210 2975
rect 17244 2964 17282 2975
rect 17316 2964 17354 2975
rect 17388 2964 17426 2975
rect 17460 2964 17498 2975
rect 17532 2964 17570 2975
rect 17604 2964 17642 2975
rect 17676 2964 17714 2975
rect 17748 2964 17786 2975
rect 17820 2964 17858 2975
rect 17892 2964 17930 2975
rect 17964 2964 18002 2975
rect 18036 2964 18074 2975
rect 18108 2964 18146 2975
rect 18180 2964 18218 2975
rect 18252 2964 18290 2975
rect 18324 2964 18362 2975
rect 18396 2964 18434 2975
rect 18468 2964 18597 2975
rect 18631 2964 18669 2975
rect 18703 2964 18741 2975
rect 18775 2964 18813 2975
rect 18847 2964 18885 2975
rect 18919 2964 18957 2975
rect 18991 2964 19029 2975
rect 19063 2964 19101 2975
rect 19135 2964 19173 2975
rect 19207 2964 19245 2975
rect 19279 2964 19317 2975
rect 19351 2964 19389 2975
rect 19423 2964 19461 2975
rect 19495 2964 19533 2975
rect 19567 2964 19605 2975
rect 19639 2964 19677 2975
rect 19711 2964 19749 2975
rect 19783 2964 19821 2975
rect 19855 2964 19893 2975
rect 19927 2964 19965 2975
rect 19999 2964 20037 2975
rect 20071 2964 20109 2975
rect 20143 2964 20181 2975
rect 20215 2964 20253 2975
rect 20287 2964 20325 2975
rect 20359 2964 20397 2975
rect 20431 2964 20469 2975
rect 20503 2964 20541 2975
rect 20575 2964 20613 2975
rect 20647 2964 20685 2975
rect 20719 2964 20757 2975
rect 20791 2964 20829 2975
rect 20863 2964 20901 2975
rect 20935 2964 20973 2975
rect 21007 2964 21045 2975
rect 21079 2964 21117 2975
rect 21151 2964 21189 2975
rect 21223 2964 21261 2975
rect 21295 2964 21333 2975
rect 21367 2964 21405 2975
rect 21439 2964 21477 2975
rect 21511 2964 21549 2975
rect 21583 2964 21621 2975
rect 21655 2964 21693 2975
rect 21727 2964 21765 2975
rect 21799 2964 21837 2975
rect 21871 2964 21909 2975
rect 21943 2964 21981 2975
rect 22015 2964 22053 2975
rect 22087 2964 22125 2975
rect 22159 2964 22197 2975
rect 22231 2964 22269 2975
rect 22303 2964 22341 2975
rect 22375 2964 22413 2975
rect 22447 2964 22485 2975
rect 22519 2964 22557 2975
rect 22591 2964 22629 2975
rect 22663 2964 22701 2975
rect 22735 2964 22773 2975
rect 22807 2964 22845 2975
rect 22879 2964 22917 2975
rect 22951 2964 22989 2975
rect 23023 2964 23061 2975
rect 23095 2964 23133 2975
rect 23167 2964 23205 2975
rect 23239 2964 23277 2975
rect 23311 2964 23349 2975
rect 23383 2964 23421 2975
rect 23455 2964 23493 2975
rect 23527 2964 23565 2975
rect 23599 2964 23637 2975
rect 23671 2964 23709 2975
rect 23743 2964 23781 2975
rect 23815 2964 23853 2975
rect 23887 2964 23925 2975
rect 23959 2964 23997 2975
rect 24031 2964 24069 2975
rect 24103 2964 24141 2975
rect 24175 2964 24213 2975
rect 24247 2964 24285 2975
rect 24319 2964 24357 2975
rect 24391 2964 24429 2975
rect 24463 2964 24501 2975
rect 24535 2964 24573 2975
rect 24607 2964 25079 2975
rect 3012 2912 3038 2964
rect 3090 2912 3120 2964
rect 3172 2912 3201 2964
rect 3253 2912 3282 2964
rect 3334 2912 3363 2964
rect 3415 2912 3444 2964
rect 3496 2912 3525 2964
rect 3577 2912 3606 2964
rect 3658 2912 3688 2964
rect 3740 2912 3769 2964
rect 3821 2912 3850 2964
rect 3902 2912 3931 2964
rect 3983 2912 4012 2964
rect 4064 2912 4093 2964
rect 4145 2912 4174 2964
rect 4226 2912 4256 2964
rect 4308 2912 4337 2964
rect 4389 2912 4418 2964
rect 4470 2912 4499 2964
rect 4551 2912 4580 2964
rect 4632 2912 4661 2964
rect 4713 2912 4742 2964
rect 4802 2942 4824 2964
rect 4794 2912 4824 2942
rect 4876 2912 4905 2964
rect 4957 2942 4984 2964
rect 5038 2942 5056 2964
rect 5119 2942 5128 2964
rect 5306 2942 5310 2964
rect 5378 2942 5392 2964
rect 5450 2942 5473 2964
rect 4957 2912 4986 2942
rect 5038 2912 5067 2942
rect 5119 2912 5148 2942
rect 5200 2912 5229 2942
rect 5281 2912 5310 2942
rect 5362 2912 5392 2942
rect 5444 2912 5473 2942
rect 5525 2912 5554 2964
rect 5606 2942 5632 2964
rect 5687 2942 5704 2964
rect 5768 2942 5776 2964
rect 5954 2942 5960 2964
rect 6026 2942 6041 2964
rect 6098 2942 6122 2964
rect 5606 2912 5635 2942
rect 5687 2912 5716 2942
rect 5768 2912 5797 2942
rect 5849 2912 5878 2942
rect 5930 2912 5960 2942
rect 6012 2912 6041 2942
rect 6093 2912 6122 2942
rect 6174 2912 6203 2964
rect 6255 2942 6280 2964
rect 6336 2942 6352 2964
rect 6417 2942 6424 2964
rect 6602 2942 6609 2964
rect 6674 2942 6690 2964
rect 6746 2942 6771 2964
rect 6255 2912 6284 2942
rect 6336 2912 6365 2942
rect 6417 2912 6446 2942
rect 6498 2912 6528 2942
rect 6580 2912 6609 2942
rect 6661 2912 6690 2942
rect 6742 2912 6771 2942
rect 6823 2912 6852 2964
rect 6904 2942 6928 2964
rect 6985 2942 7000 2964
rect 7066 2942 7072 2964
rect 7250 2942 7258 2964
rect 7322 2942 7339 2964
rect 7394 2942 7420 2964
rect 6904 2912 6933 2942
rect 6985 2912 7014 2942
rect 7066 2912 7096 2942
rect 7148 2912 7177 2942
rect 7229 2912 7258 2942
rect 7310 2912 7339 2942
rect 7391 2912 7420 2942
rect 7472 2912 7501 2964
rect 7553 2942 7576 2964
rect 7634 2942 7648 2964
rect 7716 2942 7720 2964
rect 7898 2942 7907 2964
rect 7970 2942 7988 2964
rect 8042 2942 8069 2964
rect 7553 2912 7582 2942
rect 7634 2912 7664 2942
rect 7716 2912 7745 2942
rect 7797 2912 7826 2942
rect 7878 2912 7907 2942
rect 7959 2912 7988 2942
rect 8040 2912 8069 2942
rect 8121 2912 8150 2964
rect 8202 2942 8224 2964
rect 8284 2942 8296 2964
rect 8365 2942 8368 2964
rect 8474 2942 8475 2964
rect 8546 2942 8556 2964
rect 8618 2942 8637 2964
rect 8690 2942 8718 2964
rect 8202 2912 8232 2942
rect 8284 2912 8313 2942
rect 8365 2912 8394 2942
rect 8446 2912 8475 2942
rect 8527 2912 8556 2942
rect 8608 2912 8637 2942
rect 8689 2912 8718 2942
rect 8770 2912 8800 2964
rect 8852 2942 8872 2964
rect 8933 2942 8944 2964
rect 9014 2942 9016 2964
rect 9122 2942 9124 2964
rect 9194 2942 9205 2964
rect 9266 2942 9286 2964
rect 8852 2912 8881 2942
rect 8933 2912 8962 2942
rect 9014 2912 9043 2942
rect 9095 2912 9124 2942
rect 9176 2912 9205 2942
rect 9257 2912 9286 2942
rect 9338 2912 9368 2964
rect 9420 2942 9448 2964
rect 9501 2942 9520 2964
rect 9582 2942 9592 2964
rect 9663 2942 9664 2964
rect 9770 2942 9773 2964
rect 9842 2942 9854 2964
rect 9914 2942 9936 2964
rect 9420 2912 9449 2942
rect 9501 2912 9530 2942
rect 9582 2912 9611 2942
rect 9663 2912 9692 2942
rect 9744 2912 9773 2942
rect 9825 2912 9854 2942
rect 9906 2912 9936 2942
rect 9988 2912 10017 2964
rect 10069 2942 10096 2964
rect 10150 2942 10168 2964
rect 10231 2942 10240 2964
rect 10418 2942 10422 2964
rect 10490 2942 10504 2964
rect 10562 2942 10585 2964
rect 10069 2912 10098 2942
rect 10150 2912 10179 2942
rect 10231 2912 10260 2942
rect 10312 2912 10341 2942
rect 10393 2912 10422 2942
rect 10474 2912 10504 2942
rect 10556 2912 10585 2942
rect 10637 2912 10666 2964
rect 10718 2942 10744 2964
rect 10718 2912 10747 2942
rect 10799 2912 10828 2964
rect 10880 2912 10909 2964
rect 10961 2912 10990 2964
rect 11042 2912 11118 2964
rect 11170 2912 11199 2964
rect 11251 2912 11280 2964
rect 11332 2912 11361 2964
rect 11413 2912 11442 2964
rect 11494 2912 11523 2964
rect 11575 2912 11604 2964
rect 11656 2912 11686 2964
rect 11738 2912 11767 2964
rect 11819 2912 11848 2964
rect 11900 2912 11929 2964
rect 11981 2912 12010 2964
rect 12062 2912 12091 2964
rect 12143 2912 12172 2964
rect 12224 2912 12254 2964
rect 12306 2912 12335 2964
rect 12387 2912 12416 2964
rect 12492 2941 12497 2964
rect 12564 2941 12578 2964
rect 12636 2941 12659 2964
rect 12468 2912 12497 2941
rect 12549 2912 12578 2941
rect 12630 2912 12659 2941
rect 12711 2912 12740 2964
rect 12792 2941 12818 2964
rect 12874 2941 12890 2964
rect 12955 2941 12962 2964
rect 13140 2941 13146 2964
rect 13212 2941 13227 2964
rect 13284 2941 13308 2964
rect 12792 2912 12822 2941
rect 12874 2912 12903 2941
rect 12955 2912 12984 2941
rect 13036 2912 13065 2941
rect 13117 2912 13146 2941
rect 13198 2912 13227 2941
rect 13279 2912 13308 2941
rect 13360 2912 13390 2964
rect 13442 2941 13466 2964
rect 13523 2941 13538 2964
rect 13604 2941 13610 2964
rect 13788 2941 13795 2964
rect 13860 2941 13876 2964
rect 13932 2941 13958 2964
rect 13442 2912 13471 2941
rect 13523 2912 13552 2941
rect 13604 2912 13633 2941
rect 13685 2912 13714 2941
rect 13766 2912 13795 2941
rect 13847 2912 13876 2941
rect 13928 2912 13958 2941
rect 14010 2912 14039 2964
rect 14091 2941 14114 2964
rect 14172 2941 14186 2964
rect 14253 2941 14258 2964
rect 14436 2941 14444 2964
rect 14508 2941 14526 2964
rect 14580 2941 14607 2964
rect 14091 2912 14120 2941
rect 14172 2912 14201 2941
rect 14253 2912 14282 2941
rect 14334 2912 14363 2941
rect 14415 2912 14444 2941
rect 14496 2912 14526 2941
rect 14578 2912 14607 2941
rect 14659 2912 14688 2964
rect 14740 2941 14762 2964
rect 14821 2941 14834 2964
rect 14902 2941 14906 2964
rect 15084 2941 15094 2964
rect 15156 2941 15175 2964
rect 15228 2941 15256 2964
rect 14740 2912 14769 2941
rect 14821 2912 14850 2941
rect 14902 2912 14931 2941
rect 14983 2912 15012 2941
rect 15064 2912 15094 2941
rect 15146 2912 15175 2941
rect 15227 2912 15256 2941
rect 15308 2912 15337 2964
rect 15389 2941 15410 2964
rect 15470 2941 15482 2964
rect 15551 2941 15554 2964
rect 15660 2941 15662 2964
rect 15732 2941 15743 2964
rect 15804 2941 15824 2964
rect 15389 2912 15418 2941
rect 15470 2912 15499 2941
rect 15551 2912 15580 2941
rect 15632 2912 15662 2941
rect 15714 2912 15743 2941
rect 15795 2912 15824 2941
rect 15876 2912 15905 2964
rect 15957 2912 15986 2964
rect 16038 2941 16058 2964
rect 16119 2941 16130 2964
rect 16200 2941 16202 2964
rect 16308 2941 16311 2964
rect 16380 2941 16392 2964
rect 16452 2941 16473 2964
rect 16038 2912 16067 2941
rect 16119 2912 16148 2941
rect 16200 2912 16230 2941
rect 16282 2912 16311 2941
rect 16363 2912 16392 2941
rect 16444 2912 16473 2941
rect 16525 2912 16554 2964
rect 16606 2941 16634 2964
rect 16687 2941 16706 2964
rect 16768 2941 16778 2964
rect 16956 2941 16960 2964
rect 17028 2941 17041 2964
rect 17100 2941 17122 2964
rect 16606 2912 16635 2941
rect 16687 2912 16716 2941
rect 16768 2912 16798 2941
rect 16850 2912 16879 2941
rect 16931 2912 16960 2941
rect 17012 2912 17041 2941
rect 17093 2912 17122 2941
rect 17174 2912 17203 2964
rect 17255 2941 17282 2964
rect 17336 2941 17354 2964
rect 17418 2941 17426 2964
rect 17604 2941 17609 2964
rect 17676 2941 17690 2964
rect 17748 2941 17771 2964
rect 17255 2912 17284 2941
rect 17336 2912 17366 2941
rect 17418 2912 17447 2941
rect 17499 2912 17528 2941
rect 17580 2912 17609 2941
rect 17661 2912 17690 2941
rect 17742 2912 17771 2941
rect 17823 2912 17852 2964
rect 17904 2941 17930 2964
rect 17986 2941 18002 2964
rect 18067 2941 18074 2964
rect 18252 2941 18258 2964
rect 18324 2941 18339 2964
rect 18396 2941 18420 2964
rect 17904 2912 17934 2941
rect 17986 2912 18015 2941
rect 18067 2912 18096 2941
rect 18148 2912 18177 2941
rect 18229 2912 18258 2941
rect 18310 2912 18339 2941
rect 18391 2912 18420 2941
rect 18472 2912 18502 2964
rect 18554 2912 18583 2964
rect 18635 2912 18664 2964
rect 18716 2941 18741 2964
rect 18797 2941 18813 2964
rect 18878 2941 18885 2964
rect 19063 2941 19070 2964
rect 19135 2941 19151 2964
rect 19207 2941 19232 2964
rect 18716 2912 18745 2941
rect 18797 2912 18826 2941
rect 18878 2912 18907 2941
rect 18959 2912 18988 2941
rect 19040 2912 19070 2941
rect 19122 2912 19151 2941
rect 19203 2912 19232 2941
rect 19284 2912 19313 2964
rect 19365 2941 19389 2964
rect 19446 2941 19461 2964
rect 19527 2941 19533 2964
rect 19711 2941 19719 2964
rect 19783 2941 19800 2964
rect 19855 2941 19881 2964
rect 19365 2912 19394 2941
rect 19446 2912 19475 2941
rect 19527 2912 19556 2941
rect 19608 2912 19638 2941
rect 19690 2912 19719 2941
rect 19771 2912 19800 2941
rect 19852 2912 19881 2941
rect 19933 2912 19962 2964
rect 20014 2941 20037 2964
rect 20095 2941 20109 2964
rect 20176 2941 20181 2964
rect 20359 2941 20368 2964
rect 20431 2941 20449 2964
rect 20503 2941 20530 2964
rect 20014 2912 20043 2941
rect 20095 2912 20124 2941
rect 20176 2912 20206 2941
rect 20258 2912 20287 2941
rect 20339 2912 20368 2941
rect 20420 2912 20449 2941
rect 20501 2912 20530 2941
rect 20582 2912 20611 2964
rect 20663 2941 20685 2964
rect 20744 2941 20757 2964
rect 20826 2941 20829 2964
rect 20935 2941 20936 2964
rect 21007 2941 21017 2964
rect 21079 2941 21098 2964
rect 21151 2941 21179 2964
rect 20663 2912 20692 2941
rect 20744 2912 20774 2941
rect 20826 2912 20855 2941
rect 20907 2912 20936 2941
rect 20988 2912 21017 2941
rect 21069 2912 21098 2941
rect 21150 2912 21179 2941
rect 21231 2912 21260 2964
rect 21312 2941 21333 2964
rect 21394 2941 21405 2964
rect 21475 2941 21477 2964
rect 21583 2941 21585 2964
rect 21655 2941 21666 2964
rect 21727 2941 21747 2964
rect 21312 2912 21342 2941
rect 21394 2912 21423 2941
rect 21475 2912 21504 2941
rect 21556 2912 21585 2941
rect 21637 2912 21666 2941
rect 21718 2912 21747 2941
rect 21799 2912 21828 2964
rect 21880 2941 21909 2964
rect 21962 2941 21981 2964
rect 22043 2941 22053 2964
rect 22124 2941 22125 2964
rect 22231 2941 22234 2964
rect 22303 2941 22315 2964
rect 22375 2941 22396 2964
rect 21880 2912 21910 2941
rect 21962 2912 21991 2941
rect 22043 2912 22072 2941
rect 22124 2912 22153 2941
rect 22205 2912 22234 2941
rect 22286 2912 22315 2941
rect 22367 2912 22396 2941
rect 22448 2912 22478 2964
rect 22530 2941 22557 2964
rect 22611 2941 22629 2964
rect 22692 2941 22701 2964
rect 22879 2941 22883 2964
rect 22951 2941 22964 2964
rect 23023 2941 23046 2964
rect 22530 2912 22559 2941
rect 22611 2912 22640 2941
rect 22692 2912 22721 2941
rect 22773 2912 22802 2941
rect 22854 2912 22883 2941
rect 22935 2912 22964 2941
rect 23016 2912 23046 2941
rect 23098 2912 23127 2964
rect 23179 2941 23205 2964
rect 23260 2941 23277 2964
rect 23341 2941 23349 2964
rect 23527 2941 23532 2964
rect 23599 2941 23614 2964
rect 23671 2941 23695 2964
rect 23179 2912 23208 2941
rect 23260 2912 23289 2941
rect 23341 2912 23370 2941
rect 23422 2912 23451 2941
rect 23503 2912 23532 2941
rect 23584 2912 23614 2941
rect 23666 2912 23695 2941
rect 23747 2912 23776 2964
rect 23828 2941 23853 2964
rect 23909 2941 23925 2964
rect 23990 2941 23997 2964
rect 24175 2941 24182 2964
rect 24247 2941 24263 2964
rect 24319 2941 24344 2964
rect 23828 2912 23857 2941
rect 23909 2912 23938 2941
rect 23990 2912 24019 2941
rect 24071 2912 24100 2941
rect 24152 2912 24182 2941
rect 24234 2912 24263 2941
rect 24315 2912 24344 2941
rect 24396 2912 24425 2964
rect 24477 2941 24501 2964
rect 24558 2941 24573 2964
rect 24477 2912 24506 2941
rect 24558 2912 24587 2941
rect 24639 2912 24668 2964
rect 24720 2912 25079 2964
rect 3012 2905 25079 2912
rect 4760 2883 10808 2905
rect 4760 2816 4780 2883
rect 4808 2833 4850 2837
rect 4804 2660 4850 2833
rect 5040 2687 5086 2864
rect 5276 2672 5322 2849
rect 5512 2687 5558 2876
rect 5630 2675 5676 2687
rect 5754 2675 5788 2852
rect 5984 2687 6030 2883
rect 5866 2675 5912 2687
rect 5630 2667 5636 2675
rect 5670 2667 5676 2675
rect 5866 2667 5872 2675
rect 5906 2667 5912 2675
rect 6102 2675 6148 2687
rect 6220 2684 6266 2861
rect 6102 2667 6108 2675
rect 6142 2667 6148 2675
rect 6338 2675 6384 2687
rect 6462 2675 6496 2883
rect 6574 2675 6620 2687
rect 6338 2667 6344 2675
rect 6378 2667 6384 2675
rect 6574 2667 6580 2675
rect 6614 2667 6620 2675
rect 6802 2672 6848 2849
rect 7038 2687 7084 2876
rect 7274 2684 7320 2861
rect 7510 2687 7556 2883
rect 7746 2687 7792 2864
rect 7982 2687 8028 2883
rect 8218 2687 8264 2873
rect 8454 2687 8500 2883
rect 7392 2675 7438 2687
rect 7392 2667 7398 2675
rect 7432 2667 7438 2675
rect 7864 2675 7910 2687
rect 7864 2667 7870 2675
rect 7904 2667 7910 2675
rect 8336 2675 8382 2687
rect 8336 2667 8342 2675
rect 8376 2667 8382 2675
rect 8800 2672 8846 2849
rect 9036 2687 9082 2876
rect 8918 2675 8964 2687
rect 9272 2684 9318 2861
rect 9508 2687 9554 2883
rect 9744 2687 9790 2864
rect 9980 2687 10026 2883
rect 10216 2687 10262 2873
rect 10452 2687 10498 2883
rect 12450 2881 25079 2905
rect 12450 2869 23858 2881
rect 23859 2871 25079 2881
rect 12450 2835 18598 2869
rect 18632 2835 23858 2869
rect 12450 2815 23858 2835
rect 15621 2687 16451 2815
rect 8918 2667 8924 2675
rect 8958 2667 8964 2675
rect 9390 2675 9436 2687
rect 9390 2667 9396 2675
rect 9430 2667 9436 2675
rect 9862 2675 9908 2687
rect 9862 2667 9868 2675
rect 9902 2667 9908 2675
rect 10334 2675 10380 2687
rect 10334 2667 10340 2675
rect 10374 2667 10380 2675
rect 12730 2674 12776 2686
rect 4909 2107 4919 2667
rect 4971 2107 4981 2667
rect 5145 2107 5155 2667
rect 5207 2107 5217 2667
rect 5381 2107 5391 2667
rect 5443 2107 5453 2667
rect 5617 2107 5627 2667
rect 5679 2107 5689 2667
rect 5853 2107 5863 2667
rect 5915 2107 5925 2667
rect 6089 2107 6099 2667
rect 6151 2107 6161 2667
rect 6325 2107 6335 2667
rect 6387 2107 6397 2667
rect 6561 2107 6571 2667
rect 6623 2107 6633 2667
rect 6907 2107 6917 2667
rect 6969 2107 6979 2667
rect 7143 2107 7153 2667
rect 7205 2107 7215 2667
rect 7379 2107 7389 2667
rect 7441 2107 7451 2667
rect 7615 2107 7625 2667
rect 7677 2107 7687 2667
rect 7851 2107 7861 2667
rect 7913 2107 7923 2667
rect 8087 2107 8097 2667
rect 8149 2107 8159 2667
rect 8323 2107 8333 2667
rect 8385 2107 8395 2667
rect 8559 2107 8569 2667
rect 8621 2107 8631 2667
rect 8905 2107 8915 2667
rect 8967 2107 8977 2667
rect 9141 2107 9151 2667
rect 9203 2107 9213 2667
rect 9377 2107 9387 2667
rect 9439 2107 9449 2667
rect 9613 2107 9623 2667
rect 9675 2107 9685 2667
rect 9849 2107 9859 2667
rect 9911 2107 9921 2667
rect 10085 2107 10095 2667
rect 10147 2107 10157 2667
rect 10321 2107 10331 2667
rect 10383 2107 10393 2667
rect 10557 2107 10567 2667
rect 10619 2107 10629 2667
rect 12730 2666 12736 2674
rect 12770 2666 12776 2674
rect 12848 2674 12894 2686
rect 12848 2666 12854 2674
rect 12888 2666 12894 2674
rect 12966 2674 13012 2686
rect 12966 2666 12972 2674
rect 13006 2666 13012 2674
rect 13084 2674 13130 2686
rect 13084 2666 13090 2674
rect 13124 2666 13130 2674
rect 13202 2674 13248 2686
rect 13202 2666 13208 2674
rect 13242 2666 13248 2674
rect 13320 2674 13366 2686
rect 13320 2666 13326 2674
rect 13360 2666 13366 2674
rect 13438 2674 13484 2686
rect 13438 2666 13444 2674
rect 13478 2666 13484 2674
rect 13556 2674 13602 2686
rect 13556 2666 13562 2674
rect 13596 2666 13602 2674
rect 13674 2674 13720 2686
rect 13674 2666 13680 2674
rect 13714 2666 13720 2674
rect 13792 2674 13838 2686
rect 13792 2666 13798 2674
rect 13832 2666 13838 2674
rect 13910 2674 13956 2686
rect 13910 2666 13916 2674
rect 13950 2666 13956 2674
rect 14028 2674 14074 2686
rect 14028 2666 14034 2674
rect 14068 2666 14074 2674
rect 14146 2674 14192 2686
rect 14146 2666 14152 2674
rect 14186 2666 14192 2674
rect 14264 2674 14310 2686
rect 14264 2666 14270 2674
rect 14304 2666 14310 2674
rect 14382 2674 14428 2686
rect 14382 2666 14388 2674
rect 14422 2666 14428 2674
rect 14500 2674 14546 2686
rect 14500 2666 14506 2674
rect 14540 2666 14546 2674
rect 14618 2674 14664 2686
rect 14618 2666 14624 2674
rect 14658 2666 14664 2674
rect 14736 2674 14782 2686
rect 14736 2666 14742 2674
rect 14776 2666 14782 2674
rect 14854 2674 14900 2686
rect 14854 2666 14860 2674
rect 14894 2666 14900 2674
rect 14972 2674 15018 2686
rect 14972 2666 14978 2674
rect 15012 2666 15018 2674
rect 15090 2674 15136 2686
rect 15090 2666 15096 2674
rect 15130 2666 15136 2674
rect 15208 2674 15254 2686
rect 15208 2666 15214 2674
rect 15248 2666 15254 2674
rect 15326 2674 15372 2686
rect 15326 2666 15332 2674
rect 15366 2666 15372 2674
rect 15444 2674 15490 2686
rect 15444 2666 15450 2674
rect 15484 2666 15490 2674
rect 5630 2099 5636 2107
rect 5670 2099 5676 2107
rect 5630 2087 5676 2099
rect 5866 2099 5872 2107
rect 5906 2099 5912 2107
rect 5866 2087 5912 2099
rect 6102 2099 6108 2107
rect 6142 2099 6148 2107
rect 6102 2087 6148 2099
rect 6338 2099 6344 2107
rect 6378 2099 6384 2107
rect 6338 2087 6384 2099
rect 6574 2099 6580 2107
rect 6614 2099 6620 2107
rect 6574 2087 6620 2099
rect 7392 2099 7398 2107
rect 7432 2099 7438 2107
rect 7392 2087 7438 2099
rect 7864 2099 7870 2107
rect 7904 2099 7910 2107
rect 7864 2087 7910 2099
rect 8336 2099 8342 2107
rect 8376 2099 8382 2107
rect 8336 2087 8382 2099
rect 8918 2099 8924 2107
rect 8958 2099 8964 2107
rect 8918 2087 8964 2099
rect 9390 2099 9396 2107
rect 9430 2099 9436 2107
rect 9390 2087 9436 2099
rect 9862 2099 9868 2107
rect 9902 2099 9908 2107
rect 9862 2087 9908 2099
rect 10334 2099 10340 2107
rect 10374 2099 10380 2107
rect 12481 2106 12491 2666
rect 12543 2106 12553 2666
rect 12599 2106 12609 2666
rect 12661 2106 12671 2666
rect 12717 2106 12727 2666
rect 12779 2106 12789 2666
rect 12835 2106 12845 2666
rect 12897 2106 12907 2666
rect 12953 2106 12963 2666
rect 13015 2106 13025 2666
rect 13071 2106 13081 2666
rect 13133 2106 13143 2666
rect 13189 2106 13199 2666
rect 13251 2106 13261 2666
rect 13307 2106 13317 2666
rect 13369 2106 13379 2666
rect 13425 2106 13435 2666
rect 13487 2106 13497 2666
rect 13543 2106 13553 2666
rect 13605 2106 13615 2666
rect 13661 2106 13671 2666
rect 13723 2106 13733 2666
rect 13779 2106 13789 2666
rect 13841 2106 13851 2666
rect 13897 2106 13907 2666
rect 13959 2106 13969 2666
rect 14015 2106 14025 2666
rect 14077 2106 14087 2666
rect 14133 2106 14143 2666
rect 14195 2106 14205 2666
rect 14251 2106 14261 2666
rect 14313 2106 14323 2666
rect 14369 2106 14379 2666
rect 14431 2106 14441 2666
rect 14487 2106 14497 2666
rect 14549 2106 14559 2666
rect 14605 2106 14615 2666
rect 14667 2106 14677 2666
rect 14723 2106 14733 2666
rect 14785 2106 14795 2666
rect 14841 2106 14851 2666
rect 14903 2106 14913 2666
rect 14959 2106 14969 2666
rect 15021 2106 15031 2666
rect 15077 2106 15087 2666
rect 15139 2106 15149 2666
rect 15195 2106 15205 2666
rect 15257 2106 15267 2666
rect 15313 2106 15323 2666
rect 15375 2106 15385 2666
rect 15431 2106 15441 2666
rect 15493 2106 15503 2666
rect 15621 2653 15659 2687
rect 15693 2653 15731 2687
rect 15765 2653 15803 2687
rect 15837 2653 15875 2687
rect 15909 2653 15947 2687
rect 15981 2653 16019 2687
rect 16053 2653 16091 2687
rect 16125 2653 16163 2687
rect 16197 2653 16235 2687
rect 16269 2653 16307 2687
rect 16341 2653 16379 2687
rect 16413 2653 16451 2687
rect 19744 2687 20574 2815
rect 23903 2707 25079 2871
rect 16853 2674 16899 2686
rect 16853 2666 16859 2674
rect 16893 2666 16899 2674
rect 16971 2674 17017 2686
rect 16971 2666 16977 2674
rect 17011 2666 17017 2674
rect 17089 2674 17135 2686
rect 17089 2666 17095 2674
rect 17129 2666 17135 2674
rect 17207 2674 17253 2686
rect 17207 2666 17213 2674
rect 17247 2666 17253 2674
rect 17325 2674 17371 2686
rect 17325 2666 17331 2674
rect 17365 2666 17371 2674
rect 17443 2674 17489 2686
rect 17443 2666 17449 2674
rect 17483 2666 17489 2674
rect 17561 2674 17607 2686
rect 17561 2666 17567 2674
rect 17601 2666 17607 2674
rect 17679 2674 17725 2686
rect 17679 2666 17685 2674
rect 17719 2666 17725 2674
rect 17797 2674 17843 2686
rect 17797 2666 17803 2674
rect 17837 2666 17843 2674
rect 17915 2674 17961 2686
rect 17915 2666 17921 2674
rect 17955 2666 17961 2674
rect 18033 2674 18079 2686
rect 18033 2666 18039 2674
rect 18073 2666 18079 2674
rect 18151 2674 18197 2686
rect 18151 2666 18157 2674
rect 18191 2666 18197 2674
rect 18269 2674 18315 2686
rect 18269 2666 18275 2674
rect 18309 2666 18315 2674
rect 18387 2674 18433 2686
rect 18387 2666 18393 2674
rect 18427 2666 18433 2674
rect 18505 2674 18551 2686
rect 18505 2666 18511 2674
rect 18545 2666 18551 2674
rect 18623 2674 18669 2686
rect 18623 2666 18629 2674
rect 18663 2666 18669 2674
rect 18741 2674 18787 2686
rect 18741 2666 18747 2674
rect 18781 2666 18787 2674
rect 18859 2674 18905 2686
rect 18859 2666 18865 2674
rect 18899 2666 18905 2674
rect 18977 2674 19023 2686
rect 18977 2666 18983 2674
rect 19017 2666 19023 2674
rect 19095 2674 19141 2686
rect 19095 2666 19101 2674
rect 19135 2666 19141 2674
rect 19213 2674 19259 2686
rect 19213 2666 19219 2674
rect 19253 2666 19259 2674
rect 19331 2674 19377 2686
rect 19331 2666 19337 2674
rect 19371 2666 19377 2674
rect 19449 2674 19495 2686
rect 19449 2666 19455 2674
rect 19489 2666 19495 2674
rect 19567 2674 19613 2686
rect 19567 2666 19573 2674
rect 19607 2666 19613 2674
rect 15621 2613 16451 2653
rect 15621 2579 15659 2613
rect 15693 2579 15731 2613
rect 15765 2579 15803 2613
rect 15837 2579 15875 2613
rect 15909 2579 15947 2613
rect 15981 2579 16019 2613
rect 16053 2579 16091 2613
rect 16125 2579 16163 2613
rect 16197 2579 16235 2613
rect 16269 2579 16307 2613
rect 16341 2579 16379 2613
rect 16413 2579 16451 2613
rect 15621 2539 16451 2579
rect 15621 2505 15659 2539
rect 15693 2505 15731 2539
rect 15765 2505 15803 2539
rect 15837 2505 15875 2539
rect 15909 2505 15947 2539
rect 15981 2505 16019 2539
rect 16053 2505 16091 2539
rect 16125 2505 16163 2539
rect 16197 2505 16235 2539
rect 16269 2505 16307 2539
rect 16341 2505 16379 2539
rect 16413 2505 16451 2539
rect 15621 2465 16451 2505
rect 15621 2431 15659 2465
rect 15693 2431 15731 2465
rect 15765 2431 15803 2465
rect 15837 2431 15875 2465
rect 15909 2431 15947 2465
rect 15981 2431 16019 2465
rect 16053 2431 16091 2465
rect 16125 2431 16163 2465
rect 16197 2431 16235 2465
rect 16269 2431 16307 2465
rect 16341 2431 16379 2465
rect 16413 2431 16451 2465
rect 15621 2391 16451 2431
rect 15621 2357 15659 2391
rect 15693 2357 15731 2391
rect 15765 2357 15803 2391
rect 15837 2357 15875 2391
rect 15909 2357 15947 2391
rect 15981 2357 16019 2391
rect 16053 2357 16091 2391
rect 16125 2357 16163 2391
rect 16197 2357 16235 2391
rect 16269 2357 16307 2391
rect 16341 2357 16379 2391
rect 16413 2357 16451 2391
rect 15621 2317 16451 2357
rect 15621 2283 15659 2317
rect 15693 2283 15731 2317
rect 15765 2283 15803 2317
rect 15837 2283 15875 2317
rect 15909 2283 15947 2317
rect 15981 2283 16019 2317
rect 16053 2283 16091 2317
rect 16125 2283 16163 2317
rect 16197 2283 16235 2317
rect 16269 2283 16307 2317
rect 16341 2283 16379 2317
rect 16413 2283 16451 2317
rect 15621 2243 16451 2283
rect 15621 2209 15659 2243
rect 15693 2209 15731 2243
rect 15765 2209 15803 2243
rect 15837 2209 15875 2243
rect 15909 2209 15947 2243
rect 15981 2209 16019 2243
rect 16053 2209 16091 2243
rect 16125 2209 16163 2243
rect 16197 2209 16235 2243
rect 16269 2209 16307 2243
rect 16341 2209 16379 2243
rect 16413 2209 16451 2243
rect 15621 2169 16451 2209
rect 15621 2135 15659 2169
rect 15693 2135 15731 2169
rect 15765 2135 15803 2169
rect 15837 2135 15875 2169
rect 15909 2135 15947 2169
rect 15981 2135 16019 2169
rect 16053 2135 16091 2169
rect 16125 2135 16163 2169
rect 16197 2135 16235 2169
rect 16269 2135 16307 2169
rect 16341 2135 16379 2169
rect 16413 2135 16451 2169
rect 10334 2087 10380 2099
rect 12730 2098 12736 2106
rect 12770 2098 12776 2106
rect 12730 2086 12776 2098
rect 12848 2098 12854 2106
rect 12888 2098 12894 2106
rect 12848 2086 12894 2098
rect 12966 2098 12972 2106
rect 13006 2098 13012 2106
rect 12966 2086 13012 2098
rect 13084 2098 13090 2106
rect 13124 2098 13130 2106
rect 13084 2086 13130 2098
rect 13202 2098 13208 2106
rect 13242 2098 13248 2106
rect 13202 2086 13248 2098
rect 13320 2098 13326 2106
rect 13360 2098 13366 2106
rect 13320 2086 13366 2098
rect 13438 2098 13444 2106
rect 13478 2098 13484 2106
rect 13438 2086 13484 2098
rect 13556 2098 13562 2106
rect 13596 2098 13602 2106
rect 13556 2086 13602 2098
rect 13674 2098 13680 2106
rect 13714 2098 13720 2106
rect 13674 2086 13720 2098
rect 13792 2098 13798 2106
rect 13832 2098 13838 2106
rect 13792 2086 13838 2098
rect 13910 2098 13916 2106
rect 13950 2098 13956 2106
rect 13910 2086 13956 2098
rect 14028 2098 14034 2106
rect 14068 2098 14074 2106
rect 14028 2086 14074 2098
rect 14146 2098 14152 2106
rect 14186 2098 14192 2106
rect 14146 2086 14192 2098
rect 14264 2098 14270 2106
rect 14304 2098 14310 2106
rect 14264 2086 14310 2098
rect 14382 2098 14388 2106
rect 14422 2098 14428 2106
rect 14382 2086 14428 2098
rect 14500 2098 14506 2106
rect 14540 2098 14546 2106
rect 14500 2086 14546 2098
rect 14618 2098 14624 2106
rect 14658 2098 14664 2106
rect 14618 2086 14664 2098
rect 14736 2098 14742 2106
rect 14776 2098 14782 2106
rect 14736 2086 14782 2098
rect 14854 2098 14860 2106
rect 14894 2098 14900 2106
rect 14854 2086 14900 2098
rect 14972 2098 14978 2106
rect 15012 2098 15018 2106
rect 14972 2086 15018 2098
rect 15090 2098 15096 2106
rect 15130 2098 15136 2106
rect 15090 2086 15136 2098
rect 15208 2098 15214 2106
rect 15248 2098 15254 2106
rect 15208 2086 15254 2098
rect 15326 2098 15332 2106
rect 15366 2098 15372 2106
rect 15326 2086 15372 2098
rect 15444 2098 15450 2106
rect 15484 2098 15490 2106
rect 15444 2086 15490 2098
rect 15621 2095 16451 2135
rect 16604 2106 16614 2666
rect 16666 2106 16676 2666
rect 16722 2106 16732 2666
rect 16784 2106 16794 2666
rect 16840 2106 16850 2666
rect 16902 2106 16912 2666
rect 16958 2106 16968 2666
rect 17020 2106 17030 2666
rect 17076 2106 17086 2666
rect 17138 2106 17148 2666
rect 17194 2106 17204 2666
rect 17256 2106 17266 2666
rect 17312 2106 17322 2666
rect 17374 2106 17384 2666
rect 17430 2106 17440 2666
rect 17492 2106 17502 2666
rect 17548 2106 17558 2666
rect 17610 2106 17620 2666
rect 17666 2106 17676 2666
rect 17728 2106 17738 2666
rect 17784 2106 17794 2666
rect 17846 2106 17856 2666
rect 17902 2106 17912 2666
rect 17964 2106 17974 2666
rect 18020 2106 18030 2666
rect 18082 2106 18092 2666
rect 18138 2106 18148 2666
rect 18200 2106 18210 2666
rect 18256 2106 18266 2666
rect 18318 2106 18328 2666
rect 18374 2106 18384 2666
rect 18436 2106 18446 2666
rect 18492 2106 18502 2666
rect 18554 2106 18564 2666
rect 18610 2106 18620 2666
rect 18672 2106 18682 2666
rect 18728 2106 18738 2666
rect 18790 2106 18800 2666
rect 18846 2106 18856 2666
rect 18908 2106 18918 2666
rect 18964 2106 18974 2666
rect 19026 2106 19036 2666
rect 19082 2106 19092 2666
rect 19144 2106 19154 2666
rect 19200 2106 19210 2666
rect 19262 2106 19272 2666
rect 19318 2106 19328 2666
rect 19380 2106 19390 2666
rect 19436 2106 19446 2666
rect 19498 2106 19508 2666
rect 19554 2106 19564 2666
rect 19616 2106 19626 2666
rect 19744 2653 19782 2687
rect 19816 2653 19854 2687
rect 19888 2653 19926 2687
rect 19960 2653 19998 2687
rect 20032 2653 20070 2687
rect 20104 2653 20142 2687
rect 20176 2653 20214 2687
rect 20248 2653 20286 2687
rect 20320 2653 20358 2687
rect 20392 2653 20430 2687
rect 20464 2653 20502 2687
rect 20536 2653 20574 2687
rect 23867 2687 25079 2707
rect 20976 2674 21022 2686
rect 20976 2666 20982 2674
rect 21016 2666 21022 2674
rect 21094 2674 21140 2686
rect 21094 2666 21100 2674
rect 21134 2666 21140 2674
rect 21212 2674 21258 2686
rect 21212 2666 21218 2674
rect 21252 2666 21258 2674
rect 21330 2674 21376 2686
rect 21330 2666 21336 2674
rect 21370 2666 21376 2674
rect 21448 2674 21494 2686
rect 21448 2666 21454 2674
rect 21488 2666 21494 2674
rect 21566 2674 21612 2686
rect 21566 2666 21572 2674
rect 21606 2666 21612 2674
rect 21684 2674 21730 2686
rect 21684 2666 21690 2674
rect 21724 2666 21730 2674
rect 21802 2674 21848 2686
rect 21802 2666 21808 2674
rect 21842 2666 21848 2674
rect 21920 2674 21966 2686
rect 21920 2666 21926 2674
rect 21960 2666 21966 2674
rect 22038 2674 22084 2686
rect 22038 2666 22044 2674
rect 22078 2666 22084 2674
rect 22156 2674 22202 2686
rect 22156 2666 22162 2674
rect 22196 2666 22202 2674
rect 22274 2674 22320 2686
rect 22274 2666 22280 2674
rect 22314 2666 22320 2674
rect 22392 2674 22438 2686
rect 22392 2666 22398 2674
rect 22432 2666 22438 2674
rect 22510 2674 22556 2686
rect 22510 2666 22516 2674
rect 22550 2666 22556 2674
rect 22628 2674 22674 2686
rect 22628 2666 22634 2674
rect 22668 2666 22674 2674
rect 22746 2674 22792 2686
rect 22746 2666 22752 2674
rect 22786 2666 22792 2674
rect 22864 2674 22910 2686
rect 22864 2666 22870 2674
rect 22904 2666 22910 2674
rect 22982 2674 23028 2686
rect 22982 2666 22988 2674
rect 23022 2666 23028 2674
rect 23100 2674 23146 2686
rect 23100 2666 23106 2674
rect 23140 2666 23146 2674
rect 23218 2674 23264 2686
rect 23218 2666 23224 2674
rect 23258 2666 23264 2674
rect 23336 2674 23382 2686
rect 23336 2666 23342 2674
rect 23376 2666 23382 2674
rect 23454 2674 23500 2686
rect 23454 2666 23460 2674
rect 23494 2666 23500 2674
rect 23572 2674 23618 2686
rect 23572 2666 23578 2674
rect 23612 2666 23618 2674
rect 23690 2674 23736 2686
rect 23690 2666 23696 2674
rect 23730 2666 23736 2674
rect 19744 2613 20574 2653
rect 19744 2579 19782 2613
rect 19816 2579 19854 2613
rect 19888 2579 19926 2613
rect 19960 2579 19998 2613
rect 20032 2579 20070 2613
rect 20104 2579 20142 2613
rect 20176 2579 20214 2613
rect 20248 2579 20286 2613
rect 20320 2579 20358 2613
rect 20392 2579 20430 2613
rect 20464 2579 20502 2613
rect 20536 2579 20574 2613
rect 19744 2539 20574 2579
rect 19744 2505 19782 2539
rect 19816 2505 19854 2539
rect 19888 2505 19926 2539
rect 19960 2505 19998 2539
rect 20032 2505 20070 2539
rect 20104 2505 20142 2539
rect 20176 2505 20214 2539
rect 20248 2505 20286 2539
rect 20320 2505 20358 2539
rect 20392 2505 20430 2539
rect 20464 2505 20502 2539
rect 20536 2505 20574 2539
rect 19744 2465 20574 2505
rect 19744 2431 19782 2465
rect 19816 2431 19854 2465
rect 19888 2431 19926 2465
rect 19960 2431 19998 2465
rect 20032 2431 20070 2465
rect 20104 2431 20142 2465
rect 20176 2431 20214 2465
rect 20248 2431 20286 2465
rect 20320 2431 20358 2465
rect 20392 2431 20430 2465
rect 20464 2431 20502 2465
rect 20536 2431 20574 2465
rect 19744 2391 20574 2431
rect 19744 2357 19782 2391
rect 19816 2357 19854 2391
rect 19888 2357 19926 2391
rect 19960 2357 19998 2391
rect 20032 2357 20070 2391
rect 20104 2357 20142 2391
rect 20176 2357 20214 2391
rect 20248 2357 20286 2391
rect 20320 2357 20358 2391
rect 20392 2357 20430 2391
rect 20464 2357 20502 2391
rect 20536 2357 20574 2391
rect 19744 2317 20574 2357
rect 19744 2283 19782 2317
rect 19816 2283 19854 2317
rect 19888 2283 19926 2317
rect 19960 2283 19998 2317
rect 20032 2283 20070 2317
rect 20104 2283 20142 2317
rect 20176 2283 20214 2317
rect 20248 2283 20286 2317
rect 20320 2283 20358 2317
rect 20392 2283 20430 2317
rect 20464 2283 20502 2317
rect 20536 2283 20574 2317
rect 19744 2243 20574 2283
rect 19744 2209 19782 2243
rect 19816 2209 19854 2243
rect 19888 2209 19926 2243
rect 19960 2209 19998 2243
rect 20032 2209 20070 2243
rect 20104 2209 20142 2243
rect 20176 2209 20214 2243
rect 20248 2209 20286 2243
rect 20320 2209 20358 2243
rect 20392 2209 20430 2243
rect 20464 2209 20502 2243
rect 20536 2209 20574 2243
rect 19744 2169 20574 2209
rect 19744 2135 19782 2169
rect 19816 2135 19854 2169
rect 19888 2135 19926 2169
rect 19960 2135 19998 2169
rect 20032 2135 20070 2169
rect 20104 2135 20142 2169
rect 20176 2135 20214 2169
rect 20248 2135 20286 2169
rect 20320 2135 20358 2169
rect 20392 2135 20430 2169
rect 20464 2135 20502 2169
rect 20536 2135 20574 2169
rect 15621 2061 15659 2095
rect 15693 2061 15731 2095
rect 15765 2061 15803 2095
rect 15837 2061 15875 2095
rect 15909 2061 15947 2095
rect 15981 2061 16019 2095
rect 16053 2061 16091 2095
rect 16125 2061 16163 2095
rect 16197 2061 16235 2095
rect 16269 2061 16307 2095
rect 16341 2061 16379 2095
rect 16413 2061 16451 2095
rect 16853 2098 16859 2106
rect 16893 2098 16899 2106
rect 16853 2086 16899 2098
rect 16971 2098 16977 2106
rect 17011 2098 17017 2106
rect 16971 2086 17017 2098
rect 17089 2098 17095 2106
rect 17129 2098 17135 2106
rect 17089 2086 17135 2098
rect 17207 2098 17213 2106
rect 17247 2098 17253 2106
rect 17207 2086 17253 2098
rect 17325 2098 17331 2106
rect 17365 2098 17371 2106
rect 17325 2086 17371 2098
rect 17443 2098 17449 2106
rect 17483 2098 17489 2106
rect 17443 2086 17489 2098
rect 17561 2098 17567 2106
rect 17601 2098 17607 2106
rect 17561 2086 17607 2098
rect 17679 2098 17685 2106
rect 17719 2098 17725 2106
rect 17679 2086 17725 2098
rect 17797 2098 17803 2106
rect 17837 2098 17843 2106
rect 17797 2086 17843 2098
rect 17915 2098 17921 2106
rect 17955 2098 17961 2106
rect 17915 2086 17961 2098
rect 18033 2098 18039 2106
rect 18073 2098 18079 2106
rect 18033 2086 18079 2098
rect 18151 2098 18157 2106
rect 18191 2098 18197 2106
rect 18151 2086 18197 2098
rect 18269 2098 18275 2106
rect 18309 2098 18315 2106
rect 18269 2086 18315 2098
rect 18387 2098 18393 2106
rect 18427 2098 18433 2106
rect 18387 2086 18433 2098
rect 18505 2098 18511 2106
rect 18545 2098 18551 2106
rect 18505 2086 18551 2098
rect 18623 2098 18629 2106
rect 18663 2098 18669 2106
rect 18623 2086 18669 2098
rect 18741 2098 18747 2106
rect 18781 2098 18787 2106
rect 18741 2086 18787 2098
rect 18859 2098 18865 2106
rect 18899 2098 18905 2106
rect 18859 2086 18905 2098
rect 18977 2098 18983 2106
rect 19017 2098 19023 2106
rect 18977 2086 19023 2098
rect 19095 2098 19101 2106
rect 19135 2098 19141 2106
rect 19095 2086 19141 2098
rect 19213 2098 19219 2106
rect 19253 2098 19259 2106
rect 19213 2086 19259 2098
rect 19331 2098 19337 2106
rect 19371 2098 19377 2106
rect 19331 2086 19377 2098
rect 19449 2098 19455 2106
rect 19489 2098 19495 2106
rect 19449 2086 19495 2098
rect 19567 2098 19573 2106
rect 19607 2098 19613 2106
rect 19567 2086 19613 2098
rect 19744 2095 20574 2135
rect 20727 2106 20737 2666
rect 20789 2106 20799 2666
rect 20845 2106 20855 2666
rect 20907 2106 20917 2666
rect 20963 2106 20973 2666
rect 21025 2106 21035 2666
rect 21081 2106 21091 2666
rect 21143 2106 21153 2666
rect 21199 2106 21209 2666
rect 21261 2106 21271 2666
rect 21317 2106 21327 2666
rect 21379 2106 21389 2666
rect 21435 2106 21445 2666
rect 21497 2106 21507 2666
rect 21553 2106 21563 2666
rect 21615 2106 21625 2666
rect 21671 2106 21681 2666
rect 21733 2106 21743 2666
rect 21789 2106 21799 2666
rect 21851 2106 21861 2666
rect 21907 2106 21917 2666
rect 21969 2106 21979 2666
rect 22025 2106 22035 2666
rect 22087 2106 22097 2666
rect 22143 2106 22153 2666
rect 22205 2106 22215 2666
rect 22261 2106 22271 2666
rect 22323 2106 22333 2666
rect 22379 2106 22389 2666
rect 22441 2106 22451 2666
rect 22497 2106 22507 2666
rect 22559 2106 22569 2666
rect 22615 2106 22625 2666
rect 22677 2106 22687 2666
rect 22733 2106 22743 2666
rect 22795 2106 22805 2666
rect 22851 2106 22861 2666
rect 22913 2106 22923 2666
rect 22969 2106 22979 2666
rect 23031 2106 23041 2666
rect 23087 2106 23097 2666
rect 23149 2106 23159 2666
rect 23205 2106 23215 2666
rect 23267 2106 23277 2666
rect 23323 2106 23333 2666
rect 23385 2106 23395 2666
rect 23441 2106 23451 2666
rect 23503 2106 23513 2666
rect 23559 2106 23569 2666
rect 23621 2106 23631 2666
rect 23677 2106 23687 2666
rect 23739 2106 23749 2666
rect 23867 2653 23905 2687
rect 23939 2653 23977 2687
rect 24011 2653 24049 2687
rect 24083 2653 24121 2687
rect 24155 2653 24193 2687
rect 24227 2653 24265 2687
rect 24299 2653 24337 2687
rect 24371 2653 24409 2687
rect 24443 2653 24481 2687
rect 24515 2653 24553 2687
rect 24587 2653 24625 2687
rect 24659 2667 25079 2687
rect 24659 2653 25081 2667
rect 23867 2601 23895 2653
rect 23947 2601 23975 2653
rect 24027 2613 24055 2653
rect 24107 2613 24135 2653
rect 24187 2613 24215 2653
rect 24267 2613 24295 2653
rect 24347 2613 24375 2653
rect 24427 2613 24455 2653
rect 24507 2613 24535 2653
rect 24027 2601 24049 2613
rect 24107 2601 24121 2613
rect 24187 2601 24193 2613
rect 24371 2601 24375 2613
rect 24443 2601 24455 2613
rect 24515 2601 24535 2613
rect 24587 2601 24615 2653
rect 24667 2601 24695 2653
rect 24747 2601 24775 2653
rect 24827 2601 24855 2653
rect 24907 2601 24935 2653
rect 24987 2601 25015 2653
rect 25067 2601 25081 2653
rect 23867 2579 23905 2601
rect 23939 2579 23977 2601
rect 24011 2579 24049 2601
rect 24083 2579 24121 2601
rect 24155 2579 24193 2601
rect 24227 2579 24265 2601
rect 24299 2579 24337 2601
rect 24371 2579 24409 2601
rect 24443 2579 24481 2601
rect 24515 2579 24553 2601
rect 24587 2579 24625 2601
rect 24659 2579 25081 2601
rect 23867 2573 25081 2579
rect 23867 2521 23895 2573
rect 23947 2521 23975 2573
rect 24027 2539 24055 2573
rect 24107 2539 24135 2573
rect 24187 2539 24215 2573
rect 24267 2539 24295 2573
rect 24347 2539 24375 2573
rect 24427 2539 24455 2573
rect 24507 2539 24535 2573
rect 24027 2521 24049 2539
rect 24107 2521 24121 2539
rect 24187 2521 24193 2539
rect 24371 2521 24375 2539
rect 24443 2521 24455 2539
rect 24515 2521 24535 2539
rect 24587 2521 24615 2573
rect 24667 2521 24695 2573
rect 24747 2521 24775 2573
rect 24827 2521 24855 2573
rect 24907 2521 24935 2573
rect 24987 2521 25015 2573
rect 25067 2521 25081 2573
rect 23867 2505 23905 2521
rect 23939 2505 23977 2521
rect 24011 2505 24049 2521
rect 24083 2505 24121 2521
rect 24155 2505 24193 2521
rect 24227 2505 24265 2521
rect 24299 2505 24337 2521
rect 24371 2505 24409 2521
rect 24443 2505 24481 2521
rect 24515 2505 24553 2521
rect 24587 2505 24625 2521
rect 24659 2505 25081 2521
rect 23867 2493 25081 2505
rect 23867 2441 23895 2493
rect 23947 2441 23975 2493
rect 24027 2465 24055 2493
rect 24107 2465 24135 2493
rect 24187 2465 24215 2493
rect 24267 2465 24295 2493
rect 24347 2465 24375 2493
rect 24427 2465 24455 2493
rect 24507 2465 24535 2493
rect 24027 2441 24049 2465
rect 24107 2441 24121 2465
rect 24187 2441 24193 2465
rect 24371 2441 24375 2465
rect 24443 2441 24455 2465
rect 24515 2441 24535 2465
rect 24587 2441 24615 2493
rect 24667 2441 24695 2493
rect 24747 2441 24775 2493
rect 24827 2441 24855 2493
rect 24907 2441 24935 2493
rect 24987 2441 25015 2493
rect 25067 2441 25081 2493
rect 23867 2431 23905 2441
rect 23939 2431 23977 2441
rect 24011 2431 24049 2441
rect 24083 2431 24121 2441
rect 24155 2431 24193 2441
rect 24227 2431 24265 2441
rect 24299 2431 24337 2441
rect 24371 2431 24409 2441
rect 24443 2431 24481 2441
rect 24515 2431 24553 2441
rect 24587 2431 24625 2441
rect 24659 2431 25081 2441
rect 23867 2413 25081 2431
rect 23867 2361 23895 2413
rect 23947 2361 23975 2413
rect 24027 2391 24055 2413
rect 24107 2391 24135 2413
rect 24187 2391 24215 2413
rect 24267 2391 24295 2413
rect 24347 2391 24375 2413
rect 24427 2391 24455 2413
rect 24507 2391 24535 2413
rect 24027 2361 24049 2391
rect 24107 2361 24121 2391
rect 24187 2361 24193 2391
rect 24371 2361 24375 2391
rect 24443 2361 24455 2391
rect 24515 2361 24535 2391
rect 24587 2361 24615 2413
rect 24667 2361 24695 2413
rect 24747 2361 24775 2413
rect 24827 2361 24855 2413
rect 24907 2361 24935 2413
rect 24987 2361 25015 2413
rect 25067 2361 25081 2413
rect 23867 2357 23905 2361
rect 23939 2357 23977 2361
rect 24011 2357 24049 2361
rect 24083 2357 24121 2361
rect 24155 2357 24193 2361
rect 24227 2357 24265 2361
rect 24299 2357 24337 2361
rect 24371 2357 24409 2361
rect 24443 2357 24481 2361
rect 24515 2357 24553 2361
rect 24587 2357 24625 2361
rect 24659 2357 25081 2361
rect 23867 2333 25081 2357
rect 23867 2281 23895 2333
rect 23947 2281 23975 2333
rect 24027 2317 24055 2333
rect 24107 2317 24135 2333
rect 24187 2317 24215 2333
rect 24267 2317 24295 2333
rect 24347 2317 24375 2333
rect 24427 2317 24455 2333
rect 24507 2317 24535 2333
rect 24027 2283 24049 2317
rect 24107 2283 24121 2317
rect 24187 2283 24193 2317
rect 24371 2283 24375 2317
rect 24443 2283 24455 2317
rect 24515 2283 24535 2317
rect 24027 2281 24055 2283
rect 24107 2281 24135 2283
rect 24187 2281 24215 2283
rect 24267 2281 24295 2283
rect 24347 2281 24375 2283
rect 24427 2281 24455 2283
rect 24507 2281 24535 2283
rect 24587 2281 24615 2333
rect 24667 2281 24695 2333
rect 24747 2281 24775 2333
rect 24827 2281 24855 2333
rect 24907 2281 24935 2333
rect 24987 2281 25015 2333
rect 25067 2281 25081 2333
rect 23867 2253 25081 2281
rect 23867 2201 23895 2253
rect 23947 2201 23975 2253
rect 24027 2243 24055 2253
rect 24107 2243 24135 2253
rect 24187 2243 24215 2253
rect 24267 2243 24295 2253
rect 24347 2243 24375 2253
rect 24427 2243 24455 2253
rect 24507 2243 24535 2253
rect 24027 2209 24049 2243
rect 24107 2209 24121 2243
rect 24187 2209 24193 2243
rect 24371 2209 24375 2243
rect 24443 2209 24455 2243
rect 24515 2209 24535 2243
rect 24027 2201 24055 2209
rect 24107 2201 24135 2209
rect 24187 2201 24215 2209
rect 24267 2201 24295 2209
rect 24347 2201 24375 2209
rect 24427 2201 24455 2209
rect 24507 2201 24535 2209
rect 24587 2201 24615 2253
rect 24667 2201 24695 2253
rect 24747 2201 24775 2253
rect 24827 2201 24855 2253
rect 24907 2201 24935 2253
rect 24987 2201 25015 2253
rect 25067 2201 25081 2253
rect 23867 2173 25081 2201
rect 23867 2121 23895 2173
rect 23947 2121 23975 2173
rect 24027 2169 24055 2173
rect 24107 2169 24135 2173
rect 24187 2169 24215 2173
rect 24267 2169 24295 2173
rect 24347 2169 24375 2173
rect 24427 2169 24455 2173
rect 24507 2169 24535 2173
rect 24027 2135 24049 2169
rect 24107 2135 24121 2169
rect 24187 2135 24193 2169
rect 24371 2135 24375 2169
rect 24443 2135 24455 2169
rect 24515 2135 24535 2169
rect 24027 2121 24055 2135
rect 24107 2121 24135 2135
rect 24187 2121 24215 2135
rect 24267 2121 24295 2135
rect 24347 2121 24375 2135
rect 24427 2121 24455 2135
rect 24507 2121 24535 2135
rect 24587 2121 24615 2173
rect 24667 2121 24695 2173
rect 24747 2121 24775 2173
rect 24827 2121 24855 2173
rect 24907 2121 24935 2173
rect 24987 2121 25015 2173
rect 25067 2121 25081 2173
rect 4857 2044 4915 2046
rect 4975 2044 5033 2046
rect 5093 2044 5151 2046
rect 5211 2044 5269 2046
rect 5329 2044 5387 2046
rect 5447 2044 5505 2046
rect 5565 2044 5623 2046
rect 5683 2044 5741 2046
rect 5801 2044 5859 2046
rect 5919 2044 5977 2046
rect 6037 2044 6095 2046
rect 6155 2044 6213 2046
rect 6273 2044 6331 2046
rect 6391 2044 6449 2046
rect 6509 2044 6567 2046
rect 7091 2044 7149 2046
rect 7209 2044 7267 2046
rect 7327 2044 7385 2046
rect 7445 2044 7503 2046
rect 7563 2044 7621 2046
rect 7681 2044 7739 2046
rect 7799 2044 7857 2046
rect 7917 2044 7975 2046
rect 8035 2044 8093 2046
rect 8153 2044 8211 2046
rect 8271 2044 8329 2046
rect 8389 2044 8447 2046
rect 8507 2044 8565 2046
rect 8853 2044 8911 2046
rect 8971 2044 9029 2046
rect 9089 2044 9147 2046
rect 9207 2044 9265 2046
rect 9325 2044 9383 2046
rect 9443 2044 9501 2046
rect 9561 2044 9619 2046
rect 9679 2044 9737 2046
rect 9797 2044 9855 2046
rect 9915 2044 9973 2046
rect 10033 2044 10091 2046
rect 10151 2044 10209 2046
rect 10269 2044 10327 2046
rect 10387 2044 10445 2046
rect 10505 2044 10563 2046
rect 4847 1952 4857 2044
rect 4915 1952 4925 2044
rect 4965 1952 4975 2044
rect 5033 1952 5043 2044
rect 5083 1952 5093 2044
rect 5151 1952 5161 2044
rect 5201 1952 5211 2044
rect 5269 1952 5279 2044
rect 5319 1952 5329 2044
rect 5387 1952 5397 2044
rect 5437 1952 5447 2044
rect 5505 1952 5515 2044
rect 5555 1952 5565 2044
rect 5623 1952 5633 2044
rect 5673 1952 5683 2044
rect 5741 1952 5751 2044
rect 5791 1952 5801 2044
rect 5859 1952 5869 2044
rect 5909 1952 5919 2044
rect 5977 1952 5987 2044
rect 6027 1952 6037 2044
rect 6095 1952 6105 2044
rect 6145 1952 6155 2044
rect 6213 1952 6223 2044
rect 6263 1952 6273 2044
rect 6331 1952 6341 2044
rect 6381 1952 6391 2044
rect 6449 1952 6459 2044
rect 6499 1952 6509 2044
rect 6567 1952 6577 2044
rect 6845 1952 6855 2044
rect 6913 1952 6923 2044
rect 6963 1952 6973 2044
rect 7031 1952 7041 2044
rect 7081 1952 7091 2044
rect 7149 1952 7159 2044
rect 7199 1952 7209 2044
rect 7267 1952 7277 2044
rect 7317 1952 7327 2044
rect 7385 1952 7395 2044
rect 7435 1952 7445 2044
rect 7503 1952 7513 2044
rect 7553 1952 7563 2044
rect 7621 1952 7631 2044
rect 7671 1952 7681 2044
rect 7739 1952 7749 2044
rect 7789 1952 7799 2044
rect 7857 1952 7867 2044
rect 7907 1952 7917 2044
rect 7975 1952 7985 2044
rect 8025 1952 8035 2044
rect 8093 1952 8103 2044
rect 8143 1952 8153 2044
rect 8211 1952 8221 2044
rect 8261 1952 8271 2044
rect 8329 1952 8339 2044
rect 8379 1952 8389 2044
rect 8447 1952 8457 2044
rect 8497 1952 8507 2044
rect 8565 1952 8575 2044
rect 8843 1952 8853 2044
rect 8911 1952 8921 2044
rect 8961 1952 8971 2044
rect 9029 1952 9039 2044
rect 9079 1952 9089 2044
rect 9147 1952 9157 2044
rect 9197 1952 9207 2044
rect 9265 1952 9275 2044
rect 9315 1952 9325 2044
rect 9383 1952 9393 2044
rect 9433 1952 9443 2044
rect 9501 1952 9511 2044
rect 9551 1952 9561 2044
rect 9619 1952 9629 2044
rect 9669 1952 9679 2044
rect 9737 1952 9747 2044
rect 9787 1952 9797 2044
rect 9855 1952 9865 2044
rect 9905 1952 9915 2044
rect 9973 1952 9983 2044
rect 10023 1952 10033 2044
rect 10091 1952 10101 2044
rect 10141 1952 10151 2044
rect 10209 1952 10219 2044
rect 10259 1952 10269 2044
rect 10327 1952 10337 2044
rect 10377 1952 10387 2044
rect 10445 1952 10455 2044
rect 10495 1952 10505 2044
rect 10563 1952 10573 2044
rect 12537 1891 12547 2045
rect 12605 1891 12615 2045
rect 12655 1891 12665 2045
rect 12723 1891 12733 2045
rect 12773 1891 12783 2045
rect 12841 1891 12851 2045
rect 12891 1891 12901 2045
rect 12959 1891 12969 2045
rect 13009 1891 13019 2045
rect 13077 1891 13087 2045
rect 13127 1891 13137 2045
rect 13195 1891 13205 2045
rect 13245 1891 13255 2045
rect 13313 1891 13323 2045
rect 13363 1891 13373 2045
rect 13431 1891 13441 2045
rect 13481 1891 13491 2045
rect 13549 1891 13559 2045
rect 13599 1891 13609 2045
rect 13667 1891 13677 2045
rect 13717 1891 13727 2045
rect 13785 1891 13795 2045
rect 13835 1891 13845 2045
rect 13903 1891 13913 2045
rect 13953 1891 13963 2045
rect 14021 1891 14031 2045
rect 14071 1891 14081 2045
rect 14139 1891 14149 2045
rect 14189 1891 14199 2045
rect 14257 1891 14267 2045
rect 14307 1891 14317 2045
rect 14375 1891 14385 2045
rect 14425 1891 14435 2045
rect 14493 1891 14503 2045
rect 14543 1891 14553 2045
rect 14611 1891 14621 2045
rect 14661 1891 14671 2045
rect 14729 1891 14739 2045
rect 14779 1891 14789 2045
rect 14847 1891 14857 2045
rect 14897 1891 14907 2045
rect 14965 1891 14975 2045
rect 15015 1891 15025 2045
rect 15083 1891 15093 2045
rect 15133 1891 15143 2045
rect 15201 1891 15211 2045
rect 15251 1891 15261 2045
rect 15319 1891 15329 2045
rect 15369 1891 15379 2045
rect 15437 1891 15447 2045
rect 15621 2021 16451 2061
rect 19744 2061 19782 2095
rect 19816 2061 19854 2095
rect 19888 2061 19926 2095
rect 19960 2061 19998 2095
rect 20032 2061 20070 2095
rect 20104 2061 20142 2095
rect 20176 2061 20214 2095
rect 20248 2061 20286 2095
rect 20320 2061 20358 2095
rect 20392 2061 20430 2095
rect 20464 2061 20502 2095
rect 20536 2061 20574 2095
rect 20976 2098 20982 2106
rect 21016 2098 21022 2106
rect 20976 2086 21022 2098
rect 21094 2098 21100 2106
rect 21134 2098 21140 2106
rect 21094 2086 21140 2098
rect 21212 2098 21218 2106
rect 21252 2098 21258 2106
rect 21212 2086 21258 2098
rect 21330 2098 21336 2106
rect 21370 2098 21376 2106
rect 21330 2086 21376 2098
rect 21448 2098 21454 2106
rect 21488 2098 21494 2106
rect 21448 2086 21494 2098
rect 21566 2098 21572 2106
rect 21606 2098 21612 2106
rect 21566 2086 21612 2098
rect 21684 2098 21690 2106
rect 21724 2098 21730 2106
rect 21684 2086 21730 2098
rect 21802 2098 21808 2106
rect 21842 2098 21848 2106
rect 21802 2086 21848 2098
rect 21920 2098 21926 2106
rect 21960 2098 21966 2106
rect 21920 2086 21966 2098
rect 22038 2098 22044 2106
rect 22078 2098 22084 2106
rect 22038 2086 22084 2098
rect 22156 2098 22162 2106
rect 22196 2098 22202 2106
rect 22156 2086 22202 2098
rect 22274 2098 22280 2106
rect 22314 2098 22320 2106
rect 22274 2086 22320 2098
rect 22392 2098 22398 2106
rect 22432 2098 22438 2106
rect 22392 2086 22438 2098
rect 22510 2098 22516 2106
rect 22550 2098 22556 2106
rect 22510 2086 22556 2098
rect 22628 2098 22634 2106
rect 22668 2098 22674 2106
rect 22628 2086 22674 2098
rect 22746 2098 22752 2106
rect 22786 2098 22792 2106
rect 22746 2086 22792 2098
rect 22864 2098 22870 2106
rect 22904 2098 22910 2106
rect 22864 2086 22910 2098
rect 22982 2098 22988 2106
rect 23022 2098 23028 2106
rect 22982 2086 23028 2098
rect 23100 2098 23106 2106
rect 23140 2098 23146 2106
rect 23100 2086 23146 2098
rect 23218 2098 23224 2106
rect 23258 2098 23264 2106
rect 23218 2086 23264 2098
rect 23336 2098 23342 2106
rect 23376 2098 23382 2106
rect 23336 2086 23382 2098
rect 23454 2098 23460 2106
rect 23494 2098 23500 2106
rect 23454 2086 23500 2098
rect 23572 2098 23578 2106
rect 23612 2098 23618 2106
rect 23572 2086 23618 2098
rect 23690 2098 23696 2106
rect 23730 2098 23736 2106
rect 23690 2086 23736 2098
rect 23867 2095 25081 2121
rect 23867 2093 23905 2095
rect 23939 2093 23977 2095
rect 24011 2093 24049 2095
rect 24083 2093 24121 2095
rect 24155 2093 24193 2095
rect 24227 2093 24265 2095
rect 24299 2093 24337 2095
rect 24371 2093 24409 2095
rect 24443 2093 24481 2095
rect 24515 2093 24553 2095
rect 24587 2093 24625 2095
rect 24659 2093 25081 2095
rect 15621 1987 15659 2021
rect 15693 1987 15731 2021
rect 15765 1987 15803 2021
rect 15837 1987 15875 2021
rect 15909 1987 15947 2021
rect 15981 1987 16019 2021
rect 16053 1987 16091 2021
rect 16125 1987 16163 2021
rect 16197 1987 16235 2021
rect 16269 1987 16307 2021
rect 16341 1987 16379 2021
rect 16413 1987 16451 2021
rect 15621 1947 16451 1987
rect 15621 1913 15659 1947
rect 15693 1913 15731 1947
rect 15765 1913 15803 1947
rect 15837 1913 15875 1947
rect 15909 1913 15947 1947
rect 15981 1913 16019 1947
rect 16053 1913 16091 1947
rect 16125 1913 16163 1947
rect 16197 1913 16235 1947
rect 16269 1913 16307 1947
rect 16341 1913 16379 1947
rect 16413 1913 16451 1947
rect 15621 1873 16451 1913
rect 16660 1891 16670 2045
rect 16728 1891 16738 2045
rect 16778 1891 16788 2045
rect 16846 1891 16856 2045
rect 16896 1891 16906 2045
rect 16964 1891 16974 2045
rect 17014 1891 17024 2045
rect 17082 1891 17092 2045
rect 17132 1891 17142 2045
rect 17200 1891 17210 2045
rect 17250 1891 17260 2045
rect 17318 1891 17328 2045
rect 17368 1891 17378 2045
rect 17436 1891 17446 2045
rect 17486 1891 17496 2045
rect 17554 1891 17564 2045
rect 17604 1891 17614 2045
rect 17672 1891 17682 2045
rect 17722 1891 17732 2045
rect 17790 1891 17800 2045
rect 17840 1891 17850 2045
rect 17908 1891 17918 2045
rect 17958 1891 17968 2045
rect 18026 1891 18036 2045
rect 18076 1891 18086 2045
rect 18144 1891 18154 2045
rect 18194 1891 18204 2045
rect 18262 1891 18272 2045
rect 18312 1891 18322 2045
rect 18380 1891 18390 2045
rect 18430 1891 18440 2045
rect 18498 1891 18508 2045
rect 18548 1891 18558 2045
rect 18616 1891 18626 2045
rect 18666 1891 18676 2045
rect 18734 1891 18744 2045
rect 18784 1891 18794 2045
rect 18852 1891 18862 2045
rect 18902 1891 18912 2045
rect 18970 1891 18980 2045
rect 19020 1891 19030 2045
rect 19088 1891 19098 2045
rect 19138 1891 19148 2045
rect 19206 1891 19216 2045
rect 19256 1891 19266 2045
rect 19324 1891 19334 2045
rect 19374 1891 19384 2045
rect 19442 1891 19452 2045
rect 19492 1891 19502 2045
rect 19560 1891 19570 2045
rect 19744 2021 20574 2061
rect 19744 1987 19782 2021
rect 19816 1987 19854 2021
rect 19888 1987 19926 2021
rect 19960 1987 19998 2021
rect 20032 1987 20070 2021
rect 20104 1987 20142 2021
rect 20176 1987 20214 2021
rect 20248 1987 20286 2021
rect 20320 1987 20358 2021
rect 20392 1987 20430 2021
rect 20464 1987 20502 2021
rect 20536 1987 20574 2021
rect 19744 1947 20574 1987
rect 19744 1913 19782 1947
rect 19816 1913 19854 1947
rect 19888 1913 19926 1947
rect 19960 1913 19998 1947
rect 20032 1913 20070 1947
rect 20104 1913 20142 1947
rect 20176 1913 20214 1947
rect 20248 1913 20286 1947
rect 20320 1913 20358 1947
rect 20392 1913 20430 1947
rect 20464 1913 20502 1947
rect 20536 1913 20574 1947
rect 12494 1838 12540 1850
rect 12494 1830 12500 1838
rect 12534 1830 12540 1838
rect 12612 1838 12658 1850
rect 12612 1830 12618 1838
rect 12652 1830 12658 1838
rect 12730 1838 12776 1850
rect 12730 1830 12736 1838
rect 12770 1830 12776 1838
rect 12848 1838 12894 1850
rect 12848 1830 12854 1838
rect 12888 1830 12894 1838
rect 12966 1838 13012 1850
rect 12966 1830 12972 1838
rect 13006 1830 13012 1838
rect 13084 1838 13130 1850
rect 13084 1830 13090 1838
rect 13124 1830 13130 1838
rect 13202 1838 13248 1850
rect 13202 1830 13208 1838
rect 13242 1830 13248 1838
rect 13320 1838 13366 1850
rect 13320 1830 13326 1838
rect 13360 1830 13366 1838
rect 13438 1838 13484 1850
rect 13438 1830 13444 1838
rect 13478 1830 13484 1838
rect 13556 1838 13602 1850
rect 13556 1830 13562 1838
rect 13596 1830 13602 1838
rect 13674 1838 13720 1850
rect 13674 1830 13680 1838
rect 13714 1830 13720 1838
rect 13792 1838 13838 1850
rect 13792 1830 13798 1838
rect 13832 1830 13838 1838
rect 13910 1838 13956 1850
rect 13910 1830 13916 1838
rect 13950 1830 13956 1838
rect 14028 1838 14074 1850
rect 14028 1830 14034 1838
rect 14068 1830 14074 1838
rect 14146 1838 14192 1850
rect 14146 1830 14152 1838
rect 14186 1830 14192 1838
rect 14264 1838 14310 1850
rect 14264 1830 14270 1838
rect 14304 1830 14310 1838
rect 14382 1838 14428 1850
rect 14382 1830 14388 1838
rect 14422 1830 14428 1838
rect 14500 1838 14546 1850
rect 14500 1830 14506 1838
rect 14540 1830 14546 1838
rect 14618 1838 14664 1850
rect 14618 1830 14624 1838
rect 14658 1830 14664 1838
rect 14736 1838 14782 1850
rect 14736 1830 14742 1838
rect 14776 1830 14782 1838
rect 14854 1838 14900 1850
rect 14854 1830 14860 1838
rect 14894 1830 14900 1838
rect 14972 1838 15018 1850
rect 14972 1830 14978 1838
rect 15012 1830 15018 1838
rect 15090 1838 15136 1850
rect 15090 1830 15096 1838
rect 15130 1830 15136 1838
rect 15208 1838 15254 1850
rect 15208 1830 15214 1838
rect 15248 1830 15254 1838
rect 15326 1838 15372 1850
rect 15326 1830 15332 1838
rect 15366 1830 15372 1838
rect 15444 1838 15490 1850
rect 15444 1830 15450 1838
rect 15484 1830 15490 1838
rect 15621 1839 15659 1873
rect 15693 1839 15731 1873
rect 15765 1839 15803 1873
rect 15837 1839 15875 1873
rect 15909 1839 15947 1873
rect 15981 1839 16019 1873
rect 16053 1839 16091 1873
rect 16125 1839 16163 1873
rect 16197 1839 16235 1873
rect 16269 1839 16307 1873
rect 16341 1839 16379 1873
rect 16413 1839 16451 1873
rect 19744 1873 20574 1913
rect 20783 1891 20793 2045
rect 20851 1891 20861 2045
rect 20901 1891 20911 2045
rect 20969 1891 20979 2045
rect 21019 1891 21029 2045
rect 21087 1891 21097 2045
rect 21137 1891 21147 2045
rect 21205 1891 21215 2045
rect 21255 1891 21265 2045
rect 21323 1891 21333 2045
rect 21373 1891 21383 2045
rect 21441 1891 21451 2045
rect 21491 1891 21501 2045
rect 21559 1891 21569 2045
rect 21609 1891 21619 2045
rect 21677 1891 21687 2045
rect 21727 1891 21737 2045
rect 21795 1891 21805 2045
rect 21845 1891 21855 2045
rect 21913 1891 21923 2045
rect 21963 1891 21973 2045
rect 22031 1891 22041 2045
rect 22081 1891 22091 2045
rect 22149 1891 22159 2045
rect 22199 1891 22209 2045
rect 22267 1891 22277 2045
rect 22317 1891 22327 2045
rect 22385 1891 22395 2045
rect 22435 1891 22445 2045
rect 22503 1891 22513 2045
rect 22553 1891 22563 2045
rect 22621 1891 22631 2045
rect 22671 1891 22681 2045
rect 22739 1891 22749 2045
rect 22789 1891 22799 2045
rect 22857 1891 22867 2045
rect 22907 1891 22917 2045
rect 22975 1891 22985 2045
rect 23025 1891 23035 2045
rect 23093 1891 23103 2045
rect 23143 1891 23153 2045
rect 23211 1891 23221 2045
rect 23261 1891 23271 2045
rect 23329 1891 23339 2045
rect 23379 1891 23389 2045
rect 23447 1891 23457 2045
rect 23497 1891 23507 2045
rect 23565 1891 23575 2045
rect 23615 1891 23625 2045
rect 23683 1891 23693 2045
rect 23867 2041 23895 2093
rect 23947 2041 23975 2093
rect 24027 2061 24049 2093
rect 24107 2061 24121 2093
rect 24187 2061 24193 2093
rect 24371 2061 24375 2093
rect 24443 2061 24455 2093
rect 24515 2061 24535 2093
rect 24027 2041 24055 2061
rect 24107 2041 24135 2061
rect 24187 2041 24215 2061
rect 24267 2041 24295 2061
rect 24347 2041 24375 2061
rect 24427 2041 24455 2061
rect 24507 2041 24535 2061
rect 24587 2041 24615 2093
rect 24667 2041 24695 2093
rect 24747 2041 24775 2093
rect 24827 2041 24855 2093
rect 24907 2041 24935 2093
rect 24987 2041 25015 2093
rect 25067 2041 25081 2093
rect 23867 2021 25081 2041
rect 23867 2013 23905 2021
rect 23939 2013 23977 2021
rect 24011 2013 24049 2021
rect 24083 2013 24121 2021
rect 24155 2013 24193 2021
rect 24227 2013 24265 2021
rect 24299 2013 24337 2021
rect 24371 2013 24409 2021
rect 24443 2013 24481 2021
rect 24515 2013 24553 2021
rect 24587 2013 24625 2021
rect 24659 2013 25081 2021
rect 23867 1961 23895 2013
rect 23947 1961 23975 2013
rect 24027 1987 24049 2013
rect 24107 1987 24121 2013
rect 24187 1987 24193 2013
rect 24371 1987 24375 2013
rect 24443 1987 24455 2013
rect 24515 1987 24535 2013
rect 24027 1961 24055 1987
rect 24107 1961 24135 1987
rect 24187 1961 24215 1987
rect 24267 1961 24295 1987
rect 24347 1961 24375 1987
rect 24427 1961 24455 1987
rect 24507 1961 24535 1987
rect 24587 1961 24615 2013
rect 24667 1961 24695 2013
rect 24747 1961 24775 2013
rect 24827 1961 24855 2013
rect 24907 1961 24935 2013
rect 24987 1961 25015 2013
rect 25067 1961 25081 2013
rect 23867 1947 25081 1961
rect 23867 1933 23905 1947
rect 23939 1933 23977 1947
rect 24011 1933 24049 1947
rect 24083 1933 24121 1947
rect 24155 1933 24193 1947
rect 24227 1933 24265 1947
rect 24299 1933 24337 1947
rect 24371 1933 24409 1947
rect 24443 1933 24481 1947
rect 24515 1933 24553 1947
rect 24587 1933 24625 1947
rect 24659 1933 25081 1947
rect 4582 -6438 4611 1770
rect 4634 -6438 4698 1770
rect 4722 1495 4794 1570
rect 4722 1319 4801 1495
rect 4853 1393 5037 1499
rect 4853 1319 4863 1393
rect 5089 1393 5273 1495
rect 5325 1393 5509 1495
rect 5561 1393 5745 1495
rect 5797 1393 5981 1495
rect 6033 1393 6217 1495
rect 6269 1393 6453 1495
rect 6505 1393 6689 1495
rect 6741 1393 6925 1495
rect 6977 1393 7161 1495
rect 7213 1393 7397 1495
rect 7449 1393 7633 1495
rect 7685 1393 7869 1495
rect 7921 1393 8105 1495
rect 8157 1393 8341 1495
rect 8393 1393 8577 1495
rect 8629 1393 8813 1500
rect 8865 1393 9049 1504
rect 9101 1393 9285 1505
rect 9337 1393 9521 1504
rect 9573 1393 9757 1505
rect 9809 1393 9993 1504
rect 10045 1393 10229 1495
rect 10281 1393 10465 1495
rect 10517 1393 10701 1495
rect 10753 1393 10808 1495
rect 12481 1270 12491 1830
rect 12543 1270 12553 1830
rect 12599 1270 12609 1830
rect 12661 1270 12671 1830
rect 12717 1270 12727 1830
rect 12779 1270 12789 1830
rect 12835 1270 12845 1830
rect 12897 1270 12907 1830
rect 12953 1270 12963 1830
rect 13015 1270 13025 1830
rect 13071 1270 13081 1830
rect 13133 1270 13143 1830
rect 13189 1270 13199 1830
rect 13251 1270 13261 1830
rect 13307 1270 13317 1830
rect 13369 1270 13379 1830
rect 13425 1270 13435 1830
rect 13487 1270 13497 1830
rect 13543 1270 13553 1830
rect 13605 1270 13615 1830
rect 13661 1270 13671 1830
rect 13723 1270 13733 1830
rect 13779 1270 13789 1830
rect 13841 1270 13851 1830
rect 13897 1270 13907 1830
rect 13959 1270 13969 1830
rect 14015 1270 14025 1830
rect 14077 1270 14087 1830
rect 14133 1270 14143 1830
rect 14195 1270 14205 1830
rect 14251 1270 14261 1830
rect 14313 1270 14323 1830
rect 14369 1270 14379 1830
rect 14431 1270 14441 1830
rect 14487 1270 14497 1830
rect 14549 1270 14559 1830
rect 14605 1270 14615 1830
rect 14667 1270 14677 1830
rect 14723 1270 14733 1830
rect 14785 1270 14795 1830
rect 14841 1270 14851 1830
rect 14903 1270 14913 1830
rect 14959 1270 14969 1830
rect 15021 1270 15031 1830
rect 15077 1270 15087 1830
rect 15139 1270 15149 1830
rect 15195 1270 15205 1830
rect 15257 1270 15267 1830
rect 15313 1270 15323 1830
rect 15375 1270 15385 1830
rect 15431 1270 15441 1830
rect 15493 1270 15503 1830
rect 15621 1799 16451 1839
rect 16617 1838 16663 1850
rect 16617 1830 16623 1838
rect 16657 1830 16663 1838
rect 16735 1838 16781 1850
rect 16735 1830 16741 1838
rect 16775 1830 16781 1838
rect 16853 1838 16899 1850
rect 16853 1830 16859 1838
rect 16893 1830 16899 1838
rect 16971 1838 17017 1850
rect 16971 1830 16977 1838
rect 17011 1830 17017 1838
rect 17089 1838 17135 1850
rect 17089 1830 17095 1838
rect 17129 1830 17135 1838
rect 17207 1838 17253 1850
rect 17207 1830 17213 1838
rect 17247 1830 17253 1838
rect 17325 1838 17371 1850
rect 17325 1830 17331 1838
rect 17365 1830 17371 1838
rect 17443 1838 17489 1850
rect 17443 1830 17449 1838
rect 17483 1830 17489 1838
rect 17561 1838 17607 1850
rect 17561 1830 17567 1838
rect 17601 1830 17607 1838
rect 17679 1838 17725 1850
rect 17679 1830 17685 1838
rect 17719 1830 17725 1838
rect 17797 1838 17843 1850
rect 17797 1830 17803 1838
rect 17837 1830 17843 1838
rect 17915 1838 17961 1850
rect 17915 1830 17921 1838
rect 17955 1830 17961 1838
rect 18033 1838 18079 1850
rect 18033 1830 18039 1838
rect 18073 1830 18079 1838
rect 18151 1838 18197 1850
rect 18151 1830 18157 1838
rect 18191 1830 18197 1838
rect 18269 1838 18315 1850
rect 18269 1830 18275 1838
rect 18309 1830 18315 1838
rect 18387 1838 18433 1850
rect 18387 1830 18393 1838
rect 18427 1830 18433 1838
rect 18505 1838 18551 1850
rect 18505 1830 18511 1838
rect 18545 1830 18551 1838
rect 18623 1838 18669 1850
rect 18623 1830 18629 1838
rect 18663 1830 18669 1838
rect 18741 1838 18787 1850
rect 18741 1830 18747 1838
rect 18781 1830 18787 1838
rect 18859 1838 18905 1850
rect 18859 1830 18865 1838
rect 18899 1830 18905 1838
rect 18977 1838 19023 1850
rect 18977 1830 18983 1838
rect 19017 1830 19023 1838
rect 19095 1838 19141 1850
rect 19095 1830 19101 1838
rect 19135 1830 19141 1838
rect 19213 1838 19259 1850
rect 19213 1830 19219 1838
rect 19253 1830 19259 1838
rect 19331 1838 19377 1850
rect 19331 1830 19337 1838
rect 19371 1830 19377 1838
rect 19449 1838 19495 1850
rect 19449 1830 19455 1838
rect 19489 1830 19495 1838
rect 19567 1838 19613 1850
rect 19567 1830 19573 1838
rect 19607 1830 19613 1838
rect 19744 1839 19782 1873
rect 19816 1839 19854 1873
rect 19888 1839 19926 1873
rect 19960 1839 19998 1873
rect 20032 1839 20070 1873
rect 20104 1839 20142 1873
rect 20176 1839 20214 1873
rect 20248 1839 20286 1873
rect 20320 1839 20358 1873
rect 20392 1839 20430 1873
rect 20464 1839 20502 1873
rect 20536 1839 20574 1873
rect 23867 1881 23895 1933
rect 23947 1881 23975 1933
rect 24027 1913 24049 1933
rect 24107 1913 24121 1933
rect 24187 1913 24193 1933
rect 24371 1913 24375 1933
rect 24443 1913 24455 1933
rect 24515 1913 24535 1933
rect 24027 1881 24055 1913
rect 24107 1881 24135 1913
rect 24187 1881 24215 1913
rect 24267 1881 24295 1913
rect 24347 1881 24375 1913
rect 24427 1881 24455 1913
rect 24507 1881 24535 1913
rect 24587 1881 24615 1933
rect 24667 1881 24695 1933
rect 24747 1881 24775 1933
rect 24827 1881 24855 1933
rect 24907 1881 24935 1933
rect 24987 1881 25015 1933
rect 25067 1881 25081 1933
rect 23867 1873 25081 1881
rect 23867 1853 23905 1873
rect 23939 1853 23977 1873
rect 24011 1853 24049 1873
rect 24083 1853 24121 1873
rect 24155 1853 24193 1873
rect 24227 1853 24265 1873
rect 24299 1853 24337 1873
rect 24371 1853 24409 1873
rect 24443 1853 24481 1873
rect 24515 1853 24553 1873
rect 24587 1853 24625 1873
rect 24659 1853 25081 1873
rect 15621 1765 15659 1799
rect 15693 1765 15731 1799
rect 15765 1765 15803 1799
rect 15837 1765 15875 1799
rect 15909 1765 15947 1799
rect 15981 1765 16019 1799
rect 16053 1765 16091 1799
rect 16125 1765 16163 1799
rect 16197 1765 16235 1799
rect 16269 1765 16307 1799
rect 16341 1765 16379 1799
rect 16413 1765 16451 1799
rect 15621 1725 16451 1765
rect 15621 1691 15659 1725
rect 15693 1691 15731 1725
rect 15765 1691 15803 1725
rect 15837 1691 15875 1725
rect 15909 1691 15947 1725
rect 15981 1691 16019 1725
rect 16053 1691 16091 1725
rect 16125 1691 16163 1725
rect 16197 1691 16235 1725
rect 16269 1691 16307 1725
rect 16341 1691 16379 1725
rect 16413 1691 16451 1725
rect 15621 1651 16451 1691
rect 15621 1617 15659 1651
rect 15693 1617 15731 1651
rect 15765 1617 15803 1651
rect 15837 1617 15875 1651
rect 15909 1617 15947 1651
rect 15981 1617 16019 1651
rect 16053 1617 16091 1651
rect 16125 1617 16163 1651
rect 16197 1617 16235 1651
rect 16269 1617 16307 1651
rect 16341 1617 16379 1651
rect 16413 1617 16451 1651
rect 15621 1577 16451 1617
rect 15621 1543 15659 1577
rect 15693 1543 15731 1577
rect 15765 1543 15803 1577
rect 15837 1543 15875 1577
rect 15909 1543 15947 1577
rect 15981 1543 16019 1577
rect 16053 1543 16091 1577
rect 16125 1543 16163 1577
rect 16197 1543 16235 1577
rect 16269 1543 16307 1577
rect 16341 1543 16379 1577
rect 16413 1543 16451 1577
rect 15621 1503 16451 1543
rect 15621 1469 15659 1503
rect 15693 1469 15731 1503
rect 15765 1469 15803 1503
rect 15837 1469 15875 1503
rect 15909 1469 15947 1503
rect 15981 1469 16019 1503
rect 16053 1469 16091 1503
rect 16125 1469 16163 1503
rect 16197 1469 16235 1503
rect 16269 1469 16307 1503
rect 16341 1469 16379 1503
rect 16413 1469 16451 1503
rect 15621 1429 16451 1469
rect 15621 1395 15659 1429
rect 15693 1395 15731 1429
rect 15765 1395 15803 1429
rect 15837 1395 15875 1429
rect 15909 1395 15947 1429
rect 15981 1395 16019 1429
rect 16053 1395 16091 1429
rect 16125 1395 16163 1429
rect 16197 1395 16235 1429
rect 16269 1395 16307 1429
rect 16341 1395 16379 1429
rect 16413 1395 16451 1429
rect 15621 1375 16451 1395
rect 15619 1355 16452 1375
rect 15619 1321 15659 1355
rect 15693 1321 15731 1355
rect 15765 1321 15803 1355
rect 15837 1321 15875 1355
rect 15909 1321 15947 1355
rect 15981 1321 16019 1355
rect 16053 1321 16091 1355
rect 16125 1321 16163 1355
rect 16197 1321 16235 1355
rect 16269 1321 16307 1355
rect 16341 1321 16379 1355
rect 16413 1321 16452 1355
rect 15619 1281 16452 1321
rect 12494 1262 12500 1270
rect 12534 1262 12540 1270
rect 12494 1250 12540 1262
rect 12612 1262 12618 1270
rect 12652 1262 12658 1270
rect 12612 1250 12658 1262
rect 12730 1262 12736 1270
rect 12770 1262 12776 1270
rect 12730 1250 12776 1262
rect 12848 1262 12854 1270
rect 12888 1262 12894 1270
rect 12848 1250 12894 1262
rect 12966 1262 12972 1270
rect 13006 1262 13012 1270
rect 12966 1250 13012 1262
rect 13084 1262 13090 1270
rect 13124 1262 13130 1270
rect 13084 1250 13130 1262
rect 13202 1262 13208 1270
rect 13242 1262 13248 1270
rect 13202 1250 13248 1262
rect 13320 1262 13326 1270
rect 13360 1262 13366 1270
rect 13320 1250 13366 1262
rect 13438 1262 13444 1270
rect 13478 1262 13484 1270
rect 13438 1250 13484 1262
rect 13556 1262 13562 1270
rect 13596 1262 13602 1270
rect 13556 1250 13602 1262
rect 13674 1262 13680 1270
rect 13714 1262 13720 1270
rect 13674 1250 13720 1262
rect 13792 1262 13798 1270
rect 13832 1262 13838 1270
rect 13792 1250 13838 1262
rect 13910 1262 13916 1270
rect 13950 1262 13956 1270
rect 13910 1250 13956 1262
rect 14028 1262 14034 1270
rect 14068 1262 14074 1270
rect 14028 1250 14074 1262
rect 14146 1262 14152 1270
rect 14186 1262 14192 1270
rect 14146 1250 14192 1262
rect 14264 1262 14270 1270
rect 14304 1262 14310 1270
rect 14264 1250 14310 1262
rect 14382 1262 14388 1270
rect 14422 1262 14428 1270
rect 14382 1250 14428 1262
rect 14500 1262 14506 1270
rect 14540 1262 14546 1270
rect 14500 1250 14546 1262
rect 14618 1262 14624 1270
rect 14658 1262 14664 1270
rect 14618 1250 14664 1262
rect 14736 1262 14742 1270
rect 14776 1262 14782 1270
rect 14736 1250 14782 1262
rect 14854 1262 14860 1270
rect 14894 1262 14900 1270
rect 14854 1250 14900 1262
rect 14972 1262 14978 1270
rect 15012 1262 15018 1270
rect 14972 1250 15018 1262
rect 15090 1262 15096 1270
rect 15130 1262 15136 1270
rect 15090 1250 15136 1262
rect 15208 1262 15214 1270
rect 15248 1262 15254 1270
rect 15208 1250 15254 1262
rect 15326 1262 15332 1270
rect 15366 1262 15372 1270
rect 15326 1250 15372 1262
rect 15444 1262 15450 1270
rect 15484 1262 15490 1270
rect 15444 1250 15490 1262
rect 15619 1247 15659 1281
rect 15693 1247 15731 1281
rect 15765 1247 15803 1281
rect 15837 1247 15875 1281
rect 15909 1247 15947 1281
rect 15981 1247 16019 1281
rect 16053 1247 16091 1281
rect 16125 1247 16163 1281
rect 16197 1247 16235 1281
rect 16269 1247 16307 1281
rect 16341 1247 16379 1281
rect 16413 1247 16452 1281
rect 16604 1270 16614 1830
rect 16666 1270 16676 1830
rect 16722 1270 16732 1830
rect 16784 1270 16794 1830
rect 16840 1270 16850 1830
rect 16902 1270 16912 1830
rect 16958 1270 16968 1830
rect 17020 1270 17030 1830
rect 17076 1270 17086 1830
rect 17138 1270 17148 1830
rect 17194 1270 17204 1830
rect 17256 1270 17266 1830
rect 17312 1270 17322 1830
rect 17374 1270 17384 1830
rect 17430 1270 17440 1830
rect 17492 1270 17502 1830
rect 17548 1270 17558 1830
rect 17610 1270 17620 1830
rect 17666 1270 17676 1830
rect 17728 1270 17738 1830
rect 17784 1270 17794 1830
rect 17846 1270 17856 1830
rect 17902 1270 17912 1830
rect 17964 1270 17974 1830
rect 18020 1270 18030 1830
rect 18082 1270 18092 1830
rect 18138 1270 18148 1830
rect 18200 1270 18210 1830
rect 18256 1270 18266 1830
rect 18318 1270 18328 1830
rect 18374 1270 18384 1830
rect 18436 1270 18446 1830
rect 18492 1270 18502 1830
rect 18554 1270 18564 1830
rect 18610 1270 18620 1830
rect 18672 1270 18682 1830
rect 18728 1270 18738 1830
rect 18790 1270 18800 1830
rect 18846 1270 18856 1830
rect 18908 1270 18918 1830
rect 18964 1270 18974 1830
rect 19026 1270 19036 1830
rect 19082 1270 19092 1830
rect 19144 1270 19154 1830
rect 19200 1270 19210 1830
rect 19262 1270 19272 1830
rect 19318 1270 19328 1830
rect 19380 1270 19390 1830
rect 19436 1270 19446 1830
rect 19498 1270 19508 1830
rect 19554 1270 19564 1830
rect 19616 1270 19626 1830
rect 19744 1799 20574 1839
rect 20740 1838 20786 1850
rect 20740 1830 20746 1838
rect 20780 1830 20786 1838
rect 20858 1838 20904 1850
rect 20858 1830 20864 1838
rect 20898 1830 20904 1838
rect 20976 1838 21022 1850
rect 20976 1830 20982 1838
rect 21016 1830 21022 1838
rect 21094 1838 21140 1850
rect 21094 1830 21100 1838
rect 21134 1830 21140 1838
rect 21212 1838 21258 1850
rect 21212 1830 21218 1838
rect 21252 1830 21258 1838
rect 21330 1838 21376 1850
rect 21330 1830 21336 1838
rect 21370 1830 21376 1838
rect 21448 1838 21494 1850
rect 21448 1830 21454 1838
rect 21488 1830 21494 1838
rect 21566 1838 21612 1850
rect 21566 1830 21572 1838
rect 21606 1830 21612 1838
rect 21684 1838 21730 1850
rect 21684 1830 21690 1838
rect 21724 1830 21730 1838
rect 21802 1838 21848 1850
rect 21802 1830 21808 1838
rect 21842 1830 21848 1838
rect 21920 1838 21966 1850
rect 21920 1830 21926 1838
rect 21960 1830 21966 1838
rect 22038 1838 22084 1850
rect 22038 1830 22044 1838
rect 22078 1830 22084 1838
rect 22156 1838 22202 1850
rect 22156 1830 22162 1838
rect 22196 1830 22202 1838
rect 22274 1838 22320 1850
rect 22274 1830 22280 1838
rect 22314 1830 22320 1838
rect 22392 1838 22438 1850
rect 22392 1830 22398 1838
rect 22432 1830 22438 1838
rect 22510 1838 22556 1850
rect 22510 1830 22516 1838
rect 22550 1830 22556 1838
rect 22628 1838 22674 1850
rect 22628 1830 22634 1838
rect 22668 1830 22674 1838
rect 22746 1838 22792 1850
rect 22746 1830 22752 1838
rect 22786 1830 22792 1838
rect 22864 1838 22910 1850
rect 22864 1830 22870 1838
rect 22904 1830 22910 1838
rect 22982 1838 23028 1850
rect 22982 1830 22988 1838
rect 23022 1830 23028 1838
rect 23100 1838 23146 1850
rect 23100 1830 23106 1838
rect 23140 1830 23146 1838
rect 23218 1838 23264 1850
rect 23218 1830 23224 1838
rect 23258 1830 23264 1838
rect 23336 1838 23382 1850
rect 23336 1830 23342 1838
rect 23376 1830 23382 1838
rect 23454 1838 23500 1850
rect 23454 1830 23460 1838
rect 23494 1830 23500 1838
rect 23572 1838 23618 1850
rect 23572 1830 23578 1838
rect 23612 1830 23618 1838
rect 23690 1838 23736 1850
rect 23690 1830 23696 1838
rect 23730 1830 23736 1838
rect 19744 1765 19782 1799
rect 19816 1765 19854 1799
rect 19888 1765 19926 1799
rect 19960 1765 19998 1799
rect 20032 1765 20070 1799
rect 20104 1765 20142 1799
rect 20176 1765 20214 1799
rect 20248 1765 20286 1799
rect 20320 1765 20358 1799
rect 20392 1765 20430 1799
rect 20464 1765 20502 1799
rect 20536 1765 20574 1799
rect 19744 1725 20574 1765
rect 19744 1691 19782 1725
rect 19816 1691 19854 1725
rect 19888 1691 19926 1725
rect 19960 1691 19998 1725
rect 20032 1691 20070 1725
rect 20104 1691 20142 1725
rect 20176 1691 20214 1725
rect 20248 1691 20286 1725
rect 20320 1691 20358 1725
rect 20392 1691 20430 1725
rect 20464 1691 20502 1725
rect 20536 1691 20574 1725
rect 19744 1651 20574 1691
rect 19744 1617 19782 1651
rect 19816 1617 19854 1651
rect 19888 1617 19926 1651
rect 19960 1617 19998 1651
rect 20032 1617 20070 1651
rect 20104 1617 20142 1651
rect 20176 1617 20214 1651
rect 20248 1617 20286 1651
rect 20320 1617 20358 1651
rect 20392 1617 20430 1651
rect 20464 1617 20502 1651
rect 20536 1617 20574 1651
rect 19744 1577 20574 1617
rect 19744 1543 19782 1577
rect 19816 1543 19854 1577
rect 19888 1543 19926 1577
rect 19960 1543 19998 1577
rect 20032 1543 20070 1577
rect 20104 1543 20142 1577
rect 20176 1543 20214 1577
rect 20248 1543 20286 1577
rect 20320 1543 20358 1577
rect 20392 1543 20430 1577
rect 20464 1543 20502 1577
rect 20536 1543 20574 1577
rect 19744 1503 20574 1543
rect 19744 1469 19782 1503
rect 19816 1469 19854 1503
rect 19888 1469 19926 1503
rect 19960 1469 19998 1503
rect 20032 1469 20070 1503
rect 20104 1469 20142 1503
rect 20176 1469 20214 1503
rect 20248 1469 20286 1503
rect 20320 1469 20358 1503
rect 20392 1469 20430 1503
rect 20464 1469 20502 1503
rect 20536 1469 20574 1503
rect 19744 1429 20574 1469
rect 19744 1395 19782 1429
rect 19816 1395 19854 1429
rect 19888 1395 19926 1429
rect 19960 1395 19998 1429
rect 20032 1395 20070 1429
rect 20104 1395 20142 1429
rect 20176 1395 20214 1429
rect 20248 1395 20286 1429
rect 20320 1395 20358 1429
rect 20392 1395 20430 1429
rect 20464 1395 20502 1429
rect 20536 1395 20574 1429
rect 19744 1355 20574 1395
rect 19744 1330 19782 1355
rect 19743 1321 19782 1330
rect 19816 1321 19854 1355
rect 19888 1321 19926 1355
rect 19960 1321 19998 1355
rect 20032 1321 20070 1355
rect 20104 1321 20142 1355
rect 20176 1321 20214 1355
rect 20248 1321 20286 1355
rect 20320 1321 20358 1355
rect 20392 1321 20430 1355
rect 20464 1321 20502 1355
rect 20536 1330 20574 1355
rect 20536 1321 20575 1330
rect 19743 1281 20575 1321
rect 16617 1262 16623 1270
rect 16657 1262 16663 1270
rect 16617 1250 16663 1262
rect 16735 1262 16741 1270
rect 16775 1262 16781 1270
rect 16735 1250 16781 1262
rect 16853 1262 16859 1270
rect 16893 1262 16899 1270
rect 16853 1250 16899 1262
rect 16971 1262 16977 1270
rect 17011 1262 17017 1270
rect 16971 1250 17017 1262
rect 17089 1262 17095 1270
rect 17129 1262 17135 1270
rect 17089 1250 17135 1262
rect 17207 1262 17213 1270
rect 17247 1262 17253 1270
rect 17207 1250 17253 1262
rect 17325 1262 17331 1270
rect 17365 1262 17371 1270
rect 17325 1250 17371 1262
rect 17443 1262 17449 1270
rect 17483 1262 17489 1270
rect 17443 1250 17489 1262
rect 17561 1262 17567 1270
rect 17601 1262 17607 1270
rect 17561 1250 17607 1262
rect 17679 1262 17685 1270
rect 17719 1262 17725 1270
rect 17679 1250 17725 1262
rect 17797 1262 17803 1270
rect 17837 1262 17843 1270
rect 17797 1250 17843 1262
rect 17915 1262 17921 1270
rect 17955 1262 17961 1270
rect 17915 1250 17961 1262
rect 18033 1262 18039 1270
rect 18073 1262 18079 1270
rect 18033 1250 18079 1262
rect 18151 1262 18157 1270
rect 18191 1262 18197 1270
rect 18151 1250 18197 1262
rect 18269 1262 18275 1270
rect 18309 1262 18315 1270
rect 18269 1250 18315 1262
rect 18387 1262 18393 1270
rect 18427 1262 18433 1270
rect 18387 1250 18433 1262
rect 18505 1262 18511 1270
rect 18545 1262 18551 1270
rect 18505 1250 18551 1262
rect 18623 1262 18629 1270
rect 18663 1262 18669 1270
rect 18623 1250 18669 1262
rect 18741 1262 18747 1270
rect 18781 1262 18787 1270
rect 18741 1250 18787 1262
rect 18859 1262 18865 1270
rect 18899 1262 18905 1270
rect 18859 1250 18905 1262
rect 18977 1262 18983 1270
rect 19017 1262 19023 1270
rect 18977 1250 19023 1262
rect 19095 1262 19101 1270
rect 19135 1262 19141 1270
rect 19095 1250 19141 1262
rect 19213 1262 19219 1270
rect 19253 1262 19259 1270
rect 19213 1250 19259 1262
rect 19331 1262 19337 1270
rect 19371 1262 19377 1270
rect 19331 1250 19377 1262
rect 19449 1262 19455 1270
rect 19489 1262 19495 1270
rect 19449 1250 19495 1262
rect 19567 1262 19573 1270
rect 19607 1262 19613 1270
rect 19567 1250 19613 1262
rect 4804 1178 4850 1190
rect 4804 1170 4810 1178
rect 4844 1170 4850 1178
rect 4922 1178 4968 1190
rect 4922 1170 4928 1178
rect 4962 1170 4968 1178
rect 5040 1178 5086 1190
rect 5040 1170 5046 1178
rect 5080 1170 5086 1178
rect 5158 1178 5204 1190
rect 5158 1170 5164 1178
rect 5198 1170 5204 1178
rect 5276 1178 5322 1190
rect 5276 1170 5282 1178
rect 5316 1170 5322 1178
rect 5394 1178 5440 1190
rect 5394 1170 5400 1178
rect 5434 1170 5440 1178
rect 5512 1178 5558 1190
rect 5512 1170 5518 1178
rect 5552 1170 5558 1178
rect 5630 1178 5676 1190
rect 5630 1170 5636 1178
rect 5670 1170 5676 1178
rect 5748 1178 5794 1190
rect 5748 1170 5754 1178
rect 5788 1170 5794 1178
rect 5866 1178 5912 1190
rect 5866 1170 5872 1178
rect 5906 1170 5912 1178
rect 5984 1178 6030 1190
rect 5984 1170 5990 1178
rect 6024 1170 6030 1178
rect 6102 1178 6148 1190
rect 6102 1170 6108 1178
rect 6142 1170 6148 1178
rect 6220 1178 6266 1190
rect 6220 1170 6226 1178
rect 6260 1170 6266 1178
rect 6338 1178 6384 1190
rect 6338 1170 6344 1178
rect 6378 1170 6384 1178
rect 6456 1178 6502 1190
rect 6456 1170 6462 1178
rect 6496 1170 6502 1178
rect 6574 1178 6620 1190
rect 6574 1170 6580 1178
rect 6614 1170 6620 1178
rect 6692 1178 6738 1190
rect 6692 1170 6698 1178
rect 6732 1170 6738 1178
rect 6810 1178 6856 1190
rect 6810 1170 6816 1178
rect 6850 1170 6856 1178
rect 6928 1178 6974 1190
rect 6928 1170 6934 1178
rect 6968 1170 6974 1178
rect 7046 1178 7092 1190
rect 7046 1170 7052 1178
rect 7086 1170 7092 1178
rect 7164 1178 7210 1190
rect 7164 1170 7170 1178
rect 7204 1170 7210 1178
rect 7282 1178 7328 1190
rect 7282 1170 7288 1178
rect 7322 1170 7328 1178
rect 7400 1178 7446 1190
rect 7400 1170 7406 1178
rect 7440 1170 7446 1178
rect 7518 1178 7564 1190
rect 7518 1170 7524 1178
rect 7558 1170 7564 1178
rect 7636 1178 7682 1190
rect 7636 1170 7642 1178
rect 7676 1170 7682 1178
rect 7754 1178 7800 1190
rect 7754 1170 7760 1178
rect 7794 1170 7800 1178
rect 7872 1178 7918 1190
rect 7872 1170 7878 1178
rect 7912 1170 7918 1178
rect 7990 1178 8036 1190
rect 7990 1170 7996 1178
rect 8030 1170 8036 1178
rect 8108 1178 8154 1190
rect 8108 1170 8114 1178
rect 8148 1170 8154 1178
rect 8226 1178 8272 1190
rect 8226 1170 8232 1178
rect 8266 1170 8272 1178
rect 8344 1178 8390 1190
rect 8344 1170 8350 1178
rect 8384 1170 8390 1178
rect 8462 1178 8508 1190
rect 8462 1170 8468 1178
rect 8502 1170 8508 1178
rect 8580 1178 8626 1190
rect 8580 1170 8586 1178
rect 8620 1170 8626 1178
rect 8698 1178 8744 1190
rect 8698 1170 8704 1178
rect 8738 1170 8744 1178
rect 8816 1178 8862 1190
rect 8816 1170 8822 1178
rect 8856 1170 8862 1178
rect 8934 1178 8980 1190
rect 8934 1170 8940 1178
rect 8974 1170 8980 1178
rect 9052 1178 9098 1190
rect 9052 1170 9058 1178
rect 9092 1170 9098 1178
rect 9170 1178 9216 1190
rect 9170 1170 9176 1178
rect 9210 1170 9216 1178
rect 9288 1178 9334 1190
rect 9288 1170 9294 1178
rect 9328 1170 9334 1178
rect 9406 1178 9452 1190
rect 9406 1170 9412 1178
rect 9446 1170 9452 1178
rect 9524 1178 9570 1190
rect 9524 1170 9530 1178
rect 9564 1170 9570 1178
rect 9642 1178 9688 1190
rect 9642 1170 9648 1178
rect 9682 1170 9688 1178
rect 9760 1178 9806 1190
rect 9760 1170 9766 1178
rect 9800 1170 9806 1178
rect 9878 1178 9924 1190
rect 9878 1170 9884 1178
rect 9918 1170 9924 1178
rect 9996 1178 10042 1190
rect 9996 1170 10002 1178
rect 10036 1170 10042 1178
rect 10114 1178 10160 1190
rect 10114 1170 10120 1178
rect 10154 1170 10160 1178
rect 10232 1178 10278 1190
rect 10232 1170 10238 1178
rect 10272 1170 10278 1178
rect 10350 1178 10396 1190
rect 10350 1170 10356 1178
rect 10390 1170 10396 1178
rect 10468 1178 10514 1190
rect 10468 1170 10474 1178
rect 10508 1170 10514 1178
rect 10586 1178 10632 1190
rect 10586 1170 10592 1178
rect 10626 1170 10632 1178
rect 10704 1178 10750 1190
rect 10704 1170 10710 1178
rect 10744 1170 10750 1178
rect 4791 610 4801 1170
rect 4853 610 4863 1170
rect 4907 610 4917 1170
rect 4969 610 4979 1170
rect 5027 610 5037 1170
rect 5089 610 5099 1170
rect 5143 610 5153 1170
rect 5205 610 5215 1170
rect 5263 610 5273 1170
rect 5325 610 5335 1170
rect 5379 610 5389 1170
rect 5441 610 5451 1170
rect 5499 610 5509 1170
rect 5561 610 5571 1170
rect 5615 610 5625 1170
rect 5677 610 5687 1170
rect 5735 610 5745 1170
rect 5797 610 5807 1170
rect 5851 610 5861 1170
rect 5913 610 5923 1170
rect 5971 610 5981 1170
rect 6033 610 6043 1170
rect 6087 610 6097 1170
rect 6149 610 6159 1170
rect 6207 610 6217 1170
rect 6269 610 6279 1170
rect 6323 610 6333 1170
rect 6385 610 6395 1170
rect 6443 610 6453 1170
rect 6505 610 6515 1170
rect 6559 610 6569 1170
rect 6621 610 6631 1170
rect 6679 610 6689 1170
rect 6741 610 6751 1170
rect 6795 610 6805 1170
rect 6857 610 6867 1170
rect 6915 610 6925 1170
rect 6977 610 6987 1170
rect 7031 610 7041 1170
rect 7093 610 7103 1170
rect 7151 610 7161 1170
rect 7213 610 7223 1170
rect 7267 610 7277 1170
rect 7329 610 7339 1170
rect 7387 610 7397 1170
rect 7449 610 7459 1170
rect 7503 610 7513 1170
rect 7565 610 7575 1170
rect 7623 610 7633 1170
rect 7685 610 7695 1170
rect 7739 610 7749 1170
rect 7801 610 7811 1170
rect 7859 610 7869 1170
rect 7921 610 7931 1170
rect 7975 610 7985 1170
rect 8037 610 8047 1170
rect 8095 610 8105 1170
rect 8157 610 8167 1170
rect 8211 610 8221 1170
rect 8273 610 8283 1170
rect 8331 610 8341 1170
rect 8393 610 8403 1170
rect 8447 610 8457 1170
rect 8509 610 8519 1170
rect 8567 610 8577 1170
rect 8629 610 8639 1170
rect 8683 610 8693 1170
rect 8745 610 8755 1170
rect 8803 610 8813 1170
rect 8865 610 8875 1170
rect 8919 610 8929 1170
rect 8981 610 8991 1170
rect 9039 610 9049 1170
rect 9101 610 9111 1170
rect 9155 610 9165 1170
rect 9217 610 9227 1170
rect 9275 610 9285 1170
rect 9337 610 9347 1170
rect 9391 610 9401 1170
rect 9453 610 9463 1170
rect 9511 610 9521 1170
rect 9573 610 9583 1170
rect 9627 610 9637 1170
rect 9689 610 9699 1170
rect 9747 610 9757 1170
rect 9809 610 9819 1170
rect 9863 610 9873 1170
rect 9925 610 9935 1170
rect 9983 610 9993 1170
rect 10045 610 10055 1170
rect 10099 610 10109 1170
rect 10161 610 10171 1170
rect 10219 610 10229 1170
rect 10281 610 10291 1170
rect 10335 610 10345 1170
rect 10397 610 10407 1170
rect 10455 610 10465 1170
rect 10517 610 10527 1170
rect 10571 610 10581 1170
rect 10633 610 10643 1170
rect 10691 610 10701 1170
rect 10753 610 10763 1170
rect 15619 1163 16452 1247
rect 19743 1247 19782 1281
rect 19816 1247 19854 1281
rect 19888 1247 19926 1281
rect 19960 1247 19998 1281
rect 20032 1247 20070 1281
rect 20104 1247 20142 1281
rect 20176 1247 20214 1281
rect 20248 1247 20286 1281
rect 20320 1247 20358 1281
rect 20392 1247 20430 1281
rect 20464 1247 20502 1281
rect 20536 1247 20575 1281
rect 20727 1270 20737 1830
rect 20789 1270 20799 1830
rect 20845 1270 20855 1830
rect 20907 1270 20917 1830
rect 20963 1270 20973 1830
rect 21025 1270 21035 1830
rect 21081 1270 21091 1830
rect 21143 1270 21153 1830
rect 21199 1270 21209 1830
rect 21261 1270 21271 1830
rect 21317 1270 21327 1830
rect 21379 1270 21389 1830
rect 21435 1270 21445 1830
rect 21497 1270 21507 1830
rect 21553 1270 21563 1830
rect 21615 1270 21625 1830
rect 21671 1270 21681 1830
rect 21733 1270 21743 1830
rect 21789 1270 21799 1830
rect 21851 1270 21861 1830
rect 21907 1270 21917 1830
rect 21969 1270 21979 1830
rect 22025 1270 22035 1830
rect 22087 1270 22097 1830
rect 22143 1270 22153 1830
rect 22205 1270 22215 1830
rect 22261 1270 22271 1830
rect 22323 1270 22333 1830
rect 22379 1270 22389 1830
rect 22441 1270 22451 1830
rect 22497 1270 22507 1830
rect 22559 1270 22569 1830
rect 22615 1270 22625 1830
rect 22677 1270 22687 1830
rect 22733 1270 22743 1830
rect 22795 1270 22805 1830
rect 22851 1270 22861 1830
rect 22913 1270 22923 1830
rect 22969 1270 22979 1830
rect 23031 1270 23041 1830
rect 23087 1270 23097 1830
rect 23149 1270 23159 1830
rect 23205 1270 23215 1830
rect 23267 1270 23277 1830
rect 23323 1270 23333 1830
rect 23385 1270 23395 1830
rect 23441 1270 23451 1830
rect 23503 1270 23513 1830
rect 23559 1270 23569 1830
rect 23621 1270 23631 1830
rect 23677 1270 23687 1830
rect 23739 1270 23749 1830
rect 23867 1801 23895 1853
rect 23947 1801 23975 1853
rect 24027 1839 24049 1853
rect 24107 1839 24121 1853
rect 24187 1839 24193 1853
rect 24371 1839 24375 1853
rect 24443 1839 24455 1853
rect 24515 1839 24535 1853
rect 24027 1801 24055 1839
rect 24107 1801 24135 1839
rect 24187 1801 24215 1839
rect 24267 1801 24295 1839
rect 24347 1801 24375 1839
rect 24427 1801 24455 1839
rect 24507 1801 24535 1839
rect 24587 1801 24615 1853
rect 24667 1801 24695 1853
rect 24747 1801 24775 1853
rect 24827 1801 24855 1853
rect 24907 1801 24935 1853
rect 24987 1801 25015 1853
rect 25067 1801 25081 1853
rect 23867 1799 25081 1801
rect 23867 1773 23905 1799
rect 23939 1773 23977 1799
rect 24011 1773 24049 1799
rect 24083 1773 24121 1799
rect 24155 1773 24193 1799
rect 24227 1773 24265 1799
rect 24299 1773 24337 1799
rect 24371 1773 24409 1799
rect 24443 1773 24481 1799
rect 24515 1773 24553 1799
rect 24587 1773 24625 1799
rect 24659 1773 25081 1799
rect 23867 1721 23895 1773
rect 23947 1721 23975 1773
rect 24027 1765 24049 1773
rect 24107 1765 24121 1773
rect 24187 1765 24193 1773
rect 24371 1765 24375 1773
rect 24443 1765 24455 1773
rect 24515 1765 24535 1773
rect 24027 1725 24055 1765
rect 24107 1725 24135 1765
rect 24187 1725 24215 1765
rect 24267 1725 24295 1765
rect 24347 1725 24375 1765
rect 24427 1725 24455 1765
rect 24507 1725 24535 1765
rect 24027 1721 24049 1725
rect 24107 1721 24121 1725
rect 24187 1721 24193 1725
rect 24371 1721 24375 1725
rect 24443 1721 24455 1725
rect 24515 1721 24535 1725
rect 24587 1721 24615 1773
rect 24667 1721 24695 1773
rect 24747 1721 24775 1773
rect 24827 1721 24855 1773
rect 24907 1721 24935 1773
rect 24987 1721 25015 1773
rect 25067 1721 25081 1773
rect 23867 1693 23905 1721
rect 23939 1693 23977 1721
rect 24011 1693 24049 1721
rect 24083 1693 24121 1721
rect 24155 1693 24193 1721
rect 24227 1693 24265 1721
rect 24299 1693 24337 1721
rect 24371 1693 24409 1721
rect 24443 1693 24481 1721
rect 24515 1693 24553 1721
rect 24587 1693 24625 1721
rect 24659 1693 25081 1721
rect 23867 1641 23895 1693
rect 23947 1641 23975 1693
rect 24027 1691 24049 1693
rect 24107 1691 24121 1693
rect 24187 1691 24193 1693
rect 24371 1691 24375 1693
rect 24443 1691 24455 1693
rect 24515 1691 24535 1693
rect 24027 1651 24055 1691
rect 24107 1651 24135 1691
rect 24187 1651 24215 1691
rect 24267 1651 24295 1691
rect 24347 1651 24375 1691
rect 24427 1651 24455 1691
rect 24507 1651 24535 1691
rect 24027 1641 24049 1651
rect 24107 1641 24121 1651
rect 24187 1641 24193 1651
rect 24371 1641 24375 1651
rect 24443 1641 24455 1651
rect 24515 1641 24535 1651
rect 24587 1641 24615 1693
rect 24667 1641 24695 1693
rect 24747 1641 24775 1693
rect 24827 1641 24855 1693
rect 24907 1641 24935 1693
rect 24987 1641 25015 1693
rect 25067 1641 25081 1693
rect 23867 1617 23905 1641
rect 23939 1617 23977 1641
rect 24011 1617 24049 1641
rect 24083 1617 24121 1641
rect 24155 1617 24193 1641
rect 24227 1617 24265 1641
rect 24299 1617 24337 1641
rect 24371 1617 24409 1641
rect 24443 1617 24481 1641
rect 24515 1617 24553 1641
rect 24587 1617 24625 1641
rect 24659 1617 25081 1641
rect 23867 1613 25081 1617
rect 23867 1561 23895 1613
rect 23947 1561 23975 1613
rect 24027 1577 24055 1613
rect 24107 1577 24135 1613
rect 24187 1577 24215 1613
rect 24267 1577 24295 1613
rect 24347 1577 24375 1613
rect 24427 1577 24455 1613
rect 24507 1577 24535 1613
rect 24027 1561 24049 1577
rect 24107 1561 24121 1577
rect 24187 1561 24193 1577
rect 24371 1561 24375 1577
rect 24443 1561 24455 1577
rect 24515 1561 24535 1577
rect 24587 1561 24615 1613
rect 24667 1561 24695 1613
rect 24747 1561 24775 1613
rect 24827 1561 24855 1613
rect 24907 1561 24935 1613
rect 24987 1561 25015 1613
rect 25067 1561 25081 1613
rect 23867 1543 23905 1561
rect 23939 1543 23977 1561
rect 24011 1543 24049 1561
rect 24083 1543 24121 1561
rect 24155 1543 24193 1561
rect 24227 1543 24265 1561
rect 24299 1543 24337 1561
rect 24371 1543 24409 1561
rect 24443 1543 24481 1561
rect 24515 1543 24553 1561
rect 24587 1543 24625 1561
rect 24659 1543 25081 1561
rect 23867 1533 25081 1543
rect 23867 1481 23895 1533
rect 23947 1481 23975 1533
rect 24027 1503 24055 1533
rect 24107 1503 24135 1533
rect 24187 1503 24215 1533
rect 24267 1503 24295 1533
rect 24347 1503 24375 1533
rect 24427 1503 24455 1533
rect 24507 1503 24535 1533
rect 24027 1481 24049 1503
rect 24107 1481 24121 1503
rect 24187 1481 24193 1503
rect 24371 1481 24375 1503
rect 24443 1481 24455 1503
rect 24515 1481 24535 1503
rect 24587 1481 24615 1533
rect 24667 1481 24695 1533
rect 24747 1481 24775 1533
rect 24827 1481 24855 1533
rect 24907 1481 24935 1533
rect 24987 1481 25015 1533
rect 25067 1481 25081 1533
rect 23867 1469 23905 1481
rect 23939 1469 23977 1481
rect 24011 1469 24049 1481
rect 24083 1469 24121 1481
rect 24155 1469 24193 1481
rect 24227 1469 24265 1481
rect 24299 1469 24337 1481
rect 24371 1469 24409 1481
rect 24443 1469 24481 1481
rect 24515 1469 24553 1481
rect 24587 1469 24625 1481
rect 24659 1469 25081 1481
rect 23867 1453 25081 1469
rect 23867 1401 23895 1453
rect 23947 1401 23975 1453
rect 24027 1429 24055 1453
rect 24107 1429 24135 1453
rect 24187 1429 24215 1453
rect 24267 1429 24295 1453
rect 24347 1429 24375 1453
rect 24427 1429 24455 1453
rect 24507 1429 24535 1453
rect 24027 1401 24049 1429
rect 24107 1401 24121 1429
rect 24187 1401 24193 1429
rect 24371 1401 24375 1429
rect 24443 1401 24455 1429
rect 24515 1401 24535 1429
rect 24587 1401 24615 1453
rect 24667 1401 24695 1453
rect 24747 1401 24775 1453
rect 24827 1401 24855 1453
rect 24907 1401 24935 1453
rect 24987 1401 25015 1453
rect 25067 1401 25081 1453
rect 23867 1395 23905 1401
rect 23939 1395 23977 1401
rect 24011 1395 24049 1401
rect 24083 1395 24121 1401
rect 24155 1395 24193 1401
rect 24227 1395 24265 1401
rect 24299 1395 24337 1401
rect 24371 1395 24409 1401
rect 24443 1395 24481 1401
rect 24515 1395 24553 1401
rect 24587 1395 24625 1401
rect 24659 1395 25081 1401
rect 23867 1373 25081 1395
rect 23867 1321 23895 1373
rect 23947 1321 23975 1373
rect 24027 1355 24055 1373
rect 24107 1355 24135 1373
rect 24187 1355 24215 1373
rect 24267 1355 24295 1373
rect 24347 1355 24375 1373
rect 24427 1355 24455 1373
rect 24507 1355 24535 1373
rect 24027 1321 24049 1355
rect 24107 1321 24121 1355
rect 24187 1321 24193 1355
rect 24371 1321 24375 1355
rect 24443 1321 24455 1355
rect 24515 1321 24535 1355
rect 24587 1321 24615 1373
rect 24667 1321 24695 1373
rect 24747 1321 24775 1373
rect 24827 1321 24855 1373
rect 24907 1321 24935 1373
rect 24987 1321 25015 1373
rect 25067 1321 25081 1373
rect 23867 1293 25081 1321
rect 20740 1262 20746 1270
rect 20780 1262 20786 1270
rect 20740 1250 20786 1262
rect 20858 1262 20864 1270
rect 20898 1262 20904 1270
rect 20858 1250 20904 1262
rect 20976 1262 20982 1270
rect 21016 1262 21022 1270
rect 20976 1250 21022 1262
rect 21094 1262 21100 1270
rect 21134 1262 21140 1270
rect 21094 1250 21140 1262
rect 21212 1262 21218 1270
rect 21252 1262 21258 1270
rect 21212 1250 21258 1262
rect 21330 1262 21336 1270
rect 21370 1262 21376 1270
rect 21330 1250 21376 1262
rect 21448 1262 21454 1270
rect 21488 1262 21494 1270
rect 21448 1250 21494 1262
rect 21566 1262 21572 1270
rect 21606 1262 21612 1270
rect 21566 1250 21612 1262
rect 21684 1262 21690 1270
rect 21724 1262 21730 1270
rect 21684 1250 21730 1262
rect 21802 1262 21808 1270
rect 21842 1262 21848 1270
rect 21802 1250 21848 1262
rect 21920 1262 21926 1270
rect 21960 1262 21966 1270
rect 21920 1250 21966 1262
rect 22038 1262 22044 1270
rect 22078 1262 22084 1270
rect 22038 1250 22084 1262
rect 22156 1262 22162 1270
rect 22196 1262 22202 1270
rect 22156 1250 22202 1262
rect 22274 1262 22280 1270
rect 22314 1262 22320 1270
rect 22274 1250 22320 1262
rect 22392 1262 22398 1270
rect 22432 1262 22438 1270
rect 22392 1250 22438 1262
rect 22510 1262 22516 1270
rect 22550 1262 22556 1270
rect 22510 1250 22556 1262
rect 22628 1262 22634 1270
rect 22668 1262 22674 1270
rect 22628 1250 22674 1262
rect 22746 1262 22752 1270
rect 22786 1262 22792 1270
rect 22746 1250 22792 1262
rect 22864 1262 22870 1270
rect 22904 1262 22910 1270
rect 22864 1250 22910 1262
rect 22982 1262 22988 1270
rect 23022 1262 23028 1270
rect 22982 1250 23028 1262
rect 23100 1262 23106 1270
rect 23140 1262 23146 1270
rect 23100 1250 23146 1262
rect 23218 1262 23224 1270
rect 23258 1262 23264 1270
rect 23218 1250 23264 1262
rect 23336 1262 23342 1270
rect 23376 1262 23382 1270
rect 23336 1250 23382 1262
rect 23454 1262 23460 1270
rect 23494 1262 23500 1270
rect 23454 1250 23500 1262
rect 23572 1262 23578 1270
rect 23612 1262 23618 1270
rect 23572 1250 23618 1262
rect 23690 1262 23696 1270
rect 23730 1262 23736 1270
rect 23690 1250 23736 1262
rect 19743 1163 20575 1247
rect 23867 1241 23895 1293
rect 23947 1241 23975 1293
rect 24027 1281 24055 1293
rect 24107 1281 24135 1293
rect 24187 1281 24215 1293
rect 24267 1281 24295 1293
rect 24347 1281 24375 1293
rect 24427 1281 24455 1293
rect 24507 1281 24535 1293
rect 24027 1247 24049 1281
rect 24107 1247 24121 1281
rect 24187 1247 24193 1281
rect 24371 1247 24375 1281
rect 24443 1247 24455 1281
rect 24515 1247 24535 1281
rect 24027 1241 24055 1247
rect 24107 1241 24135 1247
rect 24187 1241 24215 1247
rect 24267 1241 24295 1247
rect 24347 1241 24375 1247
rect 24427 1241 24455 1247
rect 24507 1241 24535 1247
rect 24587 1241 24615 1293
rect 24667 1241 24695 1293
rect 24747 1241 24775 1293
rect 24827 1241 24855 1293
rect 24907 1241 24935 1293
rect 24987 1241 25015 1293
rect 25067 1241 25081 1293
rect 23867 1227 25081 1241
rect 23903 1163 25079 1227
rect 12471 1149 25079 1163
rect 12471 1101 12485 1149
rect 12471 1067 12479 1101
rect 12537 1097 12565 1149
rect 12617 1097 12645 1149
rect 12697 1097 12725 1149
rect 12777 1097 12805 1149
rect 12857 1097 12885 1149
rect 12937 1097 12965 1149
rect 13017 1097 13045 1149
rect 13097 1097 13125 1149
rect 13177 1097 13205 1149
rect 13257 1097 13285 1149
rect 13337 1097 13365 1149
rect 13417 1097 13445 1149
rect 13497 1097 13525 1149
rect 13577 1097 13605 1149
rect 13657 1097 13685 1149
rect 13737 1097 13765 1149
rect 13817 1097 13845 1149
rect 13897 1097 13925 1149
rect 13977 1097 14005 1149
rect 14057 1097 14085 1149
rect 14137 1097 14165 1149
rect 14217 1097 14245 1149
rect 14297 1097 14325 1149
rect 14377 1097 14405 1149
rect 14457 1097 14485 1149
rect 14537 1097 14565 1149
rect 14617 1097 14645 1149
rect 14697 1097 14725 1149
rect 14777 1097 14805 1149
rect 14857 1097 14885 1149
rect 14937 1097 14965 1149
rect 15017 1097 15045 1149
rect 15097 1097 15125 1149
rect 15177 1097 15205 1149
rect 15257 1097 15285 1149
rect 15337 1097 15365 1149
rect 15417 1097 15445 1149
rect 15497 1097 15525 1149
rect 15577 1097 15605 1149
rect 15657 1097 15685 1149
rect 15737 1097 15765 1149
rect 15817 1097 15845 1149
rect 15897 1097 15925 1149
rect 15977 1097 16005 1149
rect 16057 1097 16085 1149
rect 16137 1097 16165 1149
rect 16217 1097 16245 1149
rect 16297 1097 16325 1149
rect 16377 1097 16405 1149
rect 16457 1097 16485 1149
rect 16537 1097 16565 1149
rect 16617 1097 16645 1149
rect 16697 1097 16725 1149
rect 16777 1097 16805 1149
rect 16857 1097 16885 1149
rect 16937 1097 16965 1149
rect 17017 1097 17045 1149
rect 17097 1097 17125 1149
rect 17177 1097 17205 1149
rect 17257 1097 17285 1149
rect 17337 1097 17365 1149
rect 17417 1097 17445 1149
rect 17497 1097 17525 1149
rect 17577 1097 17605 1149
rect 17657 1097 17685 1149
rect 17737 1097 17765 1149
rect 17817 1097 17845 1149
rect 17897 1097 17925 1149
rect 17977 1097 18005 1149
rect 18057 1097 18085 1149
rect 18137 1097 18165 1149
rect 18217 1097 18245 1149
rect 18297 1097 18325 1149
rect 18377 1097 18405 1149
rect 18457 1097 18485 1149
rect 18537 1097 18565 1149
rect 18617 1097 18645 1149
rect 18697 1097 18725 1149
rect 18777 1097 18805 1149
rect 18857 1097 18885 1149
rect 18937 1097 18965 1149
rect 19017 1097 19045 1149
rect 19097 1097 19125 1149
rect 19177 1097 19205 1149
rect 19257 1097 19285 1149
rect 19337 1097 19365 1149
rect 19417 1097 19445 1149
rect 19497 1097 19525 1149
rect 19577 1097 19605 1149
rect 19657 1097 19685 1149
rect 19737 1097 19765 1149
rect 19817 1097 19845 1149
rect 19897 1097 19925 1149
rect 19977 1097 20005 1149
rect 20057 1097 20085 1149
rect 20137 1097 20165 1149
rect 20217 1097 20245 1149
rect 20297 1097 20325 1149
rect 20377 1097 20405 1149
rect 20457 1097 20485 1149
rect 20537 1097 20565 1149
rect 20617 1097 20645 1149
rect 20697 1097 20725 1149
rect 20777 1097 20805 1149
rect 20857 1097 20885 1149
rect 20937 1097 20965 1149
rect 21017 1097 21045 1149
rect 21097 1097 21125 1149
rect 21177 1097 21205 1149
rect 21257 1097 21285 1149
rect 21337 1097 21365 1149
rect 21417 1097 21445 1149
rect 21497 1097 21525 1149
rect 21577 1097 21605 1149
rect 21657 1097 21685 1149
rect 21737 1097 21765 1149
rect 21817 1097 21845 1149
rect 21897 1097 21925 1149
rect 21977 1097 22005 1149
rect 22057 1097 22085 1149
rect 22137 1097 22165 1149
rect 22217 1097 22245 1149
rect 22297 1097 22325 1149
rect 22377 1097 22405 1149
rect 22457 1097 22485 1149
rect 22537 1097 22565 1149
rect 22617 1097 22645 1149
rect 22697 1097 22725 1149
rect 22777 1097 22805 1149
rect 22857 1097 22885 1149
rect 22937 1097 22965 1149
rect 23017 1097 23045 1149
rect 23097 1097 23125 1149
rect 23177 1097 23205 1149
rect 23257 1097 23285 1149
rect 23337 1097 23365 1149
rect 23417 1097 23445 1149
rect 23497 1097 23525 1149
rect 23577 1097 23605 1149
rect 23657 1097 23685 1149
rect 23737 1097 23765 1149
rect 23817 1097 23845 1149
rect 23897 1097 23925 1149
rect 23977 1097 24005 1149
rect 24057 1097 24085 1149
rect 24137 1097 24165 1149
rect 24217 1097 24245 1149
rect 24297 1097 24325 1149
rect 24377 1097 24405 1149
rect 24457 1097 25079 1149
rect 12513 1069 25079 1097
rect 12471 1017 12485 1067
rect 12537 1017 12565 1069
rect 12617 1017 12645 1069
rect 12697 1017 12725 1069
rect 12777 1017 12805 1069
rect 12857 1017 12885 1069
rect 12937 1017 12965 1069
rect 13017 1017 13045 1069
rect 13097 1017 13125 1069
rect 13177 1017 13205 1069
rect 13257 1017 13285 1069
rect 13337 1017 13365 1069
rect 13417 1017 13445 1069
rect 13497 1017 13525 1069
rect 13577 1017 13605 1069
rect 13657 1017 13685 1069
rect 13737 1017 13765 1069
rect 13817 1017 13845 1069
rect 13897 1017 13925 1069
rect 13977 1017 14005 1069
rect 14057 1017 14085 1069
rect 14137 1017 14165 1069
rect 14217 1017 14245 1069
rect 14297 1017 14325 1069
rect 14377 1017 14405 1069
rect 14457 1017 14485 1069
rect 14537 1017 14565 1069
rect 14617 1017 14645 1069
rect 14697 1017 14725 1069
rect 14777 1017 14805 1069
rect 14857 1017 14885 1069
rect 14937 1017 14965 1069
rect 15017 1017 15045 1069
rect 15097 1017 15125 1069
rect 15177 1017 15205 1069
rect 15257 1017 15285 1069
rect 15337 1017 15365 1069
rect 15417 1017 15445 1069
rect 15497 1017 15525 1069
rect 15577 1017 15605 1069
rect 15657 1017 15685 1069
rect 15737 1017 15765 1069
rect 15817 1017 15845 1069
rect 15897 1017 15925 1069
rect 15977 1017 16005 1069
rect 16057 1017 16085 1069
rect 16137 1017 16165 1069
rect 16217 1017 16245 1069
rect 16297 1017 16325 1069
rect 16377 1017 16405 1069
rect 16457 1017 16485 1069
rect 16537 1017 16565 1069
rect 16617 1017 16645 1069
rect 16697 1017 16725 1069
rect 16777 1017 16805 1069
rect 16857 1017 16885 1069
rect 16937 1017 16965 1069
rect 17017 1017 17045 1069
rect 17097 1017 17125 1069
rect 17177 1017 17205 1069
rect 17257 1017 17285 1069
rect 17337 1017 17365 1069
rect 17417 1017 17445 1069
rect 17497 1017 17525 1069
rect 17577 1017 17605 1069
rect 17657 1017 17685 1069
rect 17737 1017 17765 1069
rect 17817 1017 17845 1069
rect 17897 1017 17925 1069
rect 17977 1017 18005 1069
rect 18057 1017 18085 1069
rect 18137 1017 18165 1069
rect 18217 1017 18245 1069
rect 18297 1017 18325 1069
rect 18377 1017 18405 1069
rect 18457 1017 18485 1069
rect 18537 1017 18565 1069
rect 18617 1017 18645 1069
rect 18697 1017 18725 1069
rect 18777 1017 18805 1069
rect 18857 1017 18885 1069
rect 18937 1017 18965 1069
rect 19017 1017 19045 1069
rect 19097 1017 19125 1069
rect 19177 1017 19205 1069
rect 19257 1017 19285 1069
rect 19337 1017 19365 1069
rect 19417 1017 19445 1069
rect 19497 1017 19525 1069
rect 19577 1017 19605 1069
rect 19657 1017 19685 1069
rect 19737 1017 19765 1069
rect 19817 1017 19845 1069
rect 19897 1017 19925 1069
rect 19977 1017 20005 1069
rect 20057 1017 20085 1069
rect 20137 1017 20165 1069
rect 20217 1017 20245 1069
rect 20297 1017 20325 1069
rect 20377 1017 20405 1069
rect 20457 1017 20485 1069
rect 20537 1017 20565 1069
rect 20617 1017 20645 1069
rect 20697 1017 20725 1069
rect 20777 1017 20805 1069
rect 20857 1017 20885 1069
rect 20937 1017 20965 1069
rect 21017 1017 21045 1069
rect 21097 1017 21125 1069
rect 21177 1017 21205 1069
rect 21257 1017 21285 1069
rect 21337 1017 21365 1069
rect 21417 1017 21445 1069
rect 21497 1017 21525 1069
rect 21577 1017 21605 1069
rect 21657 1017 21685 1069
rect 21737 1017 21765 1069
rect 21817 1017 21845 1069
rect 21897 1017 21925 1069
rect 21977 1017 22005 1069
rect 22057 1017 22085 1069
rect 22137 1017 22165 1069
rect 22217 1017 22245 1069
rect 22297 1017 22325 1069
rect 22377 1017 22405 1069
rect 22457 1017 22485 1069
rect 22537 1017 22565 1069
rect 22617 1017 22645 1069
rect 22697 1017 22725 1069
rect 22777 1017 22805 1069
rect 22857 1017 22885 1069
rect 22937 1017 22965 1069
rect 23017 1017 23045 1069
rect 23097 1017 23125 1069
rect 23177 1017 23205 1069
rect 23257 1017 23285 1069
rect 23337 1017 23365 1069
rect 23417 1017 23445 1069
rect 23497 1017 23525 1069
rect 23577 1017 23605 1069
rect 23657 1017 23685 1069
rect 23737 1017 23765 1069
rect 23817 1017 23845 1069
rect 23897 1017 23925 1069
rect 23977 1017 24005 1069
rect 24057 1017 24085 1069
rect 24137 1017 24165 1069
rect 24217 1017 24245 1069
rect 24297 1017 24325 1069
rect 24377 1017 24405 1069
rect 24457 1017 25079 1069
rect 12471 1004 25079 1017
rect 12471 1003 24471 1004
rect 4804 602 4810 610
rect 4844 602 4850 610
rect 4804 590 4850 602
rect 4922 602 4928 610
rect 4962 602 4968 610
rect 4922 590 4968 602
rect 5040 602 5046 610
rect 5080 602 5086 610
rect 5040 590 5086 602
rect 5158 602 5164 610
rect 5198 602 5204 610
rect 5158 590 5204 602
rect 5276 602 5282 610
rect 5316 602 5322 610
rect 5276 590 5322 602
rect 5394 602 5400 610
rect 5434 602 5440 610
rect 5394 590 5440 602
rect 5512 602 5518 610
rect 5552 602 5558 610
rect 5512 590 5558 602
rect 5630 602 5636 610
rect 5670 602 5676 610
rect 5630 590 5676 602
rect 5748 602 5754 610
rect 5788 602 5794 610
rect 5748 590 5794 602
rect 5866 602 5872 610
rect 5906 602 5912 610
rect 5866 590 5912 602
rect 5984 602 5990 610
rect 6024 602 6030 610
rect 5984 590 6030 602
rect 6102 602 6108 610
rect 6142 602 6148 610
rect 6102 590 6148 602
rect 6220 602 6226 610
rect 6260 602 6266 610
rect 6220 590 6266 602
rect 6338 602 6344 610
rect 6378 602 6384 610
rect 6338 590 6384 602
rect 6456 602 6462 610
rect 6496 602 6502 610
rect 6456 590 6502 602
rect 6574 602 6580 610
rect 6614 602 6620 610
rect 6574 590 6620 602
rect 6692 602 6698 610
rect 6732 602 6738 610
rect 6692 590 6738 602
rect 6810 602 6816 610
rect 6850 602 6856 610
rect 6810 590 6856 602
rect 6928 602 6934 610
rect 6968 602 6974 610
rect 6928 590 6974 602
rect 7046 602 7052 610
rect 7086 602 7092 610
rect 7046 590 7092 602
rect 7164 602 7170 610
rect 7204 602 7210 610
rect 7164 590 7210 602
rect 7282 602 7288 610
rect 7322 602 7328 610
rect 7282 590 7328 602
rect 7400 602 7406 610
rect 7440 602 7446 610
rect 7400 590 7446 602
rect 7518 602 7524 610
rect 7558 602 7564 610
rect 7518 590 7564 602
rect 7636 602 7642 610
rect 7676 602 7682 610
rect 7636 590 7682 602
rect 7754 602 7760 610
rect 7794 602 7800 610
rect 7754 590 7800 602
rect 7872 602 7878 610
rect 7912 602 7918 610
rect 7872 590 7918 602
rect 7990 602 7996 610
rect 8030 602 8036 610
rect 7990 590 8036 602
rect 8108 602 8114 610
rect 8148 602 8154 610
rect 8108 590 8154 602
rect 8226 602 8232 610
rect 8266 602 8272 610
rect 8226 590 8272 602
rect 8344 602 8350 610
rect 8384 602 8390 610
rect 8344 590 8390 602
rect 8462 602 8468 610
rect 8502 602 8508 610
rect 8462 590 8508 602
rect 8580 602 8586 610
rect 8620 602 8626 610
rect 8580 590 8626 602
rect 8698 602 8704 610
rect 8738 602 8744 610
rect 8698 590 8744 602
rect 8816 602 8822 610
rect 8856 602 8862 610
rect 8816 590 8862 602
rect 8934 602 8940 610
rect 8974 602 8980 610
rect 8934 590 8980 602
rect 9052 602 9058 610
rect 9092 602 9098 610
rect 9052 590 9098 602
rect 9170 602 9176 610
rect 9210 602 9216 610
rect 9170 590 9216 602
rect 9288 602 9294 610
rect 9328 602 9334 610
rect 9288 590 9334 602
rect 9406 602 9412 610
rect 9446 602 9452 610
rect 9406 590 9452 602
rect 9524 602 9530 610
rect 9564 602 9570 610
rect 9524 590 9570 602
rect 9642 602 9648 610
rect 9682 602 9688 610
rect 9642 590 9688 602
rect 9760 602 9766 610
rect 9800 602 9806 610
rect 9760 590 9806 602
rect 9878 602 9884 610
rect 9918 602 9924 610
rect 9878 590 9924 602
rect 9996 602 10002 610
rect 10036 602 10042 610
rect 9996 590 10042 602
rect 10114 602 10120 610
rect 10154 602 10160 610
rect 10114 590 10160 602
rect 10232 602 10238 610
rect 10272 602 10278 610
rect 10232 590 10278 602
rect 10350 602 10356 610
rect 10390 602 10396 610
rect 10350 590 10396 602
rect 10468 602 10474 610
rect 10508 602 10514 610
rect 10468 590 10514 602
rect 10586 602 10592 610
rect 10626 602 10632 610
rect 10586 590 10632 602
rect 10704 602 10710 610
rect 10744 602 10750 610
rect 10704 590 10750 602
rect 4847 395 4857 549
rect 4915 395 4925 549
rect 4965 395 4975 549
rect 5033 395 5043 549
rect 5083 395 5093 549
rect 5151 395 5161 549
rect 5201 395 5211 549
rect 5269 395 5279 549
rect 5319 395 5329 549
rect 5387 395 5397 549
rect 5437 395 5447 549
rect 5505 395 5515 549
rect 5555 395 5565 549
rect 5623 395 5633 549
rect 5673 395 5683 549
rect 5741 395 5751 549
rect 5791 395 5801 549
rect 5859 395 5869 549
rect 5909 395 5919 549
rect 5977 395 5987 549
rect 6027 395 6037 549
rect 6095 395 6105 549
rect 6145 395 6155 549
rect 6213 395 6223 549
rect 6263 395 6273 549
rect 6331 395 6341 549
rect 6381 395 6391 549
rect 6449 395 6459 549
rect 6499 395 6509 549
rect 6567 395 6577 549
rect 6617 395 6627 549
rect 6685 395 6695 549
rect 6735 395 6745 549
rect 6803 395 6813 549
rect 6853 395 6863 549
rect 6921 395 6931 549
rect 6971 395 6981 549
rect 7039 395 7049 549
rect 7089 395 7099 549
rect 7157 395 7167 549
rect 7207 395 7217 549
rect 7275 395 7285 549
rect 7325 395 7335 549
rect 7393 395 7403 549
rect 7443 395 7453 549
rect 7511 395 7521 549
rect 7561 395 7571 549
rect 7629 395 7639 549
rect 7679 395 7689 549
rect 7747 395 7757 549
rect 7797 395 7807 549
rect 7865 395 7875 549
rect 7915 395 7925 549
rect 7983 395 7993 549
rect 8033 395 8043 549
rect 8101 395 8111 549
rect 8151 395 8161 549
rect 8219 395 8229 549
rect 8269 395 8279 549
rect 8337 395 8347 549
rect 8387 395 8397 549
rect 8455 395 8465 549
rect 8505 395 8515 549
rect 8573 395 8583 549
rect 8623 395 8633 549
rect 8691 395 8701 549
rect 8741 395 8751 549
rect 8809 395 8819 549
rect 8859 395 8869 549
rect 8927 395 8937 549
rect 8977 395 8987 549
rect 9045 395 9055 549
rect 9095 395 9105 549
rect 9163 395 9173 549
rect 9213 395 9223 549
rect 9281 395 9291 549
rect 9331 395 9341 549
rect 9399 395 9409 549
rect 9449 395 9459 549
rect 9517 395 9527 549
rect 9567 395 9577 549
rect 9635 395 9645 549
rect 9685 395 9695 549
rect 9753 395 9763 549
rect 9803 395 9813 549
rect 9871 395 9881 549
rect 9921 395 9931 549
rect 9989 395 9999 549
rect 10039 395 10049 549
rect 10107 395 10117 549
rect 10157 395 10167 549
rect 10225 395 10235 549
rect 10275 395 10285 549
rect 10343 395 10353 549
rect 10393 395 10403 549
rect 10461 395 10471 549
rect 10511 395 10521 549
rect 10579 395 10589 549
rect 10629 395 10639 549
rect 10697 395 10707 549
rect 4804 342 4850 354
rect 4804 334 4810 342
rect 4844 334 4850 342
rect 4922 342 4968 354
rect 4922 334 4928 342
rect 4962 334 4968 342
rect 5040 342 5086 354
rect 5040 334 5046 342
rect 5080 334 5086 342
rect 5158 342 5204 354
rect 5158 334 5164 342
rect 5198 334 5204 342
rect 5276 342 5322 354
rect 5276 334 5282 342
rect 5316 334 5322 342
rect 5394 342 5440 354
rect 5394 334 5400 342
rect 5434 334 5440 342
rect 5512 342 5558 354
rect 5512 334 5518 342
rect 5552 334 5558 342
rect 5630 342 5676 354
rect 5630 334 5636 342
rect 5670 334 5676 342
rect 5748 342 5794 354
rect 5748 334 5754 342
rect 5788 334 5794 342
rect 5866 342 5912 354
rect 5866 334 5872 342
rect 5906 334 5912 342
rect 5984 342 6030 354
rect 5984 334 5990 342
rect 6024 334 6030 342
rect 6102 342 6148 354
rect 6102 334 6108 342
rect 6142 334 6148 342
rect 6220 342 6266 354
rect 6220 334 6226 342
rect 6260 334 6266 342
rect 6338 342 6384 354
rect 6338 334 6344 342
rect 6378 334 6384 342
rect 6456 342 6502 354
rect 6456 334 6462 342
rect 6496 334 6502 342
rect 6574 342 6620 354
rect 6574 334 6580 342
rect 6614 334 6620 342
rect 6692 342 6738 354
rect 6692 334 6698 342
rect 6732 334 6738 342
rect 6810 342 6856 354
rect 6810 334 6816 342
rect 6850 334 6856 342
rect 6928 342 6974 354
rect 6928 334 6934 342
rect 6968 334 6974 342
rect 7046 342 7092 354
rect 7046 334 7052 342
rect 7086 334 7092 342
rect 7164 342 7210 354
rect 7164 334 7170 342
rect 7204 334 7210 342
rect 7282 342 7328 354
rect 7282 334 7288 342
rect 7322 334 7328 342
rect 7400 342 7446 354
rect 7400 334 7406 342
rect 7440 334 7446 342
rect 7518 342 7564 354
rect 7518 334 7524 342
rect 7558 334 7564 342
rect 7636 342 7682 354
rect 7636 334 7642 342
rect 7676 334 7682 342
rect 7754 342 7800 354
rect 7754 334 7760 342
rect 7794 334 7800 342
rect 7872 342 7918 354
rect 7872 334 7878 342
rect 7912 334 7918 342
rect 7990 342 8036 354
rect 7990 334 7996 342
rect 8030 334 8036 342
rect 8108 342 8154 354
rect 8108 334 8114 342
rect 8148 334 8154 342
rect 8226 342 8272 354
rect 8226 334 8232 342
rect 8266 334 8272 342
rect 8344 342 8390 354
rect 8344 334 8350 342
rect 8384 334 8390 342
rect 8462 342 8508 354
rect 8462 334 8468 342
rect 8502 334 8508 342
rect 8580 342 8626 354
rect 8580 334 8586 342
rect 8620 334 8626 342
rect 8698 342 8744 354
rect 8698 334 8704 342
rect 8738 334 8744 342
rect 8816 342 8862 354
rect 8816 334 8822 342
rect 8856 334 8862 342
rect 8934 342 8980 354
rect 8934 334 8940 342
rect 8974 334 8980 342
rect 9052 342 9098 354
rect 9052 334 9058 342
rect 9092 334 9098 342
rect 9170 342 9216 354
rect 9170 334 9176 342
rect 9210 334 9216 342
rect 9288 342 9334 354
rect 9288 334 9294 342
rect 9328 334 9334 342
rect 9406 342 9452 354
rect 9406 334 9412 342
rect 9446 334 9452 342
rect 9524 342 9570 354
rect 9524 334 9530 342
rect 9564 334 9570 342
rect 9642 342 9688 354
rect 9642 334 9648 342
rect 9682 334 9688 342
rect 9760 342 9806 354
rect 9760 334 9766 342
rect 9800 334 9806 342
rect 9878 342 9924 354
rect 9878 334 9884 342
rect 9918 334 9924 342
rect 9996 342 10042 354
rect 9996 334 10002 342
rect 10036 334 10042 342
rect 10114 342 10160 354
rect 10114 334 10120 342
rect 10154 334 10160 342
rect 10232 342 10278 354
rect 10232 334 10238 342
rect 10272 334 10278 342
rect 10350 342 10396 354
rect 10350 334 10356 342
rect 10390 334 10396 342
rect 10468 342 10514 354
rect 10468 334 10474 342
rect 10508 334 10514 342
rect 10586 342 10632 354
rect 10586 334 10592 342
rect 10626 334 10632 342
rect 10704 342 10750 354
rect 10704 334 10710 342
rect 10744 334 10750 342
rect 4791 -226 4801 334
rect 4853 -226 4863 334
rect 4907 -226 4917 334
rect 4969 -226 4979 334
rect 5027 -226 5037 334
rect 5089 -226 5099 334
rect 5143 -226 5153 334
rect 5205 -226 5215 334
rect 5263 -226 5273 334
rect 5325 -226 5335 334
rect 5379 -226 5389 334
rect 5441 -226 5451 334
rect 5499 -226 5509 334
rect 5561 -226 5571 334
rect 5615 -226 5625 334
rect 5677 -226 5687 334
rect 5735 -226 5745 334
rect 5797 -226 5807 334
rect 5851 -226 5861 334
rect 5913 -226 5923 334
rect 5971 -226 5981 334
rect 6033 -226 6043 334
rect 6087 -226 6097 334
rect 6149 -226 6159 334
rect 6207 -226 6217 334
rect 6269 -226 6279 334
rect 6323 -226 6333 334
rect 6385 -226 6395 334
rect 6443 -226 6453 334
rect 6505 -226 6515 334
rect 6559 -226 6569 334
rect 6621 -226 6631 334
rect 6679 -226 6689 334
rect 6741 -226 6751 334
rect 6795 -226 6805 334
rect 6857 -226 6867 334
rect 6915 -226 6925 334
rect 6977 -226 6987 334
rect 7031 -226 7041 334
rect 7093 -226 7103 334
rect 7151 -226 7161 334
rect 7213 -226 7223 334
rect 7267 -226 7277 334
rect 7329 -226 7339 334
rect 7387 -226 7397 334
rect 7449 -226 7459 334
rect 7503 -226 7513 334
rect 7565 -226 7575 334
rect 7623 -226 7633 334
rect 7685 -226 7695 334
rect 7739 -226 7749 334
rect 7801 -226 7811 334
rect 7859 -226 7869 334
rect 7921 -226 7931 334
rect 7975 -226 7985 334
rect 8037 -226 8047 334
rect 8095 -226 8105 334
rect 8157 -226 8167 334
rect 8211 -226 8221 334
rect 8273 -226 8283 334
rect 8331 -226 8341 334
rect 8393 -226 8403 334
rect 8447 -226 8457 334
rect 8509 -226 8519 334
rect 8567 -226 8577 334
rect 8629 -226 8639 334
rect 8683 -226 8693 334
rect 8745 -226 8755 334
rect 8803 -226 8813 334
rect 8865 -226 8875 334
rect 8919 -226 8929 334
rect 8981 -226 8991 334
rect 9039 -226 9049 334
rect 9101 -226 9111 334
rect 9155 -226 9165 334
rect 9217 -226 9227 334
rect 9275 -226 9285 334
rect 9337 -226 9347 334
rect 9391 -226 9401 334
rect 9453 -226 9463 334
rect 9511 -226 9521 334
rect 9573 -226 9583 334
rect 9627 -226 9637 334
rect 9689 -226 9699 334
rect 9747 -226 9757 334
rect 9809 -226 9819 334
rect 9863 -226 9873 334
rect 9925 -226 9935 334
rect 9983 -226 9993 334
rect 10045 -226 10055 334
rect 10099 -226 10109 334
rect 10161 -226 10171 334
rect 10219 -226 10229 334
rect 10281 -226 10291 334
rect 10335 -226 10345 334
rect 10397 -226 10407 334
rect 10455 -226 10465 334
rect 10517 -226 10527 334
rect 10571 -226 10581 334
rect 10633 -226 10643 334
rect 10691 -226 10701 334
rect 10753 -226 10763 334
rect 4804 -234 4810 -226
rect 4844 -234 4850 -226
rect 4804 -246 4850 -234
rect 4922 -234 4928 -226
rect 4962 -234 4968 -226
rect 4922 -246 4968 -234
rect 5040 -234 5046 -226
rect 5080 -234 5086 -226
rect 5040 -246 5086 -234
rect 5158 -234 5164 -226
rect 5198 -234 5204 -226
rect 5158 -246 5204 -234
rect 5276 -234 5282 -226
rect 5316 -234 5322 -226
rect 5276 -246 5322 -234
rect 5394 -234 5400 -226
rect 5434 -234 5440 -226
rect 5394 -246 5440 -234
rect 5512 -234 5518 -226
rect 5552 -234 5558 -226
rect 5512 -246 5558 -234
rect 5630 -234 5636 -226
rect 5670 -234 5676 -226
rect 5630 -246 5676 -234
rect 5748 -234 5754 -226
rect 5788 -234 5794 -226
rect 5748 -246 5794 -234
rect 5866 -234 5872 -226
rect 5906 -234 5912 -226
rect 5866 -246 5912 -234
rect 5984 -234 5990 -226
rect 6024 -234 6030 -226
rect 5984 -246 6030 -234
rect 6102 -234 6108 -226
rect 6142 -234 6148 -226
rect 6102 -246 6148 -234
rect 6220 -234 6226 -226
rect 6260 -234 6266 -226
rect 6220 -246 6266 -234
rect 6338 -234 6344 -226
rect 6378 -234 6384 -226
rect 6338 -246 6384 -234
rect 6456 -234 6462 -226
rect 6496 -234 6502 -226
rect 6456 -246 6502 -234
rect 6574 -234 6580 -226
rect 6614 -234 6620 -226
rect 6574 -246 6620 -234
rect 6692 -234 6698 -226
rect 6732 -234 6738 -226
rect 6692 -246 6738 -234
rect 6810 -234 6816 -226
rect 6850 -234 6856 -226
rect 6810 -246 6856 -234
rect 6928 -234 6934 -226
rect 6968 -234 6974 -226
rect 6928 -246 6974 -234
rect 7046 -234 7052 -226
rect 7086 -234 7092 -226
rect 7046 -246 7092 -234
rect 7164 -234 7170 -226
rect 7204 -234 7210 -226
rect 7164 -246 7210 -234
rect 7282 -234 7288 -226
rect 7322 -234 7328 -226
rect 7282 -246 7328 -234
rect 7400 -234 7406 -226
rect 7440 -234 7446 -226
rect 7400 -246 7446 -234
rect 7518 -234 7524 -226
rect 7558 -234 7564 -226
rect 7518 -246 7564 -234
rect 7636 -234 7642 -226
rect 7676 -234 7682 -226
rect 7636 -246 7682 -234
rect 7754 -234 7760 -226
rect 7794 -234 7800 -226
rect 7754 -246 7800 -234
rect 7872 -234 7878 -226
rect 7912 -234 7918 -226
rect 7872 -246 7918 -234
rect 7990 -234 7996 -226
rect 8030 -234 8036 -226
rect 7990 -246 8036 -234
rect 8108 -234 8114 -226
rect 8148 -234 8154 -226
rect 8108 -246 8154 -234
rect 8226 -234 8232 -226
rect 8266 -234 8272 -226
rect 8226 -246 8272 -234
rect 8344 -234 8350 -226
rect 8384 -234 8390 -226
rect 8344 -246 8390 -234
rect 8462 -234 8468 -226
rect 8502 -234 8508 -226
rect 8462 -246 8508 -234
rect 8580 -234 8586 -226
rect 8620 -234 8626 -226
rect 8580 -246 8626 -234
rect 8698 -234 8704 -226
rect 8738 -234 8744 -226
rect 8698 -246 8744 -234
rect 8816 -234 8822 -226
rect 8856 -234 8862 -226
rect 8816 -246 8862 -234
rect 8934 -234 8940 -226
rect 8974 -234 8980 -226
rect 8934 -246 8980 -234
rect 9052 -234 9058 -226
rect 9092 -234 9098 -226
rect 9052 -246 9098 -234
rect 9170 -234 9176 -226
rect 9210 -234 9216 -226
rect 9170 -246 9216 -234
rect 9288 -234 9294 -226
rect 9328 -234 9334 -226
rect 9288 -246 9334 -234
rect 9406 -234 9412 -226
rect 9446 -234 9452 -226
rect 9406 -246 9452 -234
rect 9524 -234 9530 -226
rect 9564 -234 9570 -226
rect 9524 -246 9570 -234
rect 9642 -234 9648 -226
rect 9682 -234 9688 -226
rect 9642 -246 9688 -234
rect 9760 -234 9766 -226
rect 9800 -234 9806 -226
rect 9760 -246 9806 -234
rect 9878 -234 9884 -226
rect 9918 -234 9924 -226
rect 9878 -246 9924 -234
rect 9996 -234 10002 -226
rect 10036 -234 10042 -226
rect 9996 -246 10042 -234
rect 10114 -234 10120 -226
rect 10154 -234 10160 -226
rect 10114 -246 10160 -234
rect 10232 -234 10238 -226
rect 10272 -234 10278 -226
rect 10232 -246 10278 -234
rect 10350 -234 10356 -226
rect 10390 -234 10396 -226
rect 10350 -246 10396 -234
rect 10468 -234 10474 -226
rect 10508 -234 10514 -226
rect 10468 -246 10514 -234
rect 10586 -234 10592 -226
rect 10626 -234 10632 -226
rect 10586 -246 10632 -234
rect 10704 -234 10710 -226
rect 10744 -234 10750 -226
rect 10704 -246 10750 -234
rect 4746 -395 4801 -375
rect 4853 -395 5037 -375
rect 5089 -395 5273 -375
rect 5325 -395 5509 -375
rect 5561 -395 5745 -375
rect 5797 -395 5981 -375
rect 6033 -395 6217 -375
rect 6269 -395 6453 -375
rect 6505 -395 6689 -375
rect 6741 -395 6925 -375
rect 6977 -395 7161 -375
rect 7213 -395 7397 -375
rect 7449 -395 7633 -375
rect 7685 -395 7869 -375
rect 7921 -395 8105 -375
rect 8157 -395 8341 -375
rect 8393 -395 8577 -375
rect 8629 -395 8813 -375
rect 8865 -395 9049 -375
rect 9101 -395 9285 -375
rect 9337 -395 9521 -375
rect 9573 -395 9757 -375
rect 9809 -395 9993 -375
rect 10045 -395 10229 -375
rect 10281 -395 10465 -375
rect 10517 -395 10701 -375
rect 10753 -395 10794 -375
rect 4746 -429 4776 -395
rect 4882 -429 4920 -395
rect 4954 -429 4992 -395
rect 5026 -429 5037 -395
rect 5098 -429 5136 -395
rect 5170 -429 5208 -395
rect 5242 -429 5273 -395
rect 5325 -429 5352 -395
rect 5386 -429 5424 -395
rect 5458 -429 5496 -395
rect 5561 -429 5568 -395
rect 5602 -429 5640 -395
rect 5674 -429 5712 -395
rect 5818 -429 5856 -395
rect 5890 -429 5928 -395
rect 5962 -429 5981 -395
rect 6034 -429 6072 -395
rect 6106 -429 6144 -395
rect 6178 -429 6216 -395
rect 6269 -429 6288 -395
rect 6322 -429 6360 -395
rect 6394 -429 6432 -395
rect 6538 -429 6576 -395
rect 6610 -429 6648 -395
rect 6682 -429 6689 -395
rect 6754 -429 6792 -395
rect 6826 -429 6864 -395
rect 6898 -429 6925 -395
rect 6977 -429 7008 -395
rect 7042 -429 7080 -395
rect 7114 -429 7152 -395
rect 7213 -429 7224 -395
rect 7258 -429 7296 -395
rect 7330 -429 7368 -395
rect 7474 -429 7512 -395
rect 7546 -429 7584 -395
rect 7618 -429 7633 -395
rect 7690 -429 7728 -395
rect 7762 -429 7800 -395
rect 7834 -429 7869 -395
rect 7921 -429 7944 -395
rect 7978 -429 8016 -395
rect 8050 -429 8088 -395
rect 8157 -429 8160 -395
rect 8194 -429 8232 -395
rect 8266 -429 8304 -395
rect 8338 -429 8341 -395
rect 8410 -429 8448 -395
rect 8482 -429 8520 -395
rect 8554 -429 8577 -395
rect 8629 -429 8664 -395
rect 8698 -429 8736 -395
rect 8770 -429 8808 -395
rect 8865 -429 8880 -395
rect 8914 -429 8952 -395
rect 8986 -429 9024 -395
rect 9130 -429 9168 -395
rect 9202 -429 9240 -395
rect 9274 -429 9285 -395
rect 9346 -429 9384 -395
rect 9418 -429 9456 -395
rect 9490 -429 9521 -395
rect 9573 -429 9600 -395
rect 9634 -429 9672 -395
rect 9706 -429 9744 -395
rect 9809 -429 9816 -395
rect 9850 -429 9888 -395
rect 9922 -429 9960 -395
rect 10066 -429 10104 -395
rect 10138 -429 10176 -395
rect 10210 -429 10229 -395
rect 10282 -429 10320 -395
rect 10354 -429 10392 -395
rect 10426 -429 10464 -395
rect 10517 -429 10536 -395
rect 10570 -429 10608 -395
rect 10642 -429 10680 -395
rect 10786 -429 10794 -395
rect 4746 -483 4801 -429
rect 4853 -483 5037 -429
rect 5089 -483 5273 -429
rect 5325 -483 5509 -429
rect 5561 -483 5745 -429
rect 5797 -483 5981 -429
rect 6033 -483 6217 -429
rect 6269 -483 6453 -429
rect 6505 -483 6689 -429
rect 6741 -483 6925 -429
rect 6977 -483 7161 -429
rect 7213 -483 7397 -429
rect 7449 -483 7633 -429
rect 7685 -483 7869 -429
rect 7921 -483 8105 -429
rect 8157 -483 8341 -429
rect 8393 -483 8577 -429
rect 8629 -483 8813 -429
rect 8865 -483 9049 -429
rect 9101 -483 9285 -429
rect 9337 -483 9521 -429
rect 9573 -483 9757 -429
rect 9809 -483 9993 -429
rect 10045 -483 10229 -429
rect 10281 -483 10465 -429
rect 10517 -483 10701 -429
rect 10753 -483 10794 -429
rect 4746 -517 4776 -483
rect 4882 -517 4920 -483
rect 4954 -517 4992 -483
rect 5026 -517 5037 -483
rect 5098 -517 5136 -483
rect 5170 -517 5208 -483
rect 5242 -517 5273 -483
rect 5325 -517 5352 -483
rect 5386 -517 5424 -483
rect 5458 -517 5496 -483
rect 5561 -517 5568 -483
rect 5602 -517 5640 -483
rect 5674 -517 5712 -483
rect 5818 -517 5856 -483
rect 5890 -517 5928 -483
rect 5962 -517 5981 -483
rect 6034 -517 6072 -483
rect 6106 -517 6144 -483
rect 6178 -517 6216 -483
rect 6269 -517 6288 -483
rect 6322 -517 6360 -483
rect 6394 -517 6432 -483
rect 6538 -517 6576 -483
rect 6610 -517 6648 -483
rect 6682 -517 6689 -483
rect 6754 -517 6792 -483
rect 6826 -517 6864 -483
rect 6898 -517 6925 -483
rect 6977 -517 7008 -483
rect 7042 -517 7080 -483
rect 7114 -517 7152 -483
rect 7213 -517 7224 -483
rect 7258 -517 7296 -483
rect 7330 -517 7368 -483
rect 7474 -517 7512 -483
rect 7546 -517 7584 -483
rect 7618 -517 7633 -483
rect 7690 -517 7728 -483
rect 7762 -517 7800 -483
rect 7834 -517 7869 -483
rect 7921 -517 7944 -483
rect 7978 -517 8016 -483
rect 8050 -517 8088 -483
rect 8157 -517 8160 -483
rect 8194 -517 8232 -483
rect 8266 -517 8304 -483
rect 8338 -517 8341 -483
rect 8410 -517 8448 -483
rect 8482 -517 8520 -483
rect 8554 -517 8577 -483
rect 8629 -517 8664 -483
rect 8698 -517 8736 -483
rect 8770 -517 8808 -483
rect 8865 -517 8880 -483
rect 8914 -517 8952 -483
rect 8986 -517 9024 -483
rect 9130 -517 9168 -483
rect 9202 -517 9240 -483
rect 9274 -517 9285 -483
rect 9346 -517 9384 -483
rect 9418 -517 9456 -483
rect 9490 -517 9521 -483
rect 9573 -517 9600 -483
rect 9634 -517 9672 -483
rect 9706 -517 9744 -483
rect 9809 -517 9816 -483
rect 9850 -517 9888 -483
rect 9922 -517 9960 -483
rect 10066 -517 10104 -483
rect 10138 -517 10176 -483
rect 10210 -517 10229 -483
rect 10282 -517 10320 -483
rect 10354 -517 10392 -483
rect 10426 -517 10464 -483
rect 10517 -517 10536 -483
rect 10570 -517 10608 -483
rect 10642 -517 10680 -483
rect 10786 -517 10794 -483
rect 4746 -571 4801 -517
rect 4853 -571 5037 -517
rect 5089 -571 5273 -517
rect 5325 -571 5509 -517
rect 5561 -571 5745 -517
rect 5797 -571 5981 -517
rect 6033 -571 6217 -517
rect 6269 -571 6453 -517
rect 6505 -571 6689 -517
rect 6741 -571 6925 -517
rect 6977 -571 7161 -517
rect 7213 -571 7397 -517
rect 7449 -571 7633 -517
rect 7685 -571 7869 -517
rect 7921 -571 8105 -517
rect 8157 -571 8341 -517
rect 8393 -571 8577 -517
rect 8629 -571 8813 -517
rect 8865 -571 9049 -517
rect 9101 -571 9285 -517
rect 9337 -571 9521 -517
rect 9573 -571 9757 -517
rect 9809 -571 9993 -517
rect 10045 -571 10229 -517
rect 10281 -571 10465 -517
rect 10517 -571 10701 -517
rect 10753 -571 10794 -517
rect 4746 -605 4776 -571
rect 4882 -605 4920 -571
rect 4954 -605 4992 -571
rect 5026 -605 5037 -571
rect 5098 -605 5136 -571
rect 5170 -605 5208 -571
rect 5242 -605 5273 -571
rect 5325 -605 5352 -571
rect 5386 -605 5424 -571
rect 5458 -605 5496 -571
rect 5561 -605 5568 -571
rect 5602 -605 5640 -571
rect 5674 -605 5712 -571
rect 5818 -605 5856 -571
rect 5890 -605 5928 -571
rect 5962 -605 5981 -571
rect 6034 -605 6072 -571
rect 6106 -605 6144 -571
rect 6178 -605 6216 -571
rect 6269 -605 6288 -571
rect 6322 -605 6360 -571
rect 6394 -605 6432 -571
rect 6538 -605 6576 -571
rect 6610 -605 6648 -571
rect 6682 -605 6689 -571
rect 6754 -605 6792 -571
rect 6826 -605 6864 -571
rect 6898 -605 6925 -571
rect 6977 -605 7008 -571
rect 7042 -605 7080 -571
rect 7114 -605 7152 -571
rect 7213 -605 7224 -571
rect 7258 -605 7296 -571
rect 7330 -605 7368 -571
rect 7474 -605 7512 -571
rect 7546 -605 7584 -571
rect 7618 -605 7633 -571
rect 7690 -605 7728 -571
rect 7762 -605 7800 -571
rect 7834 -605 7869 -571
rect 7921 -605 7944 -571
rect 7978 -605 8016 -571
rect 8050 -605 8088 -571
rect 8157 -605 8160 -571
rect 8194 -605 8232 -571
rect 8266 -605 8304 -571
rect 8338 -605 8341 -571
rect 8410 -605 8448 -571
rect 8482 -605 8520 -571
rect 8554 -605 8577 -571
rect 8629 -605 8664 -571
rect 8698 -605 8736 -571
rect 8770 -605 8808 -571
rect 8865 -605 8880 -571
rect 8914 -605 8952 -571
rect 8986 -605 9024 -571
rect 9130 -605 9168 -571
rect 9202 -605 9240 -571
rect 9274 -605 9285 -571
rect 9346 -605 9384 -571
rect 9418 -605 9456 -571
rect 9490 -605 9521 -571
rect 9573 -605 9600 -571
rect 9634 -605 9672 -571
rect 9706 -605 9744 -571
rect 9809 -605 9816 -571
rect 9850 -605 9888 -571
rect 9922 -605 9960 -571
rect 10066 -605 10104 -571
rect 10138 -605 10176 -571
rect 10210 -605 10229 -571
rect 10282 -605 10320 -571
rect 10354 -605 10392 -571
rect 10426 -605 10464 -571
rect 10517 -605 10536 -571
rect 10570 -605 10608 -571
rect 10642 -605 10680 -571
rect 10786 -605 10794 -571
rect 4746 -625 4801 -605
rect 4853 -625 5037 -605
rect 5089 -625 5273 -605
rect 5325 -625 5509 -605
rect 5561 -625 5745 -605
rect 5797 -625 5981 -605
rect 6033 -625 6217 -605
rect 6269 -625 6453 -605
rect 6505 -625 6689 -605
rect 6741 -625 6925 -605
rect 6977 -625 7161 -605
rect 7213 -625 7397 -605
rect 7449 -625 7633 -605
rect 7685 -625 7869 -605
rect 7921 -625 8105 -605
rect 8157 -625 8341 -605
rect 8393 -625 8577 -605
rect 8629 -625 8813 -605
rect 8865 -625 9049 -605
rect 9101 -625 9285 -605
rect 9337 -625 9521 -605
rect 9573 -625 9757 -605
rect 9809 -625 9993 -605
rect 10045 -625 10229 -605
rect 10281 -625 10465 -605
rect 10517 -625 10701 -605
rect 10753 -625 10794 -605
rect 4804 -872 4850 -860
rect 4804 -880 4810 -872
rect 4844 -880 4850 -872
rect 4922 -872 4968 -860
rect 4922 -880 4928 -872
rect 4962 -880 4968 -872
rect 5040 -872 5086 -860
rect 5040 -880 5046 -872
rect 5080 -880 5086 -872
rect 5158 -872 5204 -860
rect 5394 -872 5440 -860
rect 5630 -872 5676 -860
rect 5866 -872 5912 -860
rect 6102 -872 6148 -860
rect 6338 -872 6384 -860
rect 6574 -872 6620 -860
rect 6810 -872 6856 -860
rect 7046 -872 7092 -860
rect 7282 -872 7328 -860
rect 7518 -872 7564 -860
rect 7754 -872 7800 -860
rect 7990 -872 8036 -860
rect 8226 -872 8272 -860
rect 8462 -872 8508 -860
rect 8698 -872 8744 -860
rect 8934 -872 8980 -860
rect 9170 -872 9216 -860
rect 9406 -872 9452 -860
rect 9642 -872 9688 -860
rect 9878 -872 9924 -860
rect 10114 -872 10160 -860
rect 10350 -872 10396 -860
rect 10586 -872 10632 -860
rect 5158 -880 5164 -872
rect 5198 -880 5204 -872
rect 5394 -880 5400 -872
rect 5434 -880 5440 -872
rect 5630 -880 5636 -872
rect 5670 -880 5676 -872
rect 5866 -880 5872 -872
rect 5906 -880 5912 -872
rect 6102 -880 6108 -872
rect 6142 -880 6148 -872
rect 6338 -880 6344 -872
rect 6378 -880 6384 -872
rect 6574 -880 6580 -872
rect 6614 -880 6620 -872
rect 6810 -880 6816 -872
rect 6850 -880 6856 -872
rect 7046 -880 7052 -872
rect 7086 -880 7092 -872
rect 7282 -880 7288 -872
rect 7322 -880 7328 -872
rect 7518 -880 7524 -872
rect 7558 -880 7564 -872
rect 7754 -880 7760 -872
rect 7794 -880 7800 -872
rect 7990 -880 7996 -872
rect 8030 -880 8036 -872
rect 8226 -880 8232 -872
rect 8266 -880 8272 -872
rect 8462 -880 8468 -872
rect 8502 -880 8508 -872
rect 8698 -880 8704 -872
rect 8738 -880 8744 -872
rect 8934 -880 8940 -872
rect 8974 -880 8980 -872
rect 9170 -880 9176 -872
rect 9210 -880 9216 -872
rect 9406 -880 9412 -872
rect 9446 -880 9452 -872
rect 9642 -880 9648 -872
rect 9682 -880 9688 -872
rect 9878 -880 9884 -872
rect 9918 -880 9924 -872
rect 10114 -880 10120 -872
rect 10154 -880 10160 -872
rect 10350 -880 10356 -872
rect 10390 -880 10396 -872
rect 10586 -880 10592 -872
rect 10626 -880 10632 -872
rect 4791 -1440 4801 -880
rect 4853 -1440 4863 -880
rect 4907 -1440 4917 -880
rect 4969 -1440 4979 -880
rect 5027 -1440 5037 -880
rect 5089 -1440 5099 -880
rect 5143 -1440 5153 -880
rect 5205 -1440 5215 -880
rect 5263 -1440 5273 -880
rect 5325 -1440 5335 -880
rect 5379 -1440 5389 -880
rect 5441 -1440 5451 -880
rect 5499 -1440 5509 -880
rect 5561 -1440 5571 -880
rect 5615 -1440 5625 -880
rect 5677 -1440 5687 -880
rect 5735 -1440 5745 -880
rect 5797 -1440 5807 -880
rect 5851 -1440 5861 -880
rect 5913 -1440 5923 -880
rect 5971 -1440 5981 -880
rect 6033 -1440 6043 -880
rect 6087 -1440 6097 -880
rect 6149 -1440 6159 -880
rect 6207 -1440 6217 -880
rect 6269 -1440 6279 -880
rect 6323 -1440 6333 -880
rect 6385 -1440 6395 -880
rect 6443 -1440 6453 -880
rect 6505 -1440 6515 -880
rect 6559 -1440 6569 -880
rect 6621 -1440 6631 -880
rect 6679 -1440 6689 -880
rect 6741 -1440 6751 -880
rect 6795 -1440 6805 -880
rect 6857 -1440 6867 -880
rect 6915 -1440 6925 -880
rect 6977 -1440 6987 -880
rect 7031 -1440 7041 -880
rect 7093 -1440 7103 -880
rect 7151 -1440 7161 -880
rect 7213 -1440 7223 -880
rect 7267 -1440 7277 -880
rect 7329 -1440 7339 -880
rect 7387 -1440 7397 -880
rect 7449 -1440 7459 -880
rect 7503 -1440 7513 -880
rect 7565 -1440 7575 -880
rect 7623 -1440 7633 -880
rect 7685 -1440 7695 -880
rect 7739 -1440 7749 -880
rect 7801 -1440 7811 -880
rect 7859 -1440 7869 -880
rect 7921 -1440 7931 -880
rect 7975 -1440 7985 -880
rect 8037 -1440 8047 -880
rect 8095 -1440 8105 -880
rect 8157 -1440 8167 -880
rect 8211 -1440 8221 -880
rect 8273 -1440 8283 -880
rect 8331 -1440 8341 -880
rect 8393 -1440 8403 -880
rect 8447 -1440 8457 -880
rect 8509 -1440 8519 -880
rect 8567 -1440 8577 -880
rect 8629 -1440 8639 -880
rect 8683 -1440 8693 -880
rect 8745 -1440 8755 -880
rect 8803 -1440 8813 -880
rect 8865 -1440 8875 -880
rect 8919 -1440 8929 -880
rect 8981 -1440 8991 -880
rect 9039 -1440 9049 -880
rect 9101 -1440 9111 -880
rect 9155 -1440 9165 -880
rect 9217 -1440 9227 -880
rect 9275 -1440 9285 -880
rect 9337 -1440 9347 -880
rect 9391 -1440 9401 -880
rect 9453 -1440 9463 -880
rect 9511 -1440 9521 -880
rect 9573 -1440 9583 -880
rect 9627 -1440 9637 -880
rect 9689 -1440 9699 -880
rect 9747 -1440 9757 -880
rect 9809 -1440 9819 -880
rect 9863 -1440 9873 -880
rect 9925 -1440 9935 -880
rect 9983 -1440 9993 -880
rect 10045 -1440 10055 -880
rect 10099 -1440 10109 -880
rect 10161 -1440 10171 -880
rect 10219 -1440 10229 -880
rect 10281 -1440 10291 -880
rect 10335 -1440 10345 -880
rect 10397 -1440 10407 -880
rect 10455 -1440 10465 -880
rect 10517 -1440 10527 -880
rect 10571 -1440 10581 -880
rect 10633 -1440 10643 -880
rect 10691 -1440 10701 -880
rect 10753 -1440 10763 -880
rect 4804 -1448 4810 -1440
rect 4844 -1448 4850 -1440
rect 4804 -1460 4850 -1448
rect 4922 -1448 4928 -1440
rect 4962 -1448 4968 -1440
rect 4922 -1460 4968 -1448
rect 5040 -1448 5046 -1440
rect 5080 -1448 5086 -1440
rect 5040 -1460 5086 -1448
rect 5158 -1448 5164 -1440
rect 5198 -1448 5204 -1440
rect 5158 -1460 5204 -1448
rect 5276 -1448 5282 -1440
rect 5316 -1448 5322 -1440
rect 5276 -1460 5322 -1448
rect 5394 -1448 5400 -1440
rect 5434 -1448 5440 -1440
rect 5394 -1460 5440 -1448
rect 5512 -1448 5518 -1440
rect 5552 -1448 5558 -1440
rect 5512 -1460 5558 -1448
rect 5630 -1448 5636 -1440
rect 5670 -1448 5676 -1440
rect 5630 -1460 5676 -1448
rect 5748 -1448 5754 -1440
rect 5788 -1448 5794 -1440
rect 5748 -1460 5794 -1448
rect 5866 -1448 5872 -1440
rect 5906 -1448 5912 -1440
rect 5866 -1460 5912 -1448
rect 5984 -1448 5990 -1440
rect 6024 -1448 6030 -1440
rect 5984 -1460 6030 -1448
rect 6102 -1448 6108 -1440
rect 6142 -1448 6148 -1440
rect 6102 -1460 6148 -1448
rect 6220 -1448 6226 -1440
rect 6260 -1448 6266 -1440
rect 6220 -1460 6266 -1448
rect 6338 -1448 6344 -1440
rect 6378 -1448 6384 -1440
rect 6338 -1460 6384 -1448
rect 6456 -1448 6462 -1440
rect 6496 -1448 6502 -1440
rect 6456 -1460 6502 -1448
rect 6574 -1448 6580 -1440
rect 6614 -1448 6620 -1440
rect 6574 -1460 6620 -1448
rect 6692 -1448 6698 -1440
rect 6732 -1448 6738 -1440
rect 6692 -1460 6738 -1448
rect 6810 -1448 6816 -1440
rect 6850 -1448 6856 -1440
rect 6810 -1460 6856 -1448
rect 6928 -1448 6934 -1440
rect 6968 -1448 6974 -1440
rect 6928 -1460 6974 -1448
rect 7046 -1448 7052 -1440
rect 7086 -1448 7092 -1440
rect 7046 -1460 7092 -1448
rect 7164 -1448 7170 -1440
rect 7204 -1448 7210 -1440
rect 7164 -1460 7210 -1448
rect 7282 -1448 7288 -1440
rect 7322 -1448 7328 -1440
rect 7282 -1460 7328 -1448
rect 7400 -1448 7406 -1440
rect 7440 -1448 7446 -1440
rect 7400 -1460 7446 -1448
rect 7518 -1448 7524 -1440
rect 7558 -1448 7564 -1440
rect 7518 -1460 7564 -1448
rect 7636 -1448 7642 -1440
rect 7676 -1448 7682 -1440
rect 7636 -1460 7682 -1448
rect 7754 -1448 7760 -1440
rect 7794 -1448 7800 -1440
rect 7754 -1460 7800 -1448
rect 7872 -1448 7878 -1440
rect 7912 -1448 7918 -1440
rect 7872 -1460 7918 -1448
rect 7990 -1448 7996 -1440
rect 8030 -1448 8036 -1440
rect 7990 -1460 8036 -1448
rect 8108 -1448 8114 -1440
rect 8148 -1448 8154 -1440
rect 8108 -1460 8154 -1448
rect 8226 -1448 8232 -1440
rect 8266 -1448 8272 -1440
rect 8226 -1460 8272 -1448
rect 8344 -1448 8350 -1440
rect 8384 -1448 8390 -1440
rect 8344 -1460 8390 -1448
rect 8462 -1448 8468 -1440
rect 8502 -1448 8508 -1440
rect 8462 -1460 8508 -1448
rect 8580 -1448 8586 -1440
rect 8620 -1448 8626 -1440
rect 8580 -1460 8626 -1448
rect 8698 -1448 8704 -1440
rect 8738 -1448 8744 -1440
rect 8698 -1460 8744 -1448
rect 8816 -1448 8822 -1440
rect 8856 -1448 8862 -1440
rect 8816 -1460 8862 -1448
rect 8934 -1448 8940 -1440
rect 8974 -1448 8980 -1440
rect 8934 -1460 8980 -1448
rect 9052 -1448 9058 -1440
rect 9092 -1448 9098 -1440
rect 9052 -1460 9098 -1448
rect 9170 -1448 9176 -1440
rect 9210 -1448 9216 -1440
rect 9170 -1460 9216 -1448
rect 9288 -1448 9294 -1440
rect 9328 -1448 9334 -1440
rect 9288 -1460 9334 -1448
rect 9406 -1448 9412 -1440
rect 9446 -1448 9452 -1440
rect 9406 -1460 9452 -1448
rect 9524 -1448 9530 -1440
rect 9564 -1448 9570 -1440
rect 9524 -1460 9570 -1448
rect 9642 -1448 9648 -1440
rect 9682 -1448 9688 -1440
rect 9642 -1460 9688 -1448
rect 9760 -1448 9766 -1440
rect 9800 -1448 9806 -1440
rect 9760 -1460 9806 -1448
rect 9878 -1448 9884 -1440
rect 9918 -1448 9924 -1440
rect 9878 -1460 9924 -1448
rect 9996 -1448 10002 -1440
rect 10036 -1448 10042 -1440
rect 9996 -1460 10042 -1448
rect 10114 -1448 10120 -1440
rect 10154 -1448 10160 -1440
rect 10114 -1460 10160 -1448
rect 10232 -1448 10238 -1440
rect 10272 -1448 10278 -1440
rect 10232 -1460 10278 -1448
rect 10350 -1448 10356 -1440
rect 10390 -1448 10396 -1440
rect 10350 -1460 10396 -1448
rect 10468 -1448 10474 -1440
rect 10508 -1448 10514 -1440
rect 10468 -1460 10514 -1448
rect 10586 -1448 10592 -1440
rect 10626 -1448 10632 -1440
rect 10586 -1460 10632 -1448
rect 10704 -1448 10710 -1440
rect 10744 -1448 10750 -1440
rect 10704 -1460 10750 -1448
rect 4847 -1655 4857 -1501
rect 4915 -1655 4925 -1501
rect 4965 -1655 4975 -1501
rect 5033 -1655 5043 -1501
rect 5083 -1655 5093 -1501
rect 5151 -1655 5161 -1501
rect 5201 -1655 5211 -1501
rect 5269 -1655 5279 -1501
rect 5319 -1655 5329 -1501
rect 5387 -1655 5397 -1501
rect 5437 -1655 5447 -1501
rect 5505 -1655 5515 -1501
rect 5555 -1655 5565 -1501
rect 5623 -1655 5633 -1501
rect 5673 -1655 5683 -1501
rect 5741 -1655 5751 -1501
rect 5791 -1655 5801 -1501
rect 5859 -1655 5869 -1501
rect 5909 -1655 5919 -1501
rect 5977 -1655 5987 -1501
rect 6027 -1655 6037 -1501
rect 6095 -1655 6105 -1501
rect 6145 -1655 6155 -1501
rect 6213 -1655 6223 -1501
rect 6263 -1655 6273 -1501
rect 6331 -1655 6341 -1501
rect 6381 -1655 6391 -1501
rect 6449 -1655 6459 -1501
rect 6499 -1655 6509 -1501
rect 6567 -1655 6577 -1501
rect 6617 -1655 6627 -1501
rect 6685 -1655 6695 -1501
rect 6735 -1655 6745 -1501
rect 6803 -1655 6813 -1501
rect 6853 -1655 6863 -1501
rect 6921 -1655 6931 -1501
rect 6971 -1655 6981 -1501
rect 7039 -1655 7049 -1501
rect 7089 -1655 7099 -1501
rect 7157 -1655 7167 -1501
rect 7207 -1655 7217 -1501
rect 7275 -1655 7285 -1501
rect 7325 -1655 7335 -1501
rect 7393 -1655 7403 -1501
rect 7443 -1655 7453 -1501
rect 7511 -1655 7521 -1501
rect 7561 -1655 7571 -1501
rect 7629 -1655 7639 -1501
rect 7679 -1655 7689 -1501
rect 7747 -1655 7757 -1501
rect 7797 -1655 7807 -1501
rect 7865 -1655 7875 -1501
rect 7915 -1655 7925 -1501
rect 7983 -1655 7993 -1501
rect 8033 -1655 8043 -1501
rect 8101 -1655 8111 -1501
rect 8151 -1655 8161 -1501
rect 8219 -1655 8229 -1501
rect 8269 -1655 8279 -1501
rect 8337 -1655 8347 -1501
rect 8387 -1655 8397 -1501
rect 8455 -1655 8465 -1501
rect 8505 -1655 8515 -1501
rect 8573 -1655 8583 -1501
rect 8623 -1655 8633 -1501
rect 8691 -1655 8701 -1501
rect 8741 -1655 8751 -1501
rect 8809 -1655 8819 -1501
rect 8859 -1655 8869 -1501
rect 8927 -1655 8937 -1501
rect 8977 -1655 8987 -1501
rect 9045 -1655 9055 -1501
rect 9095 -1655 9105 -1501
rect 9163 -1655 9173 -1501
rect 9213 -1655 9223 -1501
rect 9281 -1655 9291 -1501
rect 9331 -1655 9341 -1501
rect 9399 -1655 9409 -1501
rect 9449 -1655 9459 -1501
rect 9517 -1655 9527 -1501
rect 9567 -1655 9577 -1501
rect 9635 -1655 9645 -1501
rect 9685 -1655 9695 -1501
rect 9753 -1655 9763 -1501
rect 9803 -1655 9813 -1501
rect 9871 -1655 9881 -1501
rect 9921 -1655 9931 -1501
rect 9989 -1655 9999 -1501
rect 10039 -1655 10049 -1501
rect 10107 -1655 10117 -1501
rect 10157 -1655 10167 -1501
rect 10225 -1655 10235 -1501
rect 10275 -1655 10285 -1501
rect 10343 -1655 10353 -1501
rect 10393 -1655 10403 -1501
rect 10461 -1655 10471 -1501
rect 10511 -1655 10521 -1501
rect 10579 -1655 10589 -1501
rect 10629 -1655 10639 -1501
rect 10697 -1655 10707 -1501
rect 4804 -1708 4850 -1696
rect 4804 -1716 4810 -1708
rect 4844 -1716 4850 -1708
rect 4922 -1708 4968 -1696
rect 4922 -1716 4928 -1708
rect 4962 -1716 4968 -1708
rect 5040 -1708 5086 -1696
rect 5040 -1716 5046 -1708
rect 5080 -1716 5086 -1708
rect 5158 -1708 5204 -1696
rect 5158 -1716 5164 -1708
rect 5198 -1716 5204 -1708
rect 5276 -1708 5322 -1696
rect 5276 -1716 5282 -1708
rect 5316 -1716 5322 -1708
rect 5394 -1708 5440 -1696
rect 5394 -1716 5400 -1708
rect 5434 -1716 5440 -1708
rect 5512 -1708 5558 -1696
rect 5512 -1716 5518 -1708
rect 5552 -1716 5558 -1708
rect 5630 -1708 5676 -1696
rect 5630 -1716 5636 -1708
rect 5670 -1716 5676 -1708
rect 5748 -1708 5794 -1696
rect 5748 -1716 5754 -1708
rect 5788 -1716 5794 -1708
rect 5866 -1708 5912 -1696
rect 5866 -1716 5872 -1708
rect 5906 -1716 5912 -1708
rect 5984 -1708 6030 -1696
rect 5984 -1716 5990 -1708
rect 6024 -1716 6030 -1708
rect 6102 -1708 6148 -1696
rect 6102 -1716 6108 -1708
rect 6142 -1716 6148 -1708
rect 6220 -1708 6266 -1696
rect 6220 -1716 6226 -1708
rect 6260 -1716 6266 -1708
rect 6338 -1708 6384 -1696
rect 6338 -1716 6344 -1708
rect 6378 -1716 6384 -1708
rect 6456 -1708 6502 -1696
rect 6456 -1716 6462 -1708
rect 6496 -1716 6502 -1708
rect 6574 -1708 6620 -1696
rect 6574 -1716 6580 -1708
rect 6614 -1716 6620 -1708
rect 6692 -1708 6738 -1696
rect 6692 -1716 6698 -1708
rect 6732 -1716 6738 -1708
rect 6810 -1708 6856 -1696
rect 6810 -1716 6816 -1708
rect 6850 -1716 6856 -1708
rect 6928 -1708 6974 -1696
rect 6928 -1716 6934 -1708
rect 6968 -1716 6974 -1708
rect 7046 -1708 7092 -1696
rect 7046 -1716 7052 -1708
rect 7086 -1716 7092 -1708
rect 7164 -1708 7210 -1696
rect 7164 -1716 7170 -1708
rect 7204 -1716 7210 -1708
rect 7282 -1708 7328 -1696
rect 7282 -1716 7288 -1708
rect 7322 -1716 7328 -1708
rect 7400 -1708 7446 -1696
rect 7400 -1716 7406 -1708
rect 7440 -1716 7446 -1708
rect 7518 -1708 7564 -1696
rect 7518 -1716 7524 -1708
rect 7558 -1716 7564 -1708
rect 7636 -1708 7682 -1696
rect 7636 -1716 7642 -1708
rect 7676 -1716 7682 -1708
rect 7754 -1708 7800 -1696
rect 7754 -1716 7760 -1708
rect 7794 -1716 7800 -1708
rect 7872 -1708 7918 -1696
rect 7872 -1716 7878 -1708
rect 7912 -1716 7918 -1708
rect 7990 -1708 8036 -1696
rect 7990 -1716 7996 -1708
rect 8030 -1716 8036 -1708
rect 8108 -1708 8154 -1696
rect 8108 -1716 8114 -1708
rect 8148 -1716 8154 -1708
rect 8226 -1708 8272 -1696
rect 8226 -1716 8232 -1708
rect 8266 -1716 8272 -1708
rect 8344 -1708 8390 -1696
rect 8344 -1716 8350 -1708
rect 8384 -1716 8390 -1708
rect 8462 -1708 8508 -1696
rect 8462 -1716 8468 -1708
rect 8502 -1716 8508 -1708
rect 8580 -1708 8626 -1696
rect 8580 -1716 8586 -1708
rect 8620 -1716 8626 -1708
rect 8698 -1708 8744 -1696
rect 8698 -1716 8704 -1708
rect 8738 -1716 8744 -1708
rect 8816 -1708 8862 -1696
rect 8816 -1716 8822 -1708
rect 8856 -1716 8862 -1708
rect 8934 -1708 8980 -1696
rect 8934 -1716 8940 -1708
rect 8974 -1716 8980 -1708
rect 9052 -1708 9098 -1696
rect 9052 -1716 9058 -1708
rect 9092 -1716 9098 -1708
rect 9170 -1708 9216 -1696
rect 9170 -1716 9176 -1708
rect 9210 -1716 9216 -1708
rect 9288 -1708 9334 -1696
rect 9288 -1716 9294 -1708
rect 9328 -1716 9334 -1708
rect 9406 -1708 9452 -1696
rect 9406 -1716 9412 -1708
rect 9446 -1716 9452 -1708
rect 9524 -1708 9570 -1696
rect 9524 -1716 9530 -1708
rect 9564 -1716 9570 -1708
rect 9642 -1708 9688 -1696
rect 9642 -1716 9648 -1708
rect 9682 -1716 9688 -1708
rect 9760 -1708 9806 -1696
rect 9760 -1716 9766 -1708
rect 9800 -1716 9806 -1708
rect 9878 -1708 9924 -1696
rect 9878 -1716 9884 -1708
rect 9918 -1716 9924 -1708
rect 9996 -1708 10042 -1696
rect 9996 -1716 10002 -1708
rect 10036 -1716 10042 -1708
rect 10114 -1708 10160 -1696
rect 10114 -1716 10120 -1708
rect 10154 -1716 10160 -1708
rect 10232 -1708 10278 -1696
rect 10232 -1716 10238 -1708
rect 10272 -1716 10278 -1708
rect 10350 -1708 10396 -1696
rect 10350 -1716 10356 -1708
rect 10390 -1716 10396 -1708
rect 10468 -1708 10514 -1696
rect 10468 -1716 10474 -1708
rect 10508 -1716 10514 -1708
rect 10586 -1708 10632 -1696
rect 10586 -1716 10592 -1708
rect 10626 -1716 10632 -1708
rect 10704 -1708 10750 -1696
rect 10704 -1716 10710 -1708
rect 10744 -1716 10750 -1708
rect 4791 -2276 4801 -1716
rect 4853 -2276 4863 -1716
rect 4907 -2276 4917 -1716
rect 4969 -2276 4979 -1716
rect 5027 -2276 5037 -1716
rect 5089 -2276 5099 -1716
rect 5143 -2276 5153 -1716
rect 5205 -2276 5215 -1716
rect 5263 -2276 5273 -1716
rect 5325 -2276 5335 -1716
rect 5379 -2276 5389 -1716
rect 5441 -2276 5451 -1716
rect 5499 -2276 5509 -1716
rect 5561 -2276 5571 -1716
rect 5615 -2276 5625 -1716
rect 5677 -2276 5687 -1716
rect 5735 -2276 5745 -1716
rect 5797 -2276 5807 -1716
rect 5851 -2276 5861 -1716
rect 5913 -2276 5923 -1716
rect 5971 -2276 5981 -1716
rect 6033 -2276 6043 -1716
rect 6087 -2276 6097 -1716
rect 6149 -2276 6159 -1716
rect 6207 -2276 6217 -1716
rect 6269 -2276 6279 -1716
rect 6323 -2276 6333 -1716
rect 6385 -2276 6395 -1716
rect 6443 -2276 6453 -1716
rect 6505 -2276 6515 -1716
rect 6559 -2276 6569 -1716
rect 6621 -2276 6631 -1716
rect 6679 -2276 6689 -1716
rect 6741 -2276 6751 -1716
rect 6795 -2276 6805 -1716
rect 6857 -2276 6867 -1716
rect 6915 -2276 6925 -1716
rect 6977 -2276 6987 -1716
rect 7031 -2276 7041 -1716
rect 7093 -2276 7103 -1716
rect 7151 -2276 7161 -1716
rect 7213 -2276 7223 -1716
rect 7267 -2276 7277 -1716
rect 7329 -2276 7339 -1716
rect 7387 -2276 7397 -1716
rect 7449 -2276 7459 -1716
rect 7503 -2276 7513 -1716
rect 7565 -2276 7575 -1716
rect 7623 -2276 7633 -1716
rect 7685 -2276 7695 -1716
rect 7739 -2276 7749 -1716
rect 7801 -2276 7811 -1716
rect 7859 -2276 7869 -1716
rect 7921 -2276 7931 -1716
rect 7975 -2276 7985 -1716
rect 8037 -2276 8047 -1716
rect 8095 -2276 8105 -1716
rect 8157 -2276 8167 -1716
rect 8211 -2276 8221 -1716
rect 8273 -2276 8283 -1716
rect 8331 -2276 8341 -1716
rect 8393 -2276 8403 -1716
rect 8447 -2276 8457 -1716
rect 8509 -2276 8519 -1716
rect 8567 -2276 8577 -1716
rect 8629 -2276 8639 -1716
rect 8683 -2276 8693 -1716
rect 8745 -2276 8755 -1716
rect 8803 -2276 8813 -1716
rect 8865 -2276 8875 -1716
rect 8919 -2276 8929 -1716
rect 8981 -2276 8991 -1716
rect 9039 -2276 9049 -1716
rect 9101 -2276 9111 -1716
rect 9155 -2276 9165 -1716
rect 9217 -2276 9227 -1716
rect 9275 -2276 9285 -1716
rect 9337 -2276 9347 -1716
rect 9391 -2276 9401 -1716
rect 9453 -2276 9463 -1716
rect 9511 -2276 9521 -1716
rect 9573 -2276 9583 -1716
rect 9627 -2276 9637 -1716
rect 9689 -2276 9699 -1716
rect 9747 -2276 9757 -1716
rect 9809 -2276 9819 -1716
rect 9863 -2276 9873 -1716
rect 9925 -2276 9935 -1716
rect 9983 -2276 9993 -1716
rect 10045 -2276 10055 -1716
rect 10099 -2276 10109 -1716
rect 10161 -2276 10171 -1716
rect 10219 -2276 10229 -1716
rect 10281 -2276 10291 -1716
rect 10335 -2276 10345 -1716
rect 10397 -2276 10407 -1716
rect 10455 -2276 10465 -1716
rect 10517 -2276 10527 -1716
rect 10571 -2276 10581 -1716
rect 10633 -2276 10643 -1716
rect 10691 -2276 10701 -1716
rect 10753 -2276 10763 -1716
rect 4804 -2284 4810 -2276
rect 4844 -2284 4850 -2276
rect 4804 -2296 4850 -2284
rect 4922 -2284 4928 -2276
rect 4962 -2284 4968 -2276
rect 4922 -2296 4968 -2284
rect 5040 -2284 5046 -2276
rect 5080 -2284 5086 -2276
rect 5040 -2296 5086 -2284
rect 5158 -2284 5164 -2276
rect 5198 -2284 5204 -2276
rect 5158 -2296 5204 -2284
rect 5276 -2284 5282 -2276
rect 5316 -2284 5322 -2276
rect 5276 -2296 5322 -2284
rect 5394 -2284 5400 -2276
rect 5434 -2284 5440 -2276
rect 5394 -2296 5440 -2284
rect 5512 -2284 5518 -2276
rect 5552 -2284 5558 -2276
rect 5512 -2296 5558 -2284
rect 5630 -2284 5636 -2276
rect 5670 -2284 5676 -2276
rect 5630 -2296 5676 -2284
rect 5748 -2284 5754 -2276
rect 5788 -2284 5794 -2276
rect 5748 -2296 5794 -2284
rect 5866 -2284 5872 -2276
rect 5906 -2284 5912 -2276
rect 5866 -2296 5912 -2284
rect 5984 -2284 5990 -2276
rect 6024 -2284 6030 -2276
rect 5984 -2296 6030 -2284
rect 6102 -2284 6108 -2276
rect 6142 -2284 6148 -2276
rect 6102 -2296 6148 -2284
rect 6220 -2284 6226 -2276
rect 6260 -2284 6266 -2276
rect 6220 -2296 6266 -2284
rect 6338 -2284 6344 -2276
rect 6378 -2284 6384 -2276
rect 6338 -2296 6384 -2284
rect 6456 -2284 6462 -2276
rect 6496 -2284 6502 -2276
rect 6456 -2296 6502 -2284
rect 6574 -2284 6580 -2276
rect 6614 -2284 6620 -2276
rect 6574 -2296 6620 -2284
rect 6692 -2284 6698 -2276
rect 6732 -2284 6738 -2276
rect 6692 -2296 6738 -2284
rect 6810 -2284 6816 -2276
rect 6850 -2284 6856 -2276
rect 6810 -2296 6856 -2284
rect 6928 -2284 6934 -2276
rect 6968 -2284 6974 -2276
rect 6928 -2296 6974 -2284
rect 7046 -2284 7052 -2276
rect 7086 -2284 7092 -2276
rect 7046 -2296 7092 -2284
rect 7164 -2284 7170 -2276
rect 7204 -2284 7210 -2276
rect 7164 -2296 7210 -2284
rect 7282 -2284 7288 -2276
rect 7322 -2284 7328 -2276
rect 7282 -2296 7328 -2284
rect 7400 -2284 7406 -2276
rect 7440 -2284 7446 -2276
rect 7400 -2296 7446 -2284
rect 7518 -2284 7524 -2276
rect 7558 -2284 7564 -2276
rect 7518 -2296 7564 -2284
rect 7636 -2284 7642 -2276
rect 7676 -2284 7682 -2276
rect 7636 -2296 7682 -2284
rect 7754 -2284 7760 -2276
rect 7794 -2284 7800 -2276
rect 7754 -2296 7800 -2284
rect 7872 -2284 7878 -2276
rect 7912 -2284 7918 -2276
rect 7872 -2296 7918 -2284
rect 7990 -2284 7996 -2276
rect 8030 -2284 8036 -2276
rect 7990 -2296 8036 -2284
rect 8108 -2284 8114 -2276
rect 8148 -2284 8154 -2276
rect 8108 -2296 8154 -2284
rect 8226 -2284 8232 -2276
rect 8266 -2284 8272 -2276
rect 8226 -2296 8272 -2284
rect 8344 -2284 8350 -2276
rect 8384 -2284 8390 -2276
rect 8344 -2296 8390 -2284
rect 8462 -2284 8468 -2276
rect 8502 -2284 8508 -2276
rect 8462 -2296 8508 -2284
rect 8580 -2284 8586 -2276
rect 8620 -2284 8626 -2276
rect 8580 -2296 8626 -2284
rect 8698 -2284 8704 -2276
rect 8738 -2284 8744 -2276
rect 8698 -2296 8744 -2284
rect 8816 -2284 8822 -2276
rect 8856 -2284 8862 -2276
rect 8816 -2296 8862 -2284
rect 8934 -2284 8940 -2276
rect 8974 -2284 8980 -2276
rect 8934 -2296 8980 -2284
rect 9052 -2284 9058 -2276
rect 9092 -2284 9098 -2276
rect 9052 -2296 9098 -2284
rect 9170 -2284 9176 -2276
rect 9210 -2284 9216 -2276
rect 9170 -2296 9216 -2284
rect 9288 -2284 9294 -2276
rect 9328 -2284 9334 -2276
rect 9288 -2296 9334 -2284
rect 9406 -2284 9412 -2276
rect 9446 -2284 9452 -2276
rect 9406 -2296 9452 -2284
rect 9524 -2284 9530 -2276
rect 9564 -2284 9570 -2276
rect 9524 -2296 9570 -2284
rect 9642 -2284 9648 -2276
rect 9682 -2284 9688 -2276
rect 9642 -2296 9688 -2284
rect 9760 -2284 9766 -2276
rect 9800 -2284 9806 -2276
rect 9760 -2296 9806 -2284
rect 9878 -2284 9884 -2276
rect 9918 -2284 9924 -2276
rect 9878 -2296 9924 -2284
rect 9996 -2284 10002 -2276
rect 10036 -2284 10042 -2276
rect 9996 -2296 10042 -2284
rect 10114 -2284 10120 -2276
rect 10154 -2284 10160 -2276
rect 10114 -2296 10160 -2284
rect 10232 -2284 10238 -2276
rect 10272 -2284 10278 -2276
rect 10232 -2296 10278 -2284
rect 10350 -2284 10356 -2276
rect 10390 -2284 10396 -2276
rect 10350 -2296 10396 -2284
rect 10468 -2284 10474 -2276
rect 10508 -2284 10514 -2276
rect 10468 -2296 10514 -2284
rect 10586 -2284 10592 -2276
rect 10626 -2284 10632 -2276
rect 10586 -2296 10632 -2284
rect 10704 -2284 10710 -2276
rect 10744 -2284 10750 -2276
rect 10704 -2296 10750 -2284
rect 4746 -2445 4801 -2425
rect 4853 -2445 5037 -2425
rect 5089 -2445 5273 -2425
rect 5325 -2445 5509 -2425
rect 5561 -2445 5745 -2425
rect 5797 -2445 5981 -2425
rect 6033 -2445 6217 -2425
rect 6269 -2445 6453 -2425
rect 6505 -2445 6689 -2425
rect 6741 -2445 6925 -2425
rect 6977 -2445 7161 -2425
rect 7213 -2445 7397 -2425
rect 7449 -2445 7633 -2425
rect 7685 -2445 7869 -2425
rect 7921 -2445 8105 -2425
rect 8157 -2445 8341 -2425
rect 8393 -2445 8577 -2425
rect 8629 -2445 8813 -2425
rect 8865 -2445 9049 -2425
rect 9101 -2445 9285 -2425
rect 9337 -2445 9521 -2425
rect 9573 -2445 9757 -2425
rect 9809 -2445 9993 -2425
rect 10045 -2445 10229 -2425
rect 10281 -2445 10465 -2425
rect 10517 -2445 10701 -2425
rect 10753 -2445 10794 -2425
rect 4746 -2479 4776 -2445
rect 4882 -2479 4920 -2445
rect 4954 -2479 4992 -2445
rect 5026 -2479 5037 -2445
rect 5098 -2479 5136 -2445
rect 5170 -2479 5208 -2445
rect 5242 -2479 5273 -2445
rect 5325 -2479 5352 -2445
rect 5386 -2479 5424 -2445
rect 5458 -2479 5496 -2445
rect 5561 -2479 5568 -2445
rect 5602 -2479 5640 -2445
rect 5674 -2479 5712 -2445
rect 5818 -2479 5856 -2445
rect 5890 -2479 5928 -2445
rect 5962 -2479 5981 -2445
rect 6034 -2479 6072 -2445
rect 6106 -2479 6144 -2445
rect 6178 -2479 6216 -2445
rect 6269 -2479 6288 -2445
rect 6322 -2479 6360 -2445
rect 6394 -2479 6432 -2445
rect 6538 -2479 6576 -2445
rect 6610 -2479 6648 -2445
rect 6682 -2479 6689 -2445
rect 6754 -2479 6792 -2445
rect 6826 -2479 6864 -2445
rect 6898 -2479 6925 -2445
rect 6977 -2479 7008 -2445
rect 7042 -2479 7080 -2445
rect 7114 -2479 7152 -2445
rect 7213 -2479 7224 -2445
rect 7258 -2479 7296 -2445
rect 7330 -2479 7368 -2445
rect 7474 -2479 7512 -2445
rect 7546 -2479 7584 -2445
rect 7618 -2479 7633 -2445
rect 7690 -2479 7728 -2445
rect 7762 -2479 7800 -2445
rect 7834 -2479 7869 -2445
rect 7921 -2479 7944 -2445
rect 7978 -2479 8016 -2445
rect 8050 -2479 8088 -2445
rect 8157 -2479 8160 -2445
rect 8194 -2479 8232 -2445
rect 8266 -2479 8304 -2445
rect 8338 -2479 8341 -2445
rect 8410 -2479 8448 -2445
rect 8482 -2479 8520 -2445
rect 8554 -2479 8577 -2445
rect 8629 -2479 8664 -2445
rect 8698 -2479 8736 -2445
rect 8770 -2479 8808 -2445
rect 8865 -2479 8880 -2445
rect 8914 -2479 8952 -2445
rect 8986 -2479 9024 -2445
rect 9130 -2479 9168 -2445
rect 9202 -2479 9240 -2445
rect 9274 -2479 9285 -2445
rect 9346 -2479 9384 -2445
rect 9418 -2479 9456 -2445
rect 9490 -2479 9521 -2445
rect 9573 -2479 9600 -2445
rect 9634 -2479 9672 -2445
rect 9706 -2479 9744 -2445
rect 9809 -2479 9816 -2445
rect 9850 -2479 9888 -2445
rect 9922 -2479 9960 -2445
rect 10066 -2479 10104 -2445
rect 10138 -2479 10176 -2445
rect 10210 -2479 10229 -2445
rect 10282 -2479 10320 -2445
rect 10354 -2479 10392 -2445
rect 10426 -2479 10464 -2445
rect 10517 -2479 10536 -2445
rect 10570 -2479 10608 -2445
rect 10642 -2479 10680 -2445
rect 10786 -2479 10794 -2445
rect 4746 -2533 4801 -2479
rect 4853 -2533 5037 -2479
rect 5089 -2533 5273 -2479
rect 5325 -2533 5509 -2479
rect 5561 -2533 5745 -2479
rect 5797 -2533 5981 -2479
rect 6033 -2533 6217 -2479
rect 6269 -2533 6453 -2479
rect 6505 -2533 6689 -2479
rect 6741 -2533 6925 -2479
rect 6977 -2533 7161 -2479
rect 7213 -2533 7397 -2479
rect 7449 -2533 7633 -2479
rect 7685 -2533 7869 -2479
rect 7921 -2533 8105 -2479
rect 8157 -2533 8341 -2479
rect 8393 -2533 8577 -2479
rect 8629 -2533 8813 -2479
rect 8865 -2533 9049 -2479
rect 9101 -2533 9285 -2479
rect 9337 -2533 9521 -2479
rect 9573 -2533 9757 -2479
rect 9809 -2533 9993 -2479
rect 10045 -2533 10229 -2479
rect 10281 -2533 10465 -2479
rect 10517 -2533 10701 -2479
rect 10753 -2533 10794 -2479
rect 4746 -2567 4776 -2533
rect 4882 -2567 4920 -2533
rect 4954 -2567 4992 -2533
rect 5026 -2567 5037 -2533
rect 5098 -2567 5136 -2533
rect 5170 -2567 5208 -2533
rect 5242 -2567 5273 -2533
rect 5325 -2567 5352 -2533
rect 5386 -2567 5424 -2533
rect 5458 -2567 5496 -2533
rect 5561 -2567 5568 -2533
rect 5602 -2567 5640 -2533
rect 5674 -2567 5712 -2533
rect 5818 -2567 5856 -2533
rect 5890 -2567 5928 -2533
rect 5962 -2567 5981 -2533
rect 6034 -2567 6072 -2533
rect 6106 -2567 6144 -2533
rect 6178 -2567 6216 -2533
rect 6269 -2567 6288 -2533
rect 6322 -2567 6360 -2533
rect 6394 -2567 6432 -2533
rect 6538 -2567 6576 -2533
rect 6610 -2567 6648 -2533
rect 6682 -2567 6689 -2533
rect 6754 -2567 6792 -2533
rect 6826 -2567 6864 -2533
rect 6898 -2567 6925 -2533
rect 6977 -2567 7008 -2533
rect 7042 -2567 7080 -2533
rect 7114 -2567 7152 -2533
rect 7213 -2567 7224 -2533
rect 7258 -2567 7296 -2533
rect 7330 -2567 7368 -2533
rect 7474 -2567 7512 -2533
rect 7546 -2567 7584 -2533
rect 7618 -2567 7633 -2533
rect 7690 -2567 7728 -2533
rect 7762 -2567 7800 -2533
rect 7834 -2567 7869 -2533
rect 7921 -2567 7944 -2533
rect 7978 -2567 8016 -2533
rect 8050 -2567 8088 -2533
rect 8157 -2567 8160 -2533
rect 8194 -2567 8232 -2533
rect 8266 -2567 8304 -2533
rect 8338 -2567 8341 -2533
rect 8410 -2567 8448 -2533
rect 8482 -2567 8520 -2533
rect 8554 -2567 8577 -2533
rect 8629 -2567 8664 -2533
rect 8698 -2567 8736 -2533
rect 8770 -2567 8808 -2533
rect 8865 -2567 8880 -2533
rect 8914 -2567 8952 -2533
rect 8986 -2567 9024 -2533
rect 9130 -2567 9168 -2533
rect 9202 -2567 9240 -2533
rect 9274 -2567 9285 -2533
rect 9346 -2567 9384 -2533
rect 9418 -2567 9456 -2533
rect 9490 -2567 9521 -2533
rect 9573 -2567 9600 -2533
rect 9634 -2567 9672 -2533
rect 9706 -2567 9744 -2533
rect 9809 -2567 9816 -2533
rect 9850 -2567 9888 -2533
rect 9922 -2567 9960 -2533
rect 10066 -2567 10104 -2533
rect 10138 -2567 10176 -2533
rect 10210 -2567 10229 -2533
rect 10282 -2567 10320 -2533
rect 10354 -2567 10392 -2533
rect 10426 -2567 10464 -2533
rect 10517 -2567 10536 -2533
rect 10570 -2567 10608 -2533
rect 10642 -2567 10680 -2533
rect 10786 -2567 10794 -2533
rect 4746 -2621 4801 -2567
rect 4853 -2621 5037 -2567
rect 5089 -2621 5273 -2567
rect 5325 -2621 5509 -2567
rect 5561 -2621 5745 -2567
rect 5797 -2621 5981 -2567
rect 6033 -2621 6217 -2567
rect 6269 -2621 6453 -2567
rect 6505 -2621 6689 -2567
rect 6741 -2621 6925 -2567
rect 6977 -2621 7161 -2567
rect 7213 -2621 7397 -2567
rect 7449 -2621 7633 -2567
rect 7685 -2621 7869 -2567
rect 7921 -2621 8105 -2567
rect 8157 -2621 8341 -2567
rect 8393 -2621 8577 -2567
rect 8629 -2621 8813 -2567
rect 8865 -2621 9049 -2567
rect 9101 -2621 9285 -2567
rect 9337 -2621 9521 -2567
rect 9573 -2621 9757 -2567
rect 9809 -2621 9993 -2567
rect 10045 -2621 10229 -2567
rect 10281 -2621 10465 -2567
rect 10517 -2621 10701 -2567
rect 10753 -2621 10794 -2567
rect 4746 -2655 4776 -2621
rect 4882 -2655 4920 -2621
rect 4954 -2655 4992 -2621
rect 5026 -2655 5037 -2621
rect 5098 -2655 5136 -2621
rect 5170 -2655 5208 -2621
rect 5242 -2655 5273 -2621
rect 5325 -2655 5352 -2621
rect 5386 -2655 5424 -2621
rect 5458 -2655 5496 -2621
rect 5561 -2655 5568 -2621
rect 5602 -2655 5640 -2621
rect 5674 -2655 5712 -2621
rect 5818 -2655 5856 -2621
rect 5890 -2655 5928 -2621
rect 5962 -2655 5981 -2621
rect 6034 -2655 6072 -2621
rect 6106 -2655 6144 -2621
rect 6178 -2655 6216 -2621
rect 6269 -2655 6288 -2621
rect 6322 -2655 6360 -2621
rect 6394 -2655 6432 -2621
rect 6538 -2655 6576 -2621
rect 6610 -2655 6648 -2621
rect 6682 -2655 6689 -2621
rect 6754 -2655 6792 -2621
rect 6826 -2655 6864 -2621
rect 6898 -2655 6925 -2621
rect 6977 -2655 7008 -2621
rect 7042 -2655 7080 -2621
rect 7114 -2655 7152 -2621
rect 7213 -2655 7224 -2621
rect 7258 -2655 7296 -2621
rect 7330 -2655 7368 -2621
rect 7474 -2655 7512 -2621
rect 7546 -2655 7584 -2621
rect 7618 -2655 7633 -2621
rect 7690 -2655 7728 -2621
rect 7762 -2655 7800 -2621
rect 7834 -2655 7869 -2621
rect 7921 -2655 7944 -2621
rect 7978 -2655 8016 -2621
rect 8050 -2655 8088 -2621
rect 8157 -2655 8160 -2621
rect 8194 -2655 8232 -2621
rect 8266 -2655 8304 -2621
rect 8338 -2655 8341 -2621
rect 8410 -2655 8448 -2621
rect 8482 -2655 8520 -2621
rect 8554 -2655 8577 -2621
rect 8629 -2655 8664 -2621
rect 8698 -2655 8736 -2621
rect 8770 -2655 8808 -2621
rect 8865 -2655 8880 -2621
rect 8914 -2655 8952 -2621
rect 8986 -2655 9024 -2621
rect 9130 -2655 9168 -2621
rect 9202 -2655 9240 -2621
rect 9274 -2655 9285 -2621
rect 9346 -2655 9384 -2621
rect 9418 -2655 9456 -2621
rect 9490 -2655 9521 -2621
rect 9573 -2655 9600 -2621
rect 9634 -2655 9672 -2621
rect 9706 -2655 9744 -2621
rect 9809 -2655 9816 -2621
rect 9850 -2655 9888 -2621
rect 9922 -2655 9960 -2621
rect 10066 -2655 10104 -2621
rect 10138 -2655 10176 -2621
rect 10210 -2655 10229 -2621
rect 10282 -2655 10320 -2621
rect 10354 -2655 10392 -2621
rect 10426 -2655 10464 -2621
rect 10517 -2655 10536 -2621
rect 10570 -2655 10608 -2621
rect 10642 -2655 10680 -2621
rect 10786 -2655 10794 -2621
rect 4746 -2675 4801 -2655
rect 4853 -2675 5037 -2655
rect 5089 -2675 5273 -2655
rect 5325 -2675 5509 -2655
rect 5561 -2675 5745 -2655
rect 5797 -2675 5981 -2655
rect 6033 -2675 6217 -2655
rect 6269 -2675 6453 -2655
rect 6505 -2675 6689 -2655
rect 6741 -2675 6925 -2655
rect 6977 -2675 7161 -2655
rect 7213 -2675 7397 -2655
rect 7449 -2675 7633 -2655
rect 7685 -2675 7869 -2655
rect 7921 -2675 8105 -2655
rect 8157 -2675 8341 -2655
rect 8393 -2675 8577 -2655
rect 8629 -2675 8813 -2655
rect 8865 -2675 9049 -2655
rect 9101 -2675 9285 -2655
rect 9337 -2675 9521 -2655
rect 9573 -2675 9757 -2655
rect 9809 -2675 9993 -2655
rect 10045 -2675 10229 -2655
rect 10281 -2675 10465 -2655
rect 10517 -2675 10701 -2655
rect 10753 -2675 10794 -2655
rect 4804 -2922 4850 -2910
rect 4804 -2930 4810 -2922
rect 4844 -2930 4850 -2922
rect 4922 -2922 4968 -2910
rect 4922 -2930 4928 -2922
rect 4962 -2930 4968 -2922
rect 5040 -2922 5086 -2910
rect 5040 -2930 5046 -2922
rect 5080 -2930 5086 -2922
rect 5158 -2922 5204 -2910
rect 5158 -2930 5164 -2922
rect 5198 -2930 5204 -2922
rect 5276 -2922 5322 -2910
rect 5276 -2930 5282 -2922
rect 5316 -2930 5322 -2922
rect 5394 -2922 5440 -2910
rect 5394 -2930 5400 -2922
rect 5434 -2930 5440 -2922
rect 5512 -2922 5558 -2910
rect 5512 -2930 5518 -2922
rect 5552 -2930 5558 -2922
rect 5630 -2922 5676 -2910
rect 5630 -2930 5636 -2922
rect 5670 -2930 5676 -2922
rect 5748 -2922 5794 -2910
rect 5748 -2930 5754 -2922
rect 5788 -2930 5794 -2922
rect 5866 -2922 5912 -2910
rect 5866 -2930 5872 -2922
rect 5906 -2930 5912 -2922
rect 5984 -2922 6030 -2910
rect 5984 -2930 5990 -2922
rect 6024 -2930 6030 -2922
rect 6102 -2922 6148 -2910
rect 6102 -2930 6108 -2922
rect 6142 -2930 6148 -2922
rect 6220 -2922 6266 -2910
rect 6220 -2930 6226 -2922
rect 6260 -2930 6266 -2922
rect 6338 -2922 6384 -2910
rect 6338 -2930 6344 -2922
rect 6378 -2930 6384 -2922
rect 6456 -2922 6502 -2910
rect 6456 -2930 6462 -2922
rect 6496 -2930 6502 -2922
rect 6574 -2922 6620 -2910
rect 6574 -2930 6580 -2922
rect 6614 -2930 6620 -2922
rect 6692 -2922 6738 -2910
rect 6692 -2930 6698 -2922
rect 6732 -2930 6738 -2922
rect 6810 -2922 6856 -2910
rect 6810 -2930 6816 -2922
rect 6850 -2930 6856 -2922
rect 6928 -2922 6974 -2910
rect 6928 -2930 6934 -2922
rect 6968 -2930 6974 -2922
rect 7046 -2922 7092 -2910
rect 7046 -2930 7052 -2922
rect 7086 -2930 7092 -2922
rect 7164 -2922 7210 -2910
rect 7164 -2930 7170 -2922
rect 7204 -2930 7210 -2922
rect 7282 -2922 7328 -2910
rect 7282 -2930 7288 -2922
rect 7322 -2930 7328 -2922
rect 7400 -2922 7446 -2910
rect 7400 -2930 7406 -2922
rect 7440 -2930 7446 -2922
rect 7518 -2922 7564 -2910
rect 7518 -2930 7524 -2922
rect 7558 -2930 7564 -2922
rect 7636 -2922 7682 -2910
rect 7636 -2930 7642 -2922
rect 7676 -2930 7682 -2922
rect 7754 -2922 7800 -2910
rect 7754 -2930 7760 -2922
rect 7794 -2930 7800 -2922
rect 7872 -2922 7918 -2910
rect 7872 -2930 7878 -2922
rect 7912 -2930 7918 -2922
rect 7990 -2922 8036 -2910
rect 7990 -2930 7996 -2922
rect 8030 -2930 8036 -2922
rect 8108 -2922 8154 -2910
rect 8108 -2930 8114 -2922
rect 8148 -2930 8154 -2922
rect 8226 -2922 8272 -2910
rect 8226 -2930 8232 -2922
rect 8266 -2930 8272 -2922
rect 8344 -2922 8390 -2910
rect 8344 -2930 8350 -2922
rect 8384 -2930 8390 -2922
rect 8462 -2922 8508 -2910
rect 8462 -2930 8468 -2922
rect 8502 -2930 8508 -2922
rect 8580 -2922 8626 -2910
rect 8580 -2930 8586 -2922
rect 8620 -2930 8626 -2922
rect 8698 -2922 8744 -2910
rect 8698 -2930 8704 -2922
rect 8738 -2930 8744 -2922
rect 8816 -2922 8862 -2910
rect 8816 -2930 8822 -2922
rect 8856 -2930 8862 -2922
rect 8934 -2922 8980 -2910
rect 8934 -2930 8940 -2922
rect 8974 -2930 8980 -2922
rect 9052 -2922 9098 -2910
rect 9052 -2930 9058 -2922
rect 9092 -2930 9098 -2922
rect 9170 -2922 9216 -2910
rect 9170 -2930 9176 -2922
rect 9210 -2930 9216 -2922
rect 9288 -2922 9334 -2910
rect 9288 -2930 9294 -2922
rect 9328 -2930 9334 -2922
rect 9406 -2922 9452 -2910
rect 9406 -2930 9412 -2922
rect 9446 -2930 9452 -2922
rect 9524 -2922 9570 -2910
rect 9524 -2930 9530 -2922
rect 9564 -2930 9570 -2922
rect 9642 -2922 9688 -2910
rect 9642 -2930 9648 -2922
rect 9682 -2930 9688 -2922
rect 9760 -2922 9806 -2910
rect 9760 -2930 9766 -2922
rect 9800 -2930 9806 -2922
rect 9878 -2922 9924 -2910
rect 9878 -2930 9884 -2922
rect 9918 -2930 9924 -2922
rect 9996 -2922 10042 -2910
rect 9996 -2930 10002 -2922
rect 10036 -2930 10042 -2922
rect 10114 -2922 10160 -2910
rect 10114 -2930 10120 -2922
rect 10154 -2930 10160 -2922
rect 10232 -2922 10278 -2910
rect 10232 -2930 10238 -2922
rect 10272 -2930 10278 -2922
rect 10350 -2922 10396 -2910
rect 10350 -2930 10356 -2922
rect 10390 -2930 10396 -2922
rect 10468 -2922 10514 -2910
rect 10468 -2930 10474 -2922
rect 10508 -2930 10514 -2922
rect 10586 -2922 10632 -2910
rect 10586 -2930 10592 -2922
rect 10626 -2930 10632 -2922
rect 10704 -2922 10750 -2910
rect 10704 -2930 10710 -2922
rect 10744 -2930 10750 -2922
rect 4791 -3490 4801 -2930
rect 4853 -3490 4863 -2930
rect 4911 -3490 4921 -2930
rect 4973 -3490 4983 -2930
rect 5027 -3490 5037 -2930
rect 5089 -3490 5099 -2930
rect 5147 -3490 5157 -2930
rect 5209 -3490 5219 -2930
rect 5263 -3490 5273 -2930
rect 5325 -3490 5335 -2930
rect 5383 -3490 5393 -2930
rect 5445 -3490 5455 -2930
rect 5499 -3490 5509 -2930
rect 5561 -3490 5571 -2930
rect 5619 -3490 5629 -2930
rect 5681 -3490 5691 -2930
rect 5735 -3490 5745 -2930
rect 5797 -3490 5807 -2930
rect 5855 -3490 5865 -2930
rect 5917 -3490 5927 -2930
rect 5971 -3490 5981 -2930
rect 6033 -3490 6043 -2930
rect 6091 -3490 6101 -2930
rect 6153 -3490 6163 -2930
rect 6207 -3490 6217 -2930
rect 6269 -3490 6279 -2930
rect 6327 -3490 6337 -2930
rect 6389 -3490 6399 -2930
rect 6443 -3490 6453 -2930
rect 6505 -3490 6515 -2930
rect 6563 -3490 6573 -2930
rect 6625 -3490 6635 -2930
rect 6679 -3490 6689 -2930
rect 6741 -3490 6751 -2930
rect 6799 -3490 6809 -2930
rect 6861 -3490 6871 -2930
rect 6915 -3490 6925 -2930
rect 6977 -3490 6987 -2930
rect 7035 -3490 7045 -2930
rect 7097 -3490 7107 -2930
rect 7151 -3490 7161 -2930
rect 7213 -3490 7223 -2930
rect 7271 -3490 7281 -2930
rect 7333 -3490 7343 -2930
rect 7387 -3490 7397 -2930
rect 7449 -3490 7459 -2930
rect 7507 -3490 7517 -2930
rect 7569 -3490 7579 -2930
rect 7623 -3490 7633 -2930
rect 7685 -3490 7695 -2930
rect 7743 -3490 7753 -2930
rect 7805 -3490 7815 -2930
rect 7859 -3490 7869 -2930
rect 7921 -3490 7931 -2930
rect 7979 -3490 7989 -2930
rect 8041 -3490 8051 -2930
rect 8095 -3490 8105 -2930
rect 8157 -3490 8167 -2930
rect 8215 -3490 8225 -2930
rect 8277 -3490 8287 -2930
rect 8331 -3490 8341 -2930
rect 8393 -3490 8403 -2930
rect 8451 -3490 8461 -2930
rect 8513 -3490 8523 -2930
rect 8567 -3490 8577 -2930
rect 8629 -3490 8639 -2930
rect 8687 -3490 8697 -2930
rect 8749 -3490 8759 -2930
rect 8803 -3490 8813 -2930
rect 8865 -3490 8875 -2930
rect 8923 -3490 8933 -2930
rect 8985 -3490 8995 -2930
rect 9039 -3490 9049 -2930
rect 9101 -3490 9111 -2930
rect 9159 -3490 9169 -2930
rect 9221 -3490 9231 -2930
rect 9275 -3490 9285 -2930
rect 9337 -3490 9347 -2930
rect 9395 -3490 9405 -2930
rect 9457 -3490 9467 -2930
rect 9511 -3490 9521 -2930
rect 9573 -3490 9583 -2930
rect 9631 -3490 9641 -2930
rect 9693 -3490 9703 -2930
rect 9747 -3490 9757 -2930
rect 9809 -3490 9819 -2930
rect 9867 -3490 9877 -2930
rect 9929 -3490 9939 -2930
rect 9983 -3490 9993 -2930
rect 10045 -3490 10055 -2930
rect 10103 -3490 10113 -2930
rect 10165 -3490 10175 -2930
rect 10219 -3490 10229 -2930
rect 10281 -3490 10291 -2930
rect 10339 -3490 10349 -2930
rect 10401 -3490 10411 -2930
rect 10455 -3490 10465 -2930
rect 10517 -3490 10527 -2930
rect 10575 -3490 10585 -2930
rect 10637 -3490 10647 -2930
rect 10691 -3490 10701 -2930
rect 10753 -3490 10763 -2930
rect 4804 -3498 4810 -3490
rect 4844 -3498 4850 -3490
rect 4804 -3510 4850 -3498
rect 4922 -3498 4928 -3490
rect 4962 -3498 4968 -3490
rect 4922 -3510 4968 -3498
rect 5040 -3498 5046 -3490
rect 5080 -3498 5086 -3490
rect 5040 -3510 5086 -3498
rect 5158 -3498 5164 -3490
rect 5198 -3498 5204 -3490
rect 5158 -3510 5204 -3498
rect 5276 -3498 5282 -3490
rect 5316 -3498 5322 -3490
rect 5276 -3510 5322 -3498
rect 5394 -3498 5400 -3490
rect 5434 -3498 5440 -3490
rect 5394 -3510 5440 -3498
rect 5512 -3498 5518 -3490
rect 5552 -3498 5558 -3490
rect 5512 -3510 5558 -3498
rect 5630 -3498 5636 -3490
rect 5670 -3498 5676 -3490
rect 5630 -3510 5676 -3498
rect 5748 -3498 5754 -3490
rect 5788 -3498 5794 -3490
rect 5748 -3510 5794 -3498
rect 5866 -3498 5872 -3490
rect 5906 -3498 5912 -3490
rect 5866 -3510 5912 -3498
rect 5984 -3498 5990 -3490
rect 6024 -3498 6030 -3490
rect 5984 -3510 6030 -3498
rect 6102 -3498 6108 -3490
rect 6142 -3498 6148 -3490
rect 6102 -3510 6148 -3498
rect 6220 -3498 6226 -3490
rect 6260 -3498 6266 -3490
rect 6220 -3510 6266 -3498
rect 6338 -3498 6344 -3490
rect 6378 -3498 6384 -3490
rect 6338 -3510 6384 -3498
rect 6456 -3498 6462 -3490
rect 6496 -3498 6502 -3490
rect 6456 -3510 6502 -3498
rect 6574 -3498 6580 -3490
rect 6614 -3498 6620 -3490
rect 6574 -3510 6620 -3498
rect 6692 -3498 6698 -3490
rect 6732 -3498 6738 -3490
rect 6692 -3510 6738 -3498
rect 6810 -3498 6816 -3490
rect 6850 -3498 6856 -3490
rect 6810 -3510 6856 -3498
rect 6928 -3498 6934 -3490
rect 6968 -3498 6974 -3490
rect 6928 -3510 6974 -3498
rect 7046 -3498 7052 -3490
rect 7086 -3498 7092 -3490
rect 7046 -3510 7092 -3498
rect 7164 -3498 7170 -3490
rect 7204 -3498 7210 -3490
rect 7164 -3510 7210 -3498
rect 7282 -3498 7288 -3490
rect 7322 -3498 7328 -3490
rect 7282 -3510 7328 -3498
rect 7400 -3498 7406 -3490
rect 7440 -3498 7446 -3490
rect 7400 -3510 7446 -3498
rect 7518 -3498 7524 -3490
rect 7558 -3498 7564 -3490
rect 7518 -3510 7564 -3498
rect 7636 -3498 7642 -3490
rect 7676 -3498 7682 -3490
rect 7636 -3510 7682 -3498
rect 7754 -3498 7760 -3490
rect 7794 -3498 7800 -3490
rect 7754 -3510 7800 -3498
rect 7872 -3498 7878 -3490
rect 7912 -3498 7918 -3490
rect 7872 -3510 7918 -3498
rect 7990 -3498 7996 -3490
rect 8030 -3498 8036 -3490
rect 7990 -3510 8036 -3498
rect 8108 -3498 8114 -3490
rect 8148 -3498 8154 -3490
rect 8108 -3510 8154 -3498
rect 8226 -3498 8232 -3490
rect 8266 -3498 8272 -3490
rect 8226 -3510 8272 -3498
rect 8344 -3498 8350 -3490
rect 8384 -3498 8390 -3490
rect 8344 -3510 8390 -3498
rect 8462 -3498 8468 -3490
rect 8502 -3498 8508 -3490
rect 8462 -3510 8508 -3498
rect 8580 -3498 8586 -3490
rect 8620 -3498 8626 -3490
rect 8580 -3510 8626 -3498
rect 8698 -3498 8704 -3490
rect 8738 -3498 8744 -3490
rect 8698 -3510 8744 -3498
rect 8816 -3498 8822 -3490
rect 8856 -3498 8862 -3490
rect 8816 -3510 8862 -3498
rect 8934 -3498 8940 -3490
rect 8974 -3498 8980 -3490
rect 8934 -3510 8980 -3498
rect 9052 -3498 9058 -3490
rect 9092 -3498 9098 -3490
rect 9052 -3510 9098 -3498
rect 9170 -3498 9176 -3490
rect 9210 -3498 9216 -3490
rect 9170 -3510 9216 -3498
rect 9288 -3498 9294 -3490
rect 9328 -3498 9334 -3490
rect 9288 -3510 9334 -3498
rect 9406 -3498 9412 -3490
rect 9446 -3498 9452 -3490
rect 9406 -3510 9452 -3498
rect 9524 -3498 9530 -3490
rect 9564 -3498 9570 -3490
rect 9524 -3510 9570 -3498
rect 9642 -3498 9648 -3490
rect 9682 -3498 9688 -3490
rect 9642 -3510 9688 -3498
rect 9760 -3498 9766 -3490
rect 9800 -3498 9806 -3490
rect 9760 -3510 9806 -3498
rect 9878 -3498 9884 -3490
rect 9918 -3498 9924 -3490
rect 9878 -3510 9924 -3498
rect 9996 -3498 10002 -3490
rect 10036 -3498 10042 -3490
rect 9996 -3510 10042 -3498
rect 10114 -3498 10120 -3490
rect 10154 -3498 10160 -3490
rect 10114 -3510 10160 -3498
rect 10232 -3498 10238 -3490
rect 10272 -3498 10278 -3490
rect 10232 -3510 10278 -3498
rect 10350 -3498 10356 -3490
rect 10390 -3498 10396 -3490
rect 10350 -3510 10396 -3498
rect 10468 -3498 10474 -3490
rect 10508 -3498 10514 -3490
rect 10468 -3510 10514 -3498
rect 10586 -3498 10592 -3490
rect 10626 -3498 10632 -3490
rect 10586 -3510 10632 -3498
rect 10704 -3498 10710 -3490
rect 10744 -3498 10750 -3490
rect 10704 -3510 10750 -3498
rect 4847 -3705 4857 -3551
rect 4915 -3705 4925 -3551
rect 4965 -3705 4975 -3551
rect 5033 -3705 5043 -3551
rect 5083 -3705 5093 -3551
rect 5151 -3705 5161 -3551
rect 5201 -3705 5211 -3551
rect 5269 -3705 5279 -3551
rect 5319 -3705 5329 -3551
rect 5387 -3705 5397 -3551
rect 5437 -3705 5447 -3551
rect 5505 -3705 5515 -3551
rect 5555 -3705 5565 -3551
rect 5623 -3705 5633 -3551
rect 5673 -3705 5683 -3551
rect 5741 -3705 5751 -3551
rect 5791 -3705 5801 -3551
rect 5859 -3705 5869 -3551
rect 5909 -3705 5919 -3551
rect 5977 -3705 5987 -3551
rect 6027 -3705 6037 -3551
rect 6095 -3705 6105 -3551
rect 6145 -3705 6155 -3551
rect 6213 -3705 6223 -3551
rect 6263 -3705 6273 -3551
rect 6331 -3705 6341 -3551
rect 6381 -3705 6391 -3551
rect 6449 -3705 6459 -3551
rect 6499 -3705 6509 -3551
rect 6567 -3705 6577 -3551
rect 6617 -3705 6627 -3551
rect 6685 -3705 6695 -3551
rect 6735 -3705 6745 -3551
rect 6803 -3705 6813 -3551
rect 6853 -3705 6863 -3551
rect 6921 -3705 6931 -3551
rect 6971 -3705 6981 -3551
rect 7039 -3705 7049 -3551
rect 7089 -3705 7099 -3551
rect 7157 -3705 7167 -3551
rect 7207 -3705 7217 -3551
rect 7275 -3705 7285 -3551
rect 7325 -3705 7335 -3551
rect 7393 -3705 7403 -3551
rect 7443 -3705 7453 -3551
rect 7511 -3705 7521 -3551
rect 7561 -3705 7571 -3551
rect 7629 -3705 7639 -3551
rect 7679 -3705 7689 -3551
rect 7747 -3705 7757 -3551
rect 7797 -3705 7807 -3551
rect 7865 -3705 7875 -3551
rect 7915 -3705 7925 -3551
rect 7983 -3705 7993 -3551
rect 8033 -3705 8043 -3551
rect 8101 -3705 8111 -3551
rect 8151 -3705 8161 -3551
rect 8219 -3705 8229 -3551
rect 8269 -3705 8279 -3551
rect 8337 -3705 8347 -3551
rect 8387 -3705 8397 -3551
rect 8455 -3705 8465 -3551
rect 8505 -3705 8515 -3551
rect 8573 -3705 8583 -3551
rect 8623 -3705 8633 -3551
rect 8691 -3705 8701 -3551
rect 8741 -3705 8751 -3551
rect 8809 -3705 8819 -3551
rect 8859 -3705 8869 -3551
rect 8927 -3705 8937 -3551
rect 8977 -3705 8987 -3551
rect 9045 -3705 9055 -3551
rect 9095 -3705 9105 -3551
rect 9163 -3705 9173 -3551
rect 9213 -3705 9223 -3551
rect 9281 -3705 9291 -3551
rect 9331 -3705 9341 -3551
rect 9399 -3705 9409 -3551
rect 9449 -3705 9459 -3551
rect 9517 -3705 9527 -3551
rect 9567 -3705 9577 -3551
rect 9635 -3705 9645 -3551
rect 9685 -3705 9695 -3551
rect 9753 -3705 9763 -3551
rect 9803 -3705 9813 -3551
rect 9871 -3705 9881 -3551
rect 9921 -3705 9931 -3551
rect 9989 -3705 9999 -3551
rect 10039 -3705 10049 -3551
rect 10107 -3705 10117 -3551
rect 10157 -3705 10167 -3551
rect 10225 -3705 10235 -3551
rect 10275 -3705 10285 -3551
rect 10343 -3705 10353 -3551
rect 10393 -3705 10403 -3551
rect 10461 -3705 10471 -3551
rect 10511 -3705 10521 -3551
rect 10579 -3705 10589 -3551
rect 10629 -3705 10639 -3551
rect 10697 -3705 10707 -3551
rect 4804 -3758 4850 -3746
rect 4804 -3766 4810 -3758
rect 4844 -3766 4850 -3758
rect 4922 -3758 4968 -3746
rect 4922 -3766 4928 -3758
rect 4962 -3766 4968 -3758
rect 5040 -3758 5086 -3746
rect 5040 -3766 5046 -3758
rect 5080 -3766 5086 -3758
rect 5158 -3758 5204 -3746
rect 5158 -3766 5164 -3758
rect 5198 -3766 5204 -3758
rect 5276 -3758 5322 -3746
rect 5276 -3766 5282 -3758
rect 5316 -3766 5322 -3758
rect 5394 -3758 5440 -3746
rect 5394 -3766 5400 -3758
rect 5434 -3766 5440 -3758
rect 5512 -3758 5558 -3746
rect 5512 -3766 5518 -3758
rect 5552 -3766 5558 -3758
rect 5630 -3758 5676 -3746
rect 5630 -3766 5636 -3758
rect 5670 -3766 5676 -3758
rect 5748 -3758 5794 -3746
rect 5748 -3766 5754 -3758
rect 5788 -3766 5794 -3758
rect 5866 -3758 5912 -3746
rect 5866 -3766 5872 -3758
rect 5906 -3766 5912 -3758
rect 5984 -3758 6030 -3746
rect 5984 -3766 5990 -3758
rect 6024 -3766 6030 -3758
rect 6102 -3758 6148 -3746
rect 6102 -3766 6108 -3758
rect 6142 -3766 6148 -3758
rect 6220 -3758 6266 -3746
rect 6220 -3766 6226 -3758
rect 6260 -3766 6266 -3758
rect 6338 -3758 6384 -3746
rect 6338 -3766 6344 -3758
rect 6378 -3766 6384 -3758
rect 6456 -3758 6502 -3746
rect 6456 -3766 6462 -3758
rect 6496 -3766 6502 -3758
rect 6574 -3758 6620 -3746
rect 6574 -3766 6580 -3758
rect 6614 -3766 6620 -3758
rect 6692 -3758 6738 -3746
rect 6692 -3766 6698 -3758
rect 6732 -3766 6738 -3758
rect 6810 -3758 6856 -3746
rect 6810 -3766 6816 -3758
rect 6850 -3766 6856 -3758
rect 6928 -3758 6974 -3746
rect 6928 -3766 6934 -3758
rect 6968 -3766 6974 -3758
rect 7046 -3758 7092 -3746
rect 7046 -3766 7052 -3758
rect 7086 -3766 7092 -3758
rect 7164 -3758 7210 -3746
rect 7164 -3766 7170 -3758
rect 7204 -3766 7210 -3758
rect 7282 -3758 7328 -3746
rect 7282 -3766 7288 -3758
rect 7322 -3766 7328 -3758
rect 7400 -3758 7446 -3746
rect 7400 -3766 7406 -3758
rect 7440 -3766 7446 -3758
rect 7518 -3758 7564 -3746
rect 7518 -3766 7524 -3758
rect 7558 -3766 7564 -3758
rect 7636 -3758 7682 -3746
rect 7636 -3766 7642 -3758
rect 7676 -3766 7682 -3758
rect 7754 -3758 7800 -3746
rect 7754 -3766 7760 -3758
rect 7794 -3766 7800 -3758
rect 7872 -3758 7918 -3746
rect 7872 -3766 7878 -3758
rect 7912 -3766 7918 -3758
rect 7990 -3758 8036 -3746
rect 7990 -3766 7996 -3758
rect 8030 -3766 8036 -3758
rect 8108 -3758 8154 -3746
rect 8108 -3766 8114 -3758
rect 8148 -3766 8154 -3758
rect 8226 -3758 8272 -3746
rect 8226 -3766 8232 -3758
rect 8266 -3766 8272 -3758
rect 8344 -3758 8390 -3746
rect 8344 -3766 8350 -3758
rect 8384 -3766 8390 -3758
rect 8462 -3758 8508 -3746
rect 8462 -3766 8468 -3758
rect 8502 -3766 8508 -3758
rect 8580 -3758 8626 -3746
rect 8580 -3766 8586 -3758
rect 8620 -3766 8626 -3758
rect 8698 -3758 8744 -3746
rect 8698 -3766 8704 -3758
rect 8738 -3766 8744 -3758
rect 8816 -3758 8862 -3746
rect 8816 -3766 8822 -3758
rect 8856 -3766 8862 -3758
rect 8934 -3758 8980 -3746
rect 8934 -3766 8940 -3758
rect 8974 -3766 8980 -3758
rect 9052 -3758 9098 -3746
rect 9052 -3766 9058 -3758
rect 9092 -3766 9098 -3758
rect 9170 -3758 9216 -3746
rect 9170 -3766 9176 -3758
rect 9210 -3766 9216 -3758
rect 9288 -3758 9334 -3746
rect 9288 -3766 9294 -3758
rect 9328 -3766 9334 -3758
rect 9406 -3758 9452 -3746
rect 9406 -3766 9412 -3758
rect 9446 -3766 9452 -3758
rect 9524 -3758 9570 -3746
rect 9524 -3766 9530 -3758
rect 9564 -3766 9570 -3758
rect 9642 -3758 9688 -3746
rect 9642 -3766 9648 -3758
rect 9682 -3766 9688 -3758
rect 9760 -3758 9806 -3746
rect 9760 -3766 9766 -3758
rect 9800 -3766 9806 -3758
rect 9878 -3758 9924 -3746
rect 9878 -3766 9884 -3758
rect 9918 -3766 9924 -3758
rect 9996 -3758 10042 -3746
rect 9996 -3766 10002 -3758
rect 10036 -3766 10042 -3758
rect 10114 -3758 10160 -3746
rect 10114 -3766 10120 -3758
rect 10154 -3766 10160 -3758
rect 10232 -3758 10278 -3746
rect 10232 -3766 10238 -3758
rect 10272 -3766 10278 -3758
rect 10350 -3758 10396 -3746
rect 10350 -3766 10356 -3758
rect 10390 -3766 10396 -3758
rect 10468 -3758 10514 -3746
rect 10468 -3766 10474 -3758
rect 10508 -3766 10514 -3758
rect 10586 -3758 10632 -3746
rect 10586 -3766 10592 -3758
rect 10626 -3766 10632 -3758
rect 10704 -3758 10750 -3746
rect 10704 -3766 10710 -3758
rect 10744 -3766 10750 -3758
rect 4791 -4326 4801 -3766
rect 4853 -4326 4863 -3766
rect 4911 -4326 4921 -3766
rect 4973 -4326 4983 -3766
rect 5027 -4326 5037 -3766
rect 5089 -4326 5099 -3766
rect 5147 -4326 5157 -3766
rect 5209 -4326 5219 -3766
rect 5263 -4326 5273 -3766
rect 5325 -4326 5335 -3766
rect 5383 -4326 5393 -3766
rect 5445 -4326 5455 -3766
rect 5499 -4326 5509 -3766
rect 5561 -4326 5571 -3766
rect 5619 -4326 5629 -3766
rect 5681 -4326 5691 -3766
rect 5735 -4326 5745 -3766
rect 5797 -4326 5807 -3766
rect 5855 -4326 5865 -3766
rect 5917 -4326 5927 -3766
rect 5971 -4326 5981 -3766
rect 6033 -4326 6043 -3766
rect 6091 -4326 6101 -3766
rect 6153 -4326 6163 -3766
rect 6207 -4326 6217 -3766
rect 6269 -4326 6279 -3766
rect 6327 -4326 6337 -3766
rect 6389 -4326 6399 -3766
rect 6443 -4326 6453 -3766
rect 6505 -4326 6515 -3766
rect 6563 -4326 6573 -3766
rect 6625 -4326 6635 -3766
rect 6679 -4326 6689 -3766
rect 6741 -4326 6751 -3766
rect 6799 -4326 6809 -3766
rect 6861 -4326 6871 -3766
rect 6915 -4326 6925 -3766
rect 6977 -4326 6987 -3766
rect 7035 -4326 7045 -3766
rect 7097 -4326 7107 -3766
rect 7151 -4326 7161 -3766
rect 7213 -4326 7223 -3766
rect 7271 -4326 7281 -3766
rect 7333 -4326 7343 -3766
rect 7387 -4326 7397 -3766
rect 7449 -4326 7459 -3766
rect 7507 -4326 7517 -3766
rect 7569 -4326 7579 -3766
rect 7623 -4326 7633 -3766
rect 7685 -4326 7695 -3766
rect 7743 -4326 7753 -3766
rect 7805 -4326 7815 -3766
rect 7859 -4326 7869 -3766
rect 7921 -4326 7931 -3766
rect 7979 -4326 7989 -3766
rect 8041 -4326 8051 -3766
rect 8095 -4326 8105 -3766
rect 8157 -4326 8167 -3766
rect 8215 -4326 8225 -3766
rect 8277 -4326 8287 -3766
rect 8331 -4326 8341 -3766
rect 8393 -4326 8403 -3766
rect 8451 -4326 8461 -3766
rect 8513 -4326 8523 -3766
rect 8567 -4326 8577 -3766
rect 8629 -4326 8639 -3766
rect 8687 -4326 8697 -3766
rect 8749 -4326 8759 -3766
rect 8803 -4326 8813 -3766
rect 8865 -4326 8875 -3766
rect 8923 -4326 8933 -3766
rect 8985 -4326 8995 -3766
rect 9039 -4326 9049 -3766
rect 9101 -4326 9111 -3766
rect 9159 -4326 9169 -3766
rect 9221 -4326 9231 -3766
rect 9275 -4326 9285 -3766
rect 9337 -4326 9347 -3766
rect 9395 -4326 9405 -3766
rect 9457 -4326 9467 -3766
rect 9511 -4326 9521 -3766
rect 9573 -4326 9583 -3766
rect 9631 -4326 9641 -3766
rect 9693 -4326 9703 -3766
rect 9747 -4326 9757 -3766
rect 9809 -4326 9819 -3766
rect 9867 -4326 9877 -3766
rect 9929 -4326 9939 -3766
rect 9983 -4326 9993 -3766
rect 10045 -4326 10055 -3766
rect 10103 -4326 10113 -3766
rect 10165 -4326 10175 -3766
rect 10219 -4326 10229 -3766
rect 10281 -4326 10291 -3766
rect 10339 -4326 10349 -3766
rect 10401 -4326 10411 -3766
rect 10455 -4326 10465 -3766
rect 10517 -4326 10527 -3766
rect 10575 -4326 10585 -3766
rect 10637 -4326 10647 -3766
rect 10691 -4326 10701 -3766
rect 10753 -4326 10763 -3766
rect 4804 -4334 4810 -4326
rect 4844 -4334 4850 -4326
rect 4804 -4346 4850 -4334
rect 4922 -4334 4928 -4326
rect 4962 -4334 4968 -4326
rect 4922 -4346 4968 -4334
rect 5040 -4334 5046 -4326
rect 5080 -4334 5086 -4326
rect 5040 -4346 5086 -4334
rect 5158 -4334 5164 -4326
rect 5198 -4334 5204 -4326
rect 5158 -4346 5204 -4334
rect 5276 -4334 5282 -4326
rect 5316 -4334 5322 -4326
rect 5276 -4346 5322 -4334
rect 5394 -4334 5400 -4326
rect 5434 -4334 5440 -4326
rect 5394 -4346 5440 -4334
rect 5512 -4334 5518 -4326
rect 5552 -4334 5558 -4326
rect 5512 -4346 5558 -4334
rect 5630 -4334 5636 -4326
rect 5670 -4334 5676 -4326
rect 5630 -4346 5676 -4334
rect 5748 -4334 5754 -4326
rect 5788 -4334 5794 -4326
rect 5748 -4346 5794 -4334
rect 5866 -4334 5872 -4326
rect 5906 -4334 5912 -4326
rect 5866 -4346 5912 -4334
rect 5984 -4334 5990 -4326
rect 6024 -4334 6030 -4326
rect 5984 -4346 6030 -4334
rect 6102 -4334 6108 -4326
rect 6142 -4334 6148 -4326
rect 6102 -4346 6148 -4334
rect 6220 -4334 6226 -4326
rect 6260 -4334 6266 -4326
rect 6220 -4346 6266 -4334
rect 6338 -4334 6344 -4326
rect 6378 -4334 6384 -4326
rect 6338 -4346 6384 -4334
rect 6456 -4334 6462 -4326
rect 6496 -4334 6502 -4326
rect 6456 -4346 6502 -4334
rect 6574 -4334 6580 -4326
rect 6614 -4334 6620 -4326
rect 6574 -4346 6620 -4334
rect 6692 -4334 6698 -4326
rect 6732 -4334 6738 -4326
rect 6692 -4346 6738 -4334
rect 6810 -4334 6816 -4326
rect 6850 -4334 6856 -4326
rect 6810 -4346 6856 -4334
rect 6928 -4334 6934 -4326
rect 6968 -4334 6974 -4326
rect 6928 -4346 6974 -4334
rect 7046 -4334 7052 -4326
rect 7086 -4334 7092 -4326
rect 7046 -4346 7092 -4334
rect 7164 -4334 7170 -4326
rect 7204 -4334 7210 -4326
rect 7164 -4346 7210 -4334
rect 7282 -4334 7288 -4326
rect 7322 -4334 7328 -4326
rect 7282 -4346 7328 -4334
rect 7400 -4334 7406 -4326
rect 7440 -4334 7446 -4326
rect 7400 -4346 7446 -4334
rect 7518 -4334 7524 -4326
rect 7558 -4334 7564 -4326
rect 7518 -4346 7564 -4334
rect 7636 -4334 7642 -4326
rect 7676 -4334 7682 -4326
rect 7636 -4346 7682 -4334
rect 7754 -4334 7760 -4326
rect 7794 -4334 7800 -4326
rect 7754 -4346 7800 -4334
rect 7872 -4334 7878 -4326
rect 7912 -4334 7918 -4326
rect 7872 -4346 7918 -4334
rect 7990 -4334 7996 -4326
rect 8030 -4334 8036 -4326
rect 7990 -4346 8036 -4334
rect 8108 -4334 8114 -4326
rect 8148 -4334 8154 -4326
rect 8108 -4346 8154 -4334
rect 8226 -4334 8232 -4326
rect 8266 -4334 8272 -4326
rect 8226 -4346 8272 -4334
rect 8344 -4334 8350 -4326
rect 8384 -4334 8390 -4326
rect 8344 -4346 8390 -4334
rect 8462 -4334 8468 -4326
rect 8502 -4334 8508 -4326
rect 8462 -4346 8508 -4334
rect 8580 -4334 8586 -4326
rect 8620 -4334 8626 -4326
rect 8580 -4346 8626 -4334
rect 8698 -4334 8704 -4326
rect 8738 -4334 8744 -4326
rect 8698 -4346 8744 -4334
rect 8816 -4334 8822 -4326
rect 8856 -4334 8862 -4326
rect 8816 -4346 8862 -4334
rect 8934 -4334 8940 -4326
rect 8974 -4334 8980 -4326
rect 8934 -4346 8980 -4334
rect 9052 -4334 9058 -4326
rect 9092 -4334 9098 -4326
rect 9052 -4346 9098 -4334
rect 9170 -4334 9176 -4326
rect 9210 -4334 9216 -4326
rect 9170 -4346 9216 -4334
rect 9288 -4334 9294 -4326
rect 9328 -4334 9334 -4326
rect 9288 -4346 9334 -4334
rect 9406 -4334 9412 -4326
rect 9446 -4334 9452 -4326
rect 9406 -4346 9452 -4334
rect 9524 -4334 9530 -4326
rect 9564 -4334 9570 -4326
rect 9524 -4346 9570 -4334
rect 9642 -4334 9648 -4326
rect 9682 -4334 9688 -4326
rect 9642 -4346 9688 -4334
rect 9760 -4334 9766 -4326
rect 9800 -4334 9806 -4326
rect 9760 -4346 9806 -4334
rect 9878 -4334 9884 -4326
rect 9918 -4334 9924 -4326
rect 9878 -4346 9924 -4334
rect 9996 -4334 10002 -4326
rect 10036 -4334 10042 -4326
rect 9996 -4346 10042 -4334
rect 10114 -4334 10120 -4326
rect 10154 -4334 10160 -4326
rect 10114 -4346 10160 -4334
rect 10232 -4334 10238 -4326
rect 10272 -4334 10278 -4326
rect 10232 -4346 10278 -4334
rect 10350 -4334 10356 -4326
rect 10390 -4334 10396 -4326
rect 10350 -4346 10396 -4334
rect 10468 -4334 10474 -4326
rect 10508 -4334 10514 -4326
rect 10468 -4346 10514 -4334
rect 10586 -4334 10592 -4326
rect 10626 -4334 10632 -4326
rect 10586 -4346 10632 -4334
rect 10704 -4334 10710 -4326
rect 10744 -4334 10750 -4326
rect 10704 -4346 10750 -4334
rect 4744 -4495 4801 -4475
rect 4853 -4495 5037 -4475
rect 5089 -4495 5273 -4475
rect 5325 -4495 5509 -4475
rect 5561 -4495 5745 -4475
rect 5797 -4495 5981 -4475
rect 6033 -4495 6217 -4475
rect 6269 -4495 6453 -4475
rect 6505 -4495 6689 -4475
rect 6741 -4495 6925 -4475
rect 6977 -4495 7161 -4475
rect 7213 -4495 7397 -4475
rect 7449 -4495 7633 -4475
rect 7685 -4495 7869 -4475
rect 7921 -4495 8105 -4475
rect 8157 -4495 8341 -4475
rect 8393 -4495 8577 -4475
rect 8629 -4495 8813 -4475
rect 8865 -4495 9049 -4475
rect 9101 -4495 9285 -4475
rect 9337 -4495 9521 -4475
rect 9573 -4495 9757 -4475
rect 9809 -4495 9993 -4475
rect 10045 -4495 10229 -4475
rect 10281 -4495 10465 -4475
rect 10517 -4495 10701 -4475
rect 10753 -4495 10808 -4475
rect 4744 -4529 4768 -4495
rect 4874 -4529 4912 -4495
rect 4946 -4529 4984 -4495
rect 5018 -4529 5037 -4495
rect 5090 -4529 5128 -4495
rect 5162 -4529 5200 -4495
rect 5234 -4529 5272 -4495
rect 5325 -4529 5344 -4495
rect 5378 -4529 5416 -4495
rect 5450 -4529 5488 -4495
rect 5594 -4529 5632 -4495
rect 5666 -4529 5704 -4495
rect 5738 -4529 5745 -4495
rect 5810 -4529 5848 -4495
rect 5882 -4529 5920 -4495
rect 5954 -4529 5981 -4495
rect 6033 -4529 6064 -4495
rect 6098 -4529 6136 -4495
rect 6170 -4529 6208 -4495
rect 6269 -4529 6280 -4495
rect 6314 -4529 6352 -4495
rect 6386 -4529 6424 -4495
rect 6530 -4529 6568 -4495
rect 6602 -4529 6640 -4495
rect 6674 -4529 6689 -4495
rect 6746 -4529 6784 -4495
rect 6818 -4529 6856 -4495
rect 6890 -4529 6925 -4495
rect 6977 -4529 7000 -4495
rect 7034 -4529 7072 -4495
rect 7106 -4529 7144 -4495
rect 7213 -4529 7216 -4495
rect 7250 -4529 7288 -4495
rect 7322 -4529 7360 -4495
rect 7394 -4529 7397 -4495
rect 7466 -4529 7504 -4495
rect 7538 -4529 7576 -4495
rect 7610 -4529 7633 -4495
rect 7685 -4529 7720 -4495
rect 7754 -4529 7792 -4495
rect 7826 -4529 7864 -4495
rect 7921 -4529 7936 -4495
rect 7970 -4529 8008 -4495
rect 8042 -4529 8080 -4495
rect 8186 -4529 8224 -4495
rect 8258 -4529 8296 -4495
rect 8330 -4529 8341 -4495
rect 8402 -4529 8440 -4495
rect 8474 -4529 8512 -4495
rect 8546 -4529 8577 -4495
rect 8629 -4529 8656 -4495
rect 8690 -4529 8728 -4495
rect 8762 -4529 8800 -4495
rect 8865 -4529 8872 -4495
rect 8906 -4529 8944 -4495
rect 8978 -4529 9016 -4495
rect 9122 -4529 9160 -4495
rect 9194 -4529 9232 -4495
rect 9266 -4529 9285 -4495
rect 9338 -4529 9376 -4495
rect 9410 -4529 9448 -4495
rect 9482 -4529 9520 -4495
rect 9573 -4529 9592 -4495
rect 9626 -4529 9664 -4495
rect 9698 -4529 9736 -4495
rect 9842 -4529 9880 -4495
rect 9914 -4529 9952 -4495
rect 9986 -4529 9993 -4495
rect 10058 -4529 10096 -4495
rect 10130 -4529 10168 -4495
rect 10202 -4529 10229 -4495
rect 10281 -4529 10312 -4495
rect 10346 -4529 10384 -4495
rect 10418 -4529 10456 -4495
rect 10517 -4529 10528 -4495
rect 10562 -4529 10600 -4495
rect 10634 -4529 10672 -4495
rect 10778 -4529 10808 -4495
rect 4744 -4583 4801 -4529
rect 4853 -4583 5037 -4529
rect 5089 -4583 5273 -4529
rect 5325 -4583 5509 -4529
rect 5561 -4583 5745 -4529
rect 5797 -4583 5981 -4529
rect 6033 -4583 6217 -4529
rect 6269 -4583 6453 -4529
rect 6505 -4583 6689 -4529
rect 6741 -4583 6925 -4529
rect 6977 -4583 7161 -4529
rect 7213 -4583 7397 -4529
rect 7449 -4583 7633 -4529
rect 7685 -4583 7869 -4529
rect 7921 -4583 8105 -4529
rect 8157 -4583 8341 -4529
rect 8393 -4583 8577 -4529
rect 8629 -4583 8813 -4529
rect 8865 -4583 9049 -4529
rect 9101 -4583 9285 -4529
rect 9337 -4583 9521 -4529
rect 9573 -4583 9757 -4529
rect 9809 -4583 9993 -4529
rect 10045 -4583 10229 -4529
rect 10281 -4583 10465 -4529
rect 10517 -4583 10701 -4529
rect 10753 -4583 10808 -4529
rect 4744 -4617 4768 -4583
rect 4874 -4617 4912 -4583
rect 4946 -4617 4984 -4583
rect 5018 -4617 5037 -4583
rect 5090 -4617 5128 -4583
rect 5162 -4617 5200 -4583
rect 5234 -4617 5272 -4583
rect 5325 -4617 5344 -4583
rect 5378 -4617 5416 -4583
rect 5450 -4617 5488 -4583
rect 5594 -4617 5632 -4583
rect 5666 -4617 5704 -4583
rect 5738 -4617 5745 -4583
rect 5810 -4617 5848 -4583
rect 5882 -4617 5920 -4583
rect 5954 -4617 5981 -4583
rect 6033 -4617 6064 -4583
rect 6098 -4617 6136 -4583
rect 6170 -4617 6208 -4583
rect 6269 -4617 6280 -4583
rect 6314 -4617 6352 -4583
rect 6386 -4617 6424 -4583
rect 6530 -4617 6568 -4583
rect 6602 -4617 6640 -4583
rect 6674 -4617 6689 -4583
rect 6746 -4617 6784 -4583
rect 6818 -4617 6856 -4583
rect 6890 -4617 6925 -4583
rect 6977 -4617 7000 -4583
rect 7034 -4617 7072 -4583
rect 7106 -4617 7144 -4583
rect 7213 -4617 7216 -4583
rect 7250 -4617 7288 -4583
rect 7322 -4617 7360 -4583
rect 7394 -4617 7397 -4583
rect 7466 -4617 7504 -4583
rect 7538 -4617 7576 -4583
rect 7610 -4617 7633 -4583
rect 7685 -4617 7720 -4583
rect 7754 -4617 7792 -4583
rect 7826 -4617 7864 -4583
rect 7921 -4617 7936 -4583
rect 7970 -4617 8008 -4583
rect 8042 -4617 8080 -4583
rect 8186 -4617 8224 -4583
rect 8258 -4617 8296 -4583
rect 8330 -4617 8341 -4583
rect 8402 -4617 8440 -4583
rect 8474 -4617 8512 -4583
rect 8546 -4617 8577 -4583
rect 8629 -4617 8656 -4583
rect 8690 -4617 8728 -4583
rect 8762 -4617 8800 -4583
rect 8865 -4617 8872 -4583
rect 8906 -4617 8944 -4583
rect 8978 -4617 9016 -4583
rect 9122 -4617 9160 -4583
rect 9194 -4617 9232 -4583
rect 9266 -4617 9285 -4583
rect 9338 -4617 9376 -4583
rect 9410 -4617 9448 -4583
rect 9482 -4617 9520 -4583
rect 9573 -4617 9592 -4583
rect 9626 -4617 9664 -4583
rect 9698 -4617 9736 -4583
rect 9842 -4617 9880 -4583
rect 9914 -4617 9952 -4583
rect 9986 -4617 9993 -4583
rect 10058 -4617 10096 -4583
rect 10130 -4617 10168 -4583
rect 10202 -4617 10229 -4583
rect 10281 -4617 10312 -4583
rect 10346 -4617 10384 -4583
rect 10418 -4617 10456 -4583
rect 10517 -4617 10528 -4583
rect 10562 -4617 10600 -4583
rect 10634 -4617 10672 -4583
rect 10778 -4617 10808 -4583
rect 4744 -4671 4801 -4617
rect 4853 -4671 5037 -4617
rect 5089 -4671 5273 -4617
rect 5325 -4671 5509 -4617
rect 5561 -4671 5745 -4617
rect 5797 -4671 5981 -4617
rect 6033 -4671 6217 -4617
rect 6269 -4671 6453 -4617
rect 6505 -4671 6689 -4617
rect 6741 -4671 6925 -4617
rect 6977 -4671 7161 -4617
rect 7213 -4671 7397 -4617
rect 7449 -4671 7633 -4617
rect 7685 -4671 7869 -4617
rect 7921 -4671 8105 -4617
rect 8157 -4671 8341 -4617
rect 8393 -4671 8577 -4617
rect 8629 -4671 8813 -4617
rect 8865 -4671 9049 -4617
rect 9101 -4671 9285 -4617
rect 9337 -4671 9521 -4617
rect 9573 -4671 9757 -4617
rect 9809 -4671 9993 -4617
rect 10045 -4671 10229 -4617
rect 10281 -4671 10465 -4617
rect 10517 -4671 10701 -4617
rect 10753 -4671 10808 -4617
rect 4744 -4705 4768 -4671
rect 4874 -4705 4912 -4671
rect 4946 -4705 4984 -4671
rect 5018 -4705 5037 -4671
rect 5090 -4705 5128 -4671
rect 5162 -4705 5200 -4671
rect 5234 -4705 5272 -4671
rect 5325 -4705 5344 -4671
rect 5378 -4705 5416 -4671
rect 5450 -4705 5488 -4671
rect 5594 -4705 5632 -4671
rect 5666 -4705 5704 -4671
rect 5738 -4705 5745 -4671
rect 5810 -4705 5848 -4671
rect 5882 -4705 5920 -4671
rect 5954 -4705 5981 -4671
rect 6033 -4705 6064 -4671
rect 6098 -4705 6136 -4671
rect 6170 -4705 6208 -4671
rect 6269 -4705 6280 -4671
rect 6314 -4705 6352 -4671
rect 6386 -4705 6424 -4671
rect 6530 -4705 6568 -4671
rect 6602 -4705 6640 -4671
rect 6674 -4705 6689 -4671
rect 6746 -4705 6784 -4671
rect 6818 -4705 6856 -4671
rect 6890 -4705 6925 -4671
rect 6977 -4705 7000 -4671
rect 7034 -4705 7072 -4671
rect 7106 -4705 7144 -4671
rect 7213 -4705 7216 -4671
rect 7250 -4705 7288 -4671
rect 7322 -4705 7360 -4671
rect 7394 -4705 7397 -4671
rect 7466 -4705 7504 -4671
rect 7538 -4705 7576 -4671
rect 7610 -4705 7633 -4671
rect 7685 -4705 7720 -4671
rect 7754 -4705 7792 -4671
rect 7826 -4705 7864 -4671
rect 7921 -4705 7936 -4671
rect 7970 -4705 8008 -4671
rect 8042 -4705 8080 -4671
rect 8186 -4705 8224 -4671
rect 8258 -4705 8296 -4671
rect 8330 -4705 8341 -4671
rect 8402 -4705 8440 -4671
rect 8474 -4705 8512 -4671
rect 8546 -4705 8577 -4671
rect 8629 -4705 8656 -4671
rect 8690 -4705 8728 -4671
rect 8762 -4705 8800 -4671
rect 8865 -4705 8872 -4671
rect 8906 -4705 8944 -4671
rect 8978 -4705 9016 -4671
rect 9122 -4705 9160 -4671
rect 9194 -4705 9232 -4671
rect 9266 -4705 9285 -4671
rect 9338 -4705 9376 -4671
rect 9410 -4705 9448 -4671
rect 9482 -4705 9520 -4671
rect 9573 -4705 9592 -4671
rect 9626 -4705 9664 -4671
rect 9698 -4705 9736 -4671
rect 9842 -4705 9880 -4671
rect 9914 -4705 9952 -4671
rect 9986 -4705 9993 -4671
rect 10058 -4705 10096 -4671
rect 10130 -4705 10168 -4671
rect 10202 -4705 10229 -4671
rect 10281 -4705 10312 -4671
rect 10346 -4705 10384 -4671
rect 10418 -4705 10456 -4671
rect 10517 -4705 10528 -4671
rect 10562 -4705 10600 -4671
rect 10634 -4705 10672 -4671
rect 10778 -4705 10808 -4671
rect 4744 -4725 4801 -4705
rect 4853 -4725 5037 -4705
rect 5089 -4725 5273 -4705
rect 5325 -4725 5509 -4705
rect 5561 -4725 5745 -4705
rect 5797 -4725 5981 -4705
rect 6033 -4725 6217 -4705
rect 6269 -4725 6453 -4705
rect 6505 -4725 6689 -4705
rect 6741 -4725 6925 -4705
rect 6977 -4725 7161 -4705
rect 7213 -4725 7397 -4705
rect 7449 -4725 7633 -4705
rect 7685 -4725 7869 -4705
rect 7921 -4725 8105 -4705
rect 8157 -4725 8341 -4705
rect 8393 -4725 8577 -4705
rect 8629 -4725 8813 -4705
rect 8865 -4725 9049 -4705
rect 9101 -4725 9285 -4705
rect 9337 -4725 9521 -4705
rect 9573 -4725 9757 -4705
rect 9809 -4725 9993 -4705
rect 10045 -4725 10229 -4705
rect 10281 -4725 10465 -4705
rect 10517 -4725 10701 -4705
rect 10753 -4725 10808 -4705
rect 5040 -4972 5086 -4960
rect 5040 -4980 5046 -4972
rect 5080 -4980 5086 -4972
rect 5158 -4972 5204 -4960
rect 5158 -4980 5164 -4972
rect 5198 -4980 5204 -4972
rect 5276 -4972 5322 -4960
rect 5276 -4980 5282 -4972
rect 5316 -4980 5322 -4972
rect 5394 -4972 5440 -4960
rect 5394 -4980 5400 -4972
rect 5434 -4980 5440 -4972
rect 5512 -4972 5558 -4960
rect 5512 -4980 5518 -4972
rect 5552 -4980 5558 -4972
rect 5630 -4972 5676 -4960
rect 5630 -4980 5636 -4972
rect 5670 -4980 5676 -4972
rect 5748 -4972 5794 -4960
rect 5748 -4980 5754 -4972
rect 5788 -4980 5794 -4972
rect 5866 -4972 5912 -4960
rect 5866 -4980 5872 -4972
rect 5906 -4980 5912 -4972
rect 5984 -4972 6030 -4960
rect 5984 -4980 5990 -4972
rect 6024 -4980 6030 -4972
rect 6102 -4972 6148 -4960
rect 6102 -4980 6108 -4972
rect 6142 -4980 6148 -4972
rect 6220 -4972 6266 -4960
rect 6220 -4980 6226 -4972
rect 6260 -4980 6266 -4972
rect 6338 -4972 6384 -4960
rect 6338 -4980 6344 -4972
rect 6378 -4980 6384 -4972
rect 6456 -4972 6502 -4960
rect 6456 -4980 6462 -4972
rect 6496 -4980 6502 -4972
rect 6574 -4972 6620 -4960
rect 6574 -4980 6580 -4972
rect 6614 -4980 6620 -4972
rect 6692 -4972 6738 -4960
rect 6692 -4980 6698 -4972
rect 6732 -4980 6738 -4972
rect 6810 -4972 6856 -4960
rect 6810 -4980 6816 -4972
rect 6850 -4980 6856 -4972
rect 6928 -4972 6974 -4960
rect 6928 -4980 6934 -4972
rect 6968 -4980 6974 -4972
rect 7046 -4972 7092 -4960
rect 7046 -4980 7052 -4972
rect 7086 -4980 7092 -4972
rect 7164 -4972 7210 -4960
rect 7164 -4980 7170 -4972
rect 7204 -4980 7210 -4972
rect 7282 -4972 7328 -4960
rect 7282 -4980 7288 -4972
rect 7322 -4980 7328 -4972
rect 7400 -4972 7446 -4960
rect 7400 -4980 7406 -4972
rect 7440 -4980 7446 -4972
rect 7518 -4972 7564 -4960
rect 7518 -4980 7524 -4972
rect 7558 -4980 7564 -4972
rect 7636 -4972 7682 -4960
rect 7636 -4980 7642 -4972
rect 7676 -4980 7682 -4972
rect 7754 -4972 7800 -4960
rect 7754 -4980 7760 -4972
rect 7794 -4980 7800 -4972
rect 7872 -4972 7918 -4960
rect 7872 -4980 7878 -4972
rect 7912 -4980 7918 -4972
rect 7990 -4972 8036 -4960
rect 7990 -4980 7996 -4972
rect 8030 -4980 8036 -4972
rect 8108 -4972 8154 -4960
rect 8108 -4980 8114 -4972
rect 8148 -4980 8154 -4972
rect 8226 -4972 8272 -4960
rect 8226 -4980 8232 -4972
rect 8266 -4980 8272 -4972
rect 8344 -4972 8390 -4960
rect 8344 -4980 8350 -4972
rect 8384 -4980 8390 -4972
rect 8462 -4972 8508 -4960
rect 8462 -4980 8468 -4972
rect 8502 -4980 8508 -4972
rect 8580 -4972 8626 -4960
rect 8580 -4980 8586 -4972
rect 8620 -4980 8626 -4972
rect 8698 -4972 8744 -4960
rect 8698 -4980 8704 -4972
rect 8738 -4980 8744 -4972
rect 8816 -4972 8862 -4960
rect 8816 -4980 8822 -4972
rect 8856 -4980 8862 -4972
rect 8934 -4972 8980 -4960
rect 8934 -4980 8940 -4972
rect 8974 -4980 8980 -4972
rect 9052 -4972 9098 -4960
rect 9052 -4980 9058 -4972
rect 9092 -4980 9098 -4972
rect 9170 -4972 9216 -4960
rect 9170 -4980 9176 -4972
rect 9210 -4980 9216 -4972
rect 9288 -4972 9334 -4960
rect 9288 -4980 9294 -4972
rect 9328 -4980 9334 -4972
rect 9406 -4972 9452 -4960
rect 9406 -4980 9412 -4972
rect 9446 -4980 9452 -4972
rect 9524 -4972 9570 -4960
rect 9524 -4980 9530 -4972
rect 9564 -4980 9570 -4972
rect 9642 -4972 9688 -4960
rect 9642 -4980 9648 -4972
rect 9682 -4980 9688 -4972
rect 9760 -4972 9806 -4960
rect 9760 -4980 9766 -4972
rect 9800 -4980 9806 -4972
rect 9878 -4972 9924 -4960
rect 9878 -4980 9884 -4972
rect 9918 -4980 9924 -4972
rect 9996 -4972 10042 -4960
rect 9996 -4980 10002 -4972
rect 10036 -4980 10042 -4972
rect 10114 -4972 10160 -4960
rect 10114 -4980 10120 -4972
rect 10154 -4980 10160 -4972
rect 10232 -4972 10278 -4960
rect 10232 -4980 10238 -4972
rect 10272 -4980 10278 -4972
rect 10350 -4972 10396 -4960
rect 10350 -4980 10356 -4972
rect 10390 -4980 10396 -4972
rect 10468 -4972 10514 -4960
rect 10468 -4980 10474 -4972
rect 10508 -4980 10514 -4972
rect 10586 -4972 10632 -4960
rect 10586 -4980 10592 -4972
rect 10626 -4980 10632 -4972
rect 10704 -4972 10750 -4960
rect 10704 -4980 10710 -4972
rect 10744 -4980 10750 -4972
rect 4791 -5540 4801 -4980
rect 4853 -5540 4863 -4980
rect 4911 -5540 4921 -4980
rect 4973 -5540 4983 -4980
rect 5027 -5540 5037 -4980
rect 5089 -5540 5099 -4980
rect 5147 -5540 5157 -4980
rect 5209 -5540 5219 -4980
rect 5263 -5540 5273 -4980
rect 5325 -5540 5335 -4980
rect 5383 -5540 5393 -4980
rect 5445 -5540 5455 -4980
rect 5499 -5540 5509 -4980
rect 5561 -5540 5571 -4980
rect 5619 -5540 5629 -4980
rect 5681 -5540 5691 -4980
rect 5735 -5540 5745 -4980
rect 5797 -5540 5807 -4980
rect 5855 -5540 5865 -4980
rect 5917 -5540 5927 -4980
rect 5971 -5540 5981 -4980
rect 6033 -5540 6043 -4980
rect 6091 -5540 6101 -4980
rect 6153 -5540 6163 -4980
rect 6207 -5540 6217 -4980
rect 6269 -5540 6279 -4980
rect 6327 -5540 6337 -4980
rect 6389 -5540 6399 -4980
rect 6443 -5540 6453 -4980
rect 6505 -5540 6515 -4980
rect 6563 -5540 6573 -4980
rect 6625 -5540 6635 -4980
rect 6679 -5540 6689 -4980
rect 6741 -5540 6751 -4980
rect 6799 -5540 6809 -4980
rect 6861 -5540 6871 -4980
rect 6915 -5540 6925 -4980
rect 6977 -5540 6987 -4980
rect 7035 -5540 7045 -4980
rect 7097 -5540 7107 -4980
rect 7151 -5540 7161 -4980
rect 7213 -5540 7223 -4980
rect 7271 -5540 7281 -4980
rect 7333 -5540 7343 -4980
rect 7387 -5540 7397 -4980
rect 7449 -5540 7459 -4980
rect 7507 -5540 7517 -4980
rect 7569 -5540 7579 -4980
rect 7623 -5540 7633 -4980
rect 7685 -5540 7695 -4980
rect 7743 -5540 7753 -4980
rect 7805 -5540 7815 -4980
rect 7859 -5540 7869 -4980
rect 7921 -5540 7931 -4980
rect 7979 -5540 7989 -4980
rect 8041 -5540 8051 -4980
rect 8095 -5540 8105 -4980
rect 8157 -5540 8167 -4980
rect 8215 -5540 8225 -4980
rect 8277 -5540 8287 -4980
rect 8331 -5540 8341 -4980
rect 8393 -5540 8403 -4980
rect 8451 -5540 8461 -4980
rect 8513 -5540 8523 -4980
rect 8567 -5540 8577 -4980
rect 8629 -5540 8639 -4980
rect 8687 -5540 8697 -4980
rect 8749 -5540 8759 -4980
rect 8803 -5540 8813 -4980
rect 8865 -5540 8875 -4980
rect 8923 -5540 8933 -4980
rect 8985 -5540 8995 -4980
rect 9039 -5540 9049 -4980
rect 9101 -5540 9111 -4980
rect 9159 -5540 9169 -4980
rect 9221 -5540 9231 -4980
rect 9275 -5540 9285 -4980
rect 9337 -5540 9347 -4980
rect 9395 -5540 9405 -4980
rect 9457 -5540 9467 -4980
rect 9511 -5540 9521 -4980
rect 9573 -5540 9583 -4980
rect 9631 -5540 9641 -4980
rect 9693 -5540 9703 -4980
rect 9747 -5540 9757 -4980
rect 9809 -5540 9819 -4980
rect 9867 -5540 9877 -4980
rect 9929 -5540 9939 -4980
rect 9983 -5540 9993 -4980
rect 10045 -5540 10055 -4980
rect 10103 -5540 10113 -4980
rect 10165 -5540 10175 -4980
rect 10219 -5540 10229 -4980
rect 10281 -5540 10291 -4980
rect 10339 -5540 10349 -4980
rect 10401 -5540 10411 -4980
rect 10455 -5540 10465 -4980
rect 10517 -5540 10527 -4980
rect 10575 -5540 10585 -4980
rect 10637 -5540 10647 -4980
rect 10691 -5540 10701 -4980
rect 10753 -5540 10763 -4980
rect 5040 -5548 5046 -5540
rect 5080 -5548 5086 -5540
rect 5040 -5560 5086 -5548
rect 5158 -5548 5164 -5540
rect 5198 -5548 5204 -5540
rect 5158 -5560 5204 -5548
rect 5276 -5548 5282 -5540
rect 5316 -5548 5322 -5540
rect 5276 -5560 5322 -5548
rect 5394 -5548 5400 -5540
rect 5434 -5548 5440 -5540
rect 5394 -5560 5440 -5548
rect 5512 -5548 5518 -5540
rect 5552 -5548 5558 -5540
rect 5512 -5560 5558 -5548
rect 5630 -5548 5636 -5540
rect 5670 -5548 5676 -5540
rect 5630 -5560 5676 -5548
rect 5748 -5548 5754 -5540
rect 5788 -5548 5794 -5540
rect 5748 -5560 5794 -5548
rect 5866 -5548 5872 -5540
rect 5906 -5548 5912 -5540
rect 5866 -5560 5912 -5548
rect 5984 -5548 5990 -5540
rect 6024 -5548 6030 -5540
rect 5984 -5560 6030 -5548
rect 6102 -5548 6108 -5540
rect 6142 -5548 6148 -5540
rect 6102 -5560 6148 -5548
rect 6220 -5548 6226 -5540
rect 6260 -5548 6266 -5540
rect 6220 -5560 6266 -5548
rect 6338 -5548 6344 -5540
rect 6378 -5548 6384 -5540
rect 6338 -5560 6384 -5548
rect 6456 -5548 6462 -5540
rect 6496 -5548 6502 -5540
rect 6456 -5560 6502 -5548
rect 6574 -5548 6580 -5540
rect 6614 -5548 6620 -5540
rect 6574 -5560 6620 -5548
rect 6692 -5548 6698 -5540
rect 6732 -5548 6738 -5540
rect 6692 -5560 6738 -5548
rect 6810 -5548 6816 -5540
rect 6850 -5548 6856 -5540
rect 6810 -5560 6856 -5548
rect 6928 -5548 6934 -5540
rect 6968 -5548 6974 -5540
rect 6928 -5560 6974 -5548
rect 7046 -5548 7052 -5540
rect 7086 -5548 7092 -5540
rect 7046 -5560 7092 -5548
rect 7164 -5548 7170 -5540
rect 7204 -5548 7210 -5540
rect 7164 -5560 7210 -5548
rect 7282 -5548 7288 -5540
rect 7322 -5548 7328 -5540
rect 7282 -5560 7328 -5548
rect 7400 -5548 7406 -5540
rect 7440 -5548 7446 -5540
rect 7400 -5560 7446 -5548
rect 7518 -5548 7524 -5540
rect 7558 -5548 7564 -5540
rect 7518 -5560 7564 -5548
rect 7636 -5548 7642 -5540
rect 7676 -5548 7682 -5540
rect 7636 -5560 7682 -5548
rect 7754 -5548 7760 -5540
rect 7794 -5548 7800 -5540
rect 7754 -5560 7800 -5548
rect 7872 -5548 7878 -5540
rect 7912 -5548 7918 -5540
rect 7872 -5560 7918 -5548
rect 7990 -5548 7996 -5540
rect 8030 -5548 8036 -5540
rect 7990 -5560 8036 -5548
rect 8108 -5548 8114 -5540
rect 8148 -5548 8154 -5540
rect 8108 -5560 8154 -5548
rect 8226 -5548 8232 -5540
rect 8266 -5548 8272 -5540
rect 8226 -5560 8272 -5548
rect 8344 -5548 8350 -5540
rect 8384 -5548 8390 -5540
rect 8344 -5560 8390 -5548
rect 8462 -5548 8468 -5540
rect 8502 -5548 8508 -5540
rect 8462 -5560 8508 -5548
rect 8580 -5548 8586 -5540
rect 8620 -5548 8626 -5540
rect 8580 -5560 8626 -5548
rect 8698 -5548 8704 -5540
rect 8738 -5548 8744 -5540
rect 8698 -5560 8744 -5548
rect 8816 -5548 8822 -5540
rect 8856 -5548 8862 -5540
rect 8816 -5560 8862 -5548
rect 8934 -5548 8940 -5540
rect 8974 -5548 8980 -5540
rect 8934 -5560 8980 -5548
rect 9052 -5548 9058 -5540
rect 9092 -5548 9098 -5540
rect 9052 -5560 9098 -5548
rect 9170 -5548 9176 -5540
rect 9210 -5548 9216 -5540
rect 9170 -5560 9216 -5548
rect 9288 -5548 9294 -5540
rect 9328 -5548 9334 -5540
rect 9288 -5560 9334 -5548
rect 9406 -5548 9412 -5540
rect 9446 -5548 9452 -5540
rect 9406 -5560 9452 -5548
rect 9524 -5548 9530 -5540
rect 9564 -5548 9570 -5540
rect 9524 -5560 9570 -5548
rect 9642 -5548 9648 -5540
rect 9682 -5548 9688 -5540
rect 9642 -5560 9688 -5548
rect 9760 -5548 9766 -5540
rect 9800 -5548 9806 -5540
rect 9760 -5560 9806 -5548
rect 9878 -5548 9884 -5540
rect 9918 -5548 9924 -5540
rect 9878 -5560 9924 -5548
rect 9996 -5548 10002 -5540
rect 10036 -5548 10042 -5540
rect 9996 -5560 10042 -5548
rect 10114 -5548 10120 -5540
rect 10154 -5548 10160 -5540
rect 10114 -5560 10160 -5548
rect 10232 -5548 10238 -5540
rect 10272 -5548 10278 -5540
rect 10232 -5560 10278 -5548
rect 10350 -5548 10356 -5540
rect 10390 -5548 10396 -5540
rect 10350 -5560 10396 -5548
rect 10468 -5548 10474 -5540
rect 10508 -5548 10514 -5540
rect 10468 -5560 10514 -5548
rect 10586 -5548 10592 -5540
rect 10626 -5548 10632 -5540
rect 10586 -5560 10632 -5548
rect 10704 -5548 10710 -5540
rect 10744 -5548 10750 -5540
rect 10704 -5560 10750 -5548
rect 4847 -5755 4857 -5601
rect 4915 -5755 4925 -5601
rect 4965 -5755 4975 -5601
rect 5033 -5755 5043 -5601
rect 5083 -5755 5093 -5601
rect 5151 -5755 5161 -5601
rect 5201 -5755 5211 -5601
rect 5269 -5755 5279 -5601
rect 5319 -5755 5329 -5601
rect 5387 -5755 5397 -5601
rect 5437 -5755 5447 -5601
rect 5505 -5755 5515 -5601
rect 5555 -5755 5565 -5601
rect 5623 -5755 5633 -5601
rect 5673 -5755 5683 -5601
rect 5741 -5755 5751 -5601
rect 5791 -5755 5801 -5601
rect 5859 -5755 5869 -5601
rect 5909 -5755 5919 -5601
rect 5977 -5755 5987 -5601
rect 6027 -5755 6037 -5601
rect 6095 -5755 6105 -5601
rect 6145 -5755 6155 -5601
rect 6213 -5755 6223 -5601
rect 6263 -5755 6273 -5601
rect 6331 -5755 6341 -5601
rect 6381 -5755 6391 -5601
rect 6449 -5755 6459 -5601
rect 6499 -5755 6509 -5601
rect 6567 -5755 6577 -5601
rect 6617 -5755 6627 -5601
rect 6685 -5755 6695 -5601
rect 6735 -5755 6745 -5601
rect 6803 -5755 6813 -5601
rect 6853 -5755 6863 -5601
rect 6921 -5755 6931 -5601
rect 6971 -5755 6981 -5601
rect 7039 -5755 7049 -5601
rect 7089 -5755 7099 -5601
rect 7157 -5755 7167 -5601
rect 7207 -5755 7217 -5601
rect 7275 -5755 7285 -5601
rect 7325 -5755 7335 -5601
rect 7393 -5755 7403 -5601
rect 7443 -5755 7453 -5601
rect 7511 -5755 7521 -5601
rect 7561 -5755 7571 -5601
rect 7629 -5755 7639 -5601
rect 7679 -5755 7689 -5601
rect 7747 -5755 7757 -5601
rect 7797 -5755 7807 -5601
rect 7865 -5755 7875 -5601
rect 7915 -5755 7925 -5601
rect 7983 -5755 7993 -5601
rect 8033 -5755 8043 -5601
rect 8101 -5755 8111 -5601
rect 8151 -5755 8161 -5601
rect 8219 -5755 8229 -5601
rect 8269 -5755 8279 -5601
rect 8337 -5755 8347 -5601
rect 8387 -5755 8397 -5601
rect 8455 -5755 8465 -5601
rect 8505 -5755 8515 -5601
rect 8573 -5755 8583 -5601
rect 8623 -5755 8633 -5601
rect 8691 -5755 8701 -5601
rect 8741 -5755 8751 -5601
rect 8809 -5755 8819 -5601
rect 8859 -5755 8869 -5601
rect 8927 -5755 8937 -5601
rect 8977 -5755 8987 -5601
rect 9045 -5755 9055 -5601
rect 9095 -5755 9105 -5601
rect 9163 -5755 9173 -5601
rect 9213 -5755 9223 -5601
rect 9281 -5755 9291 -5601
rect 9331 -5755 9341 -5601
rect 9399 -5755 9409 -5601
rect 9449 -5755 9459 -5601
rect 9517 -5755 9527 -5601
rect 9567 -5755 9577 -5601
rect 9635 -5755 9645 -5601
rect 9685 -5755 9695 -5601
rect 9753 -5755 9763 -5601
rect 9803 -5755 9813 -5601
rect 9871 -5755 9881 -5601
rect 9921 -5755 9931 -5601
rect 9989 -5755 9999 -5601
rect 10039 -5755 10049 -5601
rect 10107 -5755 10117 -5601
rect 10157 -5755 10167 -5601
rect 10225 -5755 10235 -5601
rect 10275 -5755 10285 -5601
rect 10343 -5755 10353 -5601
rect 10393 -5755 10403 -5601
rect 10461 -5755 10471 -5601
rect 10511 -5755 10521 -5601
rect 10579 -5755 10589 -5601
rect 10629 -5755 10639 -5601
rect 10697 -5755 10707 -5601
rect 4804 -5808 4850 -5796
rect 4804 -5816 4810 -5808
rect 4844 -5816 4850 -5808
rect 4922 -5808 4968 -5796
rect 4922 -5816 4928 -5808
rect 4962 -5816 4968 -5808
rect 5040 -5808 5086 -5796
rect 5040 -5816 5046 -5808
rect 5080 -5816 5086 -5808
rect 5158 -5808 5204 -5796
rect 5158 -5816 5164 -5808
rect 5198 -5816 5204 -5808
rect 5276 -5808 5322 -5796
rect 5276 -5816 5282 -5808
rect 5316 -5816 5322 -5808
rect 5394 -5808 5440 -5796
rect 5394 -5816 5400 -5808
rect 5434 -5816 5440 -5808
rect 5512 -5808 5558 -5796
rect 5512 -5816 5518 -5808
rect 5552 -5816 5558 -5808
rect 5630 -5808 5676 -5796
rect 5630 -5816 5636 -5808
rect 5670 -5816 5676 -5808
rect 5748 -5808 5794 -5796
rect 5748 -5816 5754 -5808
rect 5788 -5816 5794 -5808
rect 5866 -5808 5912 -5796
rect 5866 -5816 5872 -5808
rect 5906 -5816 5912 -5808
rect 5984 -5808 6030 -5796
rect 5984 -5816 5990 -5808
rect 6024 -5816 6030 -5808
rect 6102 -5808 6148 -5796
rect 6102 -5816 6108 -5808
rect 6142 -5816 6148 -5808
rect 6220 -5808 6266 -5796
rect 6220 -5816 6226 -5808
rect 6260 -5816 6266 -5808
rect 6338 -5808 6384 -5796
rect 6338 -5816 6344 -5808
rect 6378 -5816 6384 -5808
rect 6456 -5808 6502 -5796
rect 6456 -5816 6462 -5808
rect 6496 -5816 6502 -5808
rect 6574 -5808 6620 -5796
rect 6574 -5816 6580 -5808
rect 6614 -5816 6620 -5808
rect 6692 -5808 6738 -5796
rect 6692 -5816 6698 -5808
rect 6732 -5816 6738 -5808
rect 6810 -5808 6856 -5796
rect 6810 -5816 6816 -5808
rect 6850 -5816 6856 -5808
rect 6928 -5808 6974 -5796
rect 6928 -5816 6934 -5808
rect 6968 -5816 6974 -5808
rect 7046 -5808 7092 -5796
rect 7046 -5816 7052 -5808
rect 7086 -5816 7092 -5808
rect 7164 -5808 7210 -5796
rect 7164 -5816 7170 -5808
rect 7204 -5816 7210 -5808
rect 7282 -5808 7328 -5796
rect 7282 -5816 7288 -5808
rect 7322 -5816 7328 -5808
rect 7400 -5808 7446 -5796
rect 7400 -5816 7406 -5808
rect 7440 -5816 7446 -5808
rect 7518 -5808 7564 -5796
rect 7518 -5816 7524 -5808
rect 7558 -5816 7564 -5808
rect 7636 -5808 7682 -5796
rect 7636 -5816 7642 -5808
rect 7676 -5816 7682 -5808
rect 7754 -5808 7800 -5796
rect 7754 -5816 7760 -5808
rect 7794 -5816 7800 -5808
rect 7872 -5808 7918 -5796
rect 7872 -5816 7878 -5808
rect 7912 -5816 7918 -5808
rect 7990 -5808 8036 -5796
rect 7990 -5816 7996 -5808
rect 8030 -5816 8036 -5808
rect 8108 -5808 8154 -5796
rect 8108 -5816 8114 -5808
rect 8148 -5816 8154 -5808
rect 8226 -5808 8272 -5796
rect 8226 -5816 8232 -5808
rect 8266 -5816 8272 -5808
rect 8344 -5808 8390 -5796
rect 8344 -5816 8350 -5808
rect 8384 -5816 8390 -5808
rect 8462 -5808 8508 -5796
rect 8462 -5816 8468 -5808
rect 8502 -5816 8508 -5808
rect 8580 -5808 8626 -5796
rect 8580 -5816 8586 -5808
rect 8620 -5816 8626 -5808
rect 8698 -5808 8744 -5796
rect 8698 -5816 8704 -5808
rect 8738 -5816 8744 -5808
rect 8816 -5808 8862 -5796
rect 8816 -5816 8822 -5808
rect 8856 -5816 8862 -5808
rect 8934 -5808 8980 -5796
rect 8934 -5816 8940 -5808
rect 8974 -5816 8980 -5808
rect 9052 -5808 9098 -5796
rect 9052 -5816 9058 -5808
rect 9092 -5816 9098 -5808
rect 9170 -5808 9216 -5796
rect 9170 -5816 9176 -5808
rect 9210 -5816 9216 -5808
rect 9288 -5808 9334 -5796
rect 9288 -5816 9294 -5808
rect 9328 -5816 9334 -5808
rect 9406 -5808 9452 -5796
rect 9406 -5816 9412 -5808
rect 9446 -5816 9452 -5808
rect 9524 -5808 9570 -5796
rect 9524 -5816 9530 -5808
rect 9564 -5816 9570 -5808
rect 9642 -5808 9688 -5796
rect 9642 -5816 9648 -5808
rect 9682 -5816 9688 -5808
rect 9760 -5808 9806 -5796
rect 9760 -5816 9766 -5808
rect 9800 -5816 9806 -5808
rect 9878 -5808 9924 -5796
rect 9878 -5816 9884 -5808
rect 9918 -5816 9924 -5808
rect 9996 -5808 10042 -5796
rect 9996 -5816 10002 -5808
rect 10036 -5816 10042 -5808
rect 10114 -5808 10160 -5796
rect 10114 -5816 10120 -5808
rect 10154 -5816 10160 -5808
rect 10232 -5808 10278 -5796
rect 10232 -5816 10238 -5808
rect 10272 -5816 10278 -5808
rect 10350 -5808 10396 -5796
rect 10350 -5816 10356 -5808
rect 10390 -5816 10396 -5808
rect 10468 -5808 10514 -5796
rect 10468 -5816 10474 -5808
rect 10508 -5816 10514 -5808
rect 10586 -5808 10632 -5796
rect 10586 -5816 10592 -5808
rect 10626 -5816 10632 -5808
rect 10704 -5808 10750 -5796
rect 10704 -5816 10710 -5808
rect 10744 -5816 10750 -5808
rect 4791 -6376 4801 -5816
rect 4853 -6376 4863 -5816
rect 4911 -6376 4921 -5816
rect 4973 -6376 4983 -5816
rect 5027 -6376 5037 -5816
rect 5089 -6376 5099 -5816
rect 5147 -6376 5157 -5816
rect 5209 -6376 5219 -5816
rect 5263 -6376 5273 -5816
rect 5325 -6376 5335 -5816
rect 5383 -6376 5393 -5816
rect 5445 -6376 5455 -5816
rect 5499 -6376 5509 -5816
rect 5561 -6376 5571 -5816
rect 5619 -6376 5629 -5816
rect 5681 -6376 5691 -5816
rect 5735 -6376 5745 -5816
rect 5797 -6376 5807 -5816
rect 5855 -6376 5865 -5816
rect 5917 -6376 5927 -5816
rect 5971 -6376 5981 -5816
rect 6033 -6376 6043 -5816
rect 6091 -6376 6101 -5816
rect 6153 -6376 6163 -5816
rect 6207 -6376 6217 -5816
rect 6269 -6376 6279 -5816
rect 6327 -6376 6337 -5816
rect 6389 -6376 6399 -5816
rect 6443 -6376 6453 -5816
rect 6505 -6376 6515 -5816
rect 6563 -6376 6573 -5816
rect 6625 -6376 6635 -5816
rect 6679 -6376 6689 -5816
rect 6741 -6376 6751 -5816
rect 6799 -6376 6809 -5816
rect 6861 -6376 6871 -5816
rect 6915 -6376 6925 -5816
rect 6977 -6376 6987 -5816
rect 7035 -6376 7045 -5816
rect 7097 -6376 7107 -5816
rect 7151 -6376 7161 -5816
rect 7213 -6376 7223 -5816
rect 7271 -6376 7281 -5816
rect 7333 -6376 7343 -5816
rect 7387 -6376 7397 -5816
rect 7449 -6376 7459 -5816
rect 7507 -6376 7517 -5816
rect 7569 -6376 7579 -5816
rect 7623 -6376 7633 -5816
rect 7685 -6376 7695 -5816
rect 7743 -6376 7753 -5816
rect 7805 -6376 7815 -5816
rect 7859 -6376 7869 -5816
rect 7921 -6376 7931 -5816
rect 7979 -6376 7989 -5816
rect 8041 -6376 8051 -5816
rect 8095 -6376 8105 -5816
rect 8157 -6376 8167 -5816
rect 8215 -6376 8225 -5816
rect 8277 -6376 8287 -5816
rect 8331 -6376 8341 -5816
rect 8393 -6376 8403 -5816
rect 8451 -6376 8461 -5816
rect 8513 -6376 8523 -5816
rect 8567 -6376 8577 -5816
rect 8629 -6376 8639 -5816
rect 8687 -6376 8697 -5816
rect 8749 -6376 8759 -5816
rect 8803 -6376 8813 -5816
rect 8865 -6376 8875 -5816
rect 8923 -6376 8933 -5816
rect 8985 -6376 8995 -5816
rect 9039 -6376 9049 -5816
rect 9101 -6376 9111 -5816
rect 9159 -6376 9169 -5816
rect 9221 -6376 9231 -5816
rect 9275 -6376 9285 -5816
rect 9337 -6376 9347 -5816
rect 9395 -6376 9405 -5816
rect 9457 -6376 9467 -5816
rect 9511 -6376 9521 -5816
rect 9573 -6376 9583 -5816
rect 9631 -6376 9641 -5816
rect 9693 -6376 9703 -5816
rect 9747 -6376 9757 -5816
rect 9809 -6376 9819 -5816
rect 9867 -6376 9877 -5816
rect 9929 -6376 9939 -5816
rect 9983 -6376 9993 -5816
rect 10045 -6376 10055 -5816
rect 10103 -6376 10113 -5816
rect 10165 -6376 10175 -5816
rect 10219 -6376 10229 -5816
rect 10281 -6376 10291 -5816
rect 10339 -6376 10349 -5816
rect 10401 -6376 10411 -5816
rect 10455 -6376 10465 -5816
rect 10517 -6376 10527 -5816
rect 10575 -6376 10585 -5816
rect 10637 -6376 10647 -5816
rect 10691 -6376 10701 -5816
rect 10753 -6376 10763 -5816
rect 4804 -6384 4810 -6376
rect 4844 -6384 4850 -6376
rect 4804 -6396 4850 -6384
rect 4922 -6384 4928 -6376
rect 4962 -6384 4968 -6376
rect 4922 -6396 4968 -6384
rect 5040 -6384 5046 -6376
rect 5080 -6384 5086 -6376
rect 5040 -6396 5086 -6384
rect 5158 -6384 5164 -6376
rect 5198 -6384 5204 -6376
rect 5158 -6396 5204 -6384
rect 5276 -6384 5282 -6376
rect 5316 -6384 5322 -6376
rect 5276 -6396 5322 -6384
rect 5394 -6384 5400 -6376
rect 5434 -6384 5440 -6376
rect 5394 -6396 5440 -6384
rect 5512 -6384 5518 -6376
rect 5552 -6384 5558 -6376
rect 5512 -6396 5558 -6384
rect 5630 -6384 5636 -6376
rect 5670 -6384 5676 -6376
rect 5630 -6396 5676 -6384
rect 5748 -6384 5754 -6376
rect 5788 -6384 5794 -6376
rect 5748 -6396 5794 -6384
rect 5866 -6384 5872 -6376
rect 5906 -6384 5912 -6376
rect 5866 -6396 5912 -6384
rect 5984 -6384 5990 -6376
rect 6024 -6384 6030 -6376
rect 5984 -6396 6030 -6384
rect 6102 -6384 6108 -6376
rect 6142 -6384 6148 -6376
rect 6102 -6396 6148 -6384
rect 6220 -6384 6226 -6376
rect 6260 -6384 6266 -6376
rect 6220 -6396 6266 -6384
rect 6338 -6384 6344 -6376
rect 6378 -6384 6384 -6376
rect 6338 -6396 6384 -6384
rect 6456 -6384 6462 -6376
rect 6496 -6384 6502 -6376
rect 6456 -6396 6502 -6384
rect 6574 -6384 6580 -6376
rect 6614 -6384 6620 -6376
rect 6574 -6396 6620 -6384
rect 6692 -6384 6698 -6376
rect 6732 -6384 6738 -6376
rect 6692 -6396 6738 -6384
rect 6810 -6384 6816 -6376
rect 6850 -6384 6856 -6376
rect 6810 -6396 6856 -6384
rect 6928 -6384 6934 -6376
rect 6968 -6384 6974 -6376
rect 6928 -6396 6974 -6384
rect 7046 -6384 7052 -6376
rect 7086 -6384 7092 -6376
rect 7046 -6396 7092 -6384
rect 7164 -6384 7170 -6376
rect 7204 -6384 7210 -6376
rect 7164 -6396 7210 -6384
rect 7282 -6384 7288 -6376
rect 7322 -6384 7328 -6376
rect 7282 -6396 7328 -6384
rect 7400 -6384 7406 -6376
rect 7440 -6384 7446 -6376
rect 7400 -6396 7446 -6384
rect 7518 -6384 7524 -6376
rect 7558 -6384 7564 -6376
rect 7518 -6396 7564 -6384
rect 7636 -6384 7642 -6376
rect 7676 -6384 7682 -6376
rect 7636 -6396 7682 -6384
rect 7754 -6384 7760 -6376
rect 7794 -6384 7800 -6376
rect 7754 -6396 7800 -6384
rect 7872 -6384 7878 -6376
rect 7912 -6384 7918 -6376
rect 7872 -6396 7918 -6384
rect 7990 -6384 7996 -6376
rect 8030 -6384 8036 -6376
rect 7990 -6396 8036 -6384
rect 8108 -6384 8114 -6376
rect 8148 -6384 8154 -6376
rect 8108 -6396 8154 -6384
rect 8226 -6384 8232 -6376
rect 8266 -6384 8272 -6376
rect 8226 -6396 8272 -6384
rect 8344 -6384 8350 -6376
rect 8384 -6384 8390 -6376
rect 8344 -6396 8390 -6384
rect 8462 -6384 8468 -6376
rect 8502 -6384 8508 -6376
rect 8462 -6396 8508 -6384
rect 8580 -6384 8586 -6376
rect 8620 -6384 8626 -6376
rect 8580 -6396 8626 -6384
rect 8698 -6384 8704 -6376
rect 8738 -6384 8744 -6376
rect 8698 -6396 8744 -6384
rect 8816 -6384 8822 -6376
rect 8856 -6384 8862 -6376
rect 8816 -6396 8862 -6384
rect 8934 -6384 8940 -6376
rect 8974 -6384 8980 -6376
rect 8934 -6396 8980 -6384
rect 9052 -6384 9058 -6376
rect 9092 -6384 9098 -6376
rect 9052 -6396 9098 -6384
rect 9170 -6384 9176 -6376
rect 9210 -6384 9216 -6376
rect 9170 -6396 9216 -6384
rect 9288 -6384 9294 -6376
rect 9328 -6384 9334 -6376
rect 9288 -6396 9334 -6384
rect 9406 -6384 9412 -6376
rect 9446 -6384 9452 -6376
rect 9406 -6396 9452 -6384
rect 9524 -6384 9530 -6376
rect 9564 -6384 9570 -6376
rect 9524 -6396 9570 -6384
rect 9642 -6384 9648 -6376
rect 9682 -6384 9688 -6376
rect 9642 -6396 9688 -6384
rect 9760 -6384 9766 -6376
rect 9800 -6384 9806 -6376
rect 9760 -6396 9806 -6384
rect 9878 -6384 9884 -6376
rect 9918 -6384 9924 -6376
rect 9878 -6396 9924 -6384
rect 9996 -6384 10002 -6376
rect 10036 -6384 10042 -6376
rect 9996 -6396 10042 -6384
rect 10114 -6384 10120 -6376
rect 10154 -6384 10160 -6376
rect 10114 -6396 10160 -6384
rect 10232 -6384 10238 -6376
rect 10272 -6384 10278 -6376
rect 10232 -6396 10278 -6384
rect 10350 -6384 10356 -6376
rect 10390 -6384 10396 -6376
rect 10350 -6396 10396 -6384
rect 10468 -6384 10474 -6376
rect 10508 -6384 10514 -6376
rect 10468 -6396 10514 -6384
rect 10586 -6384 10592 -6376
rect 10626 -6384 10632 -6376
rect 10586 -6396 10632 -6384
rect 10704 -6384 10710 -6376
rect 10744 -6384 10750 -6376
rect 10704 -6396 10750 -6384
rect 4582 -6456 4740 -6438
rect 4582 -6510 4656 -6456
rect 4666 -6510 4740 -6456
rect 4675 -6599 4760 -6510
rect 4791 -6599 4801 -6525
rect 4675 -6701 4801 -6599
rect 4675 -6775 4760 -6701
rect 4791 -6775 4801 -6701
rect 4853 -6599 4863 -6525
rect 4853 -6701 5037 -6599
rect 4853 -6775 4863 -6701
rect 5089 -6701 5273 -6599
rect 5325 -6701 5509 -6599
rect 5561 -6701 5745 -6599
rect 5797 -6701 5981 -6599
rect 6033 -6701 6217 -6599
rect 6269 -6701 6453 -6599
rect 6505 -6701 6689 -6599
rect 6741 -6701 6925 -6599
rect 6977 -6701 7161 -6599
rect 7213 -6701 7397 -6599
rect 7449 -6701 7633 -6599
rect 7685 -6701 7869 -6599
rect 7921 -6701 8105 -6599
rect 8157 -6701 8341 -6599
rect 8393 -6701 8577 -6599
rect 8629 -6701 8813 -6599
rect 8865 -6701 9049 -6599
rect 9101 -6701 9285 -6599
rect 9337 -6701 9521 -6599
rect 9573 -6701 9757 -6599
rect 9809 -6701 9993 -6599
rect 10045 -6701 10229 -6599
rect 10281 -6701 10465 -6599
rect 10517 -6701 10701 -6599
rect 10805 -6599 11600 -6524
rect 10753 -6655 11600 -6599
rect 10753 -6701 10902 -6655
rect 10808 -6775 10902 -6701
rect 11054 -6752 11068 -6700
rect 11120 -6752 11149 -6700
rect 11201 -6752 11230 -6700
rect 11282 -6752 11311 -6700
rect 11363 -6752 11392 -6700
rect 11444 -6752 11473 -6700
rect 11525 -6752 11554 -6700
rect 11606 -6752 11621 -6700
rect 11054 -6804 11621 -6752
rect 11054 -6856 11068 -6804
rect 11120 -6856 11149 -6804
rect 11201 -6856 11230 -6804
rect 11282 -6856 11311 -6804
rect 11363 -6856 11392 -6804
rect 11444 -6856 11473 -6804
rect 11525 -6856 11554 -6804
rect 11606 -6856 11621 -6804
rect 9794 -6928 10626 -6860
rect 11054 -6908 11621 -6856
rect 5745 -6942 10875 -6928
rect 5745 -6994 5759 -6942
rect 5811 -6994 5839 -6942
rect 5891 -6994 5919 -6942
rect 5971 -6994 5999 -6942
rect 6051 -6994 6079 -6942
rect 6131 -6994 6159 -6942
rect 6211 -6994 6239 -6942
rect 6291 -6994 6319 -6942
rect 6371 -6994 6399 -6942
rect 6451 -6994 6479 -6942
rect 6531 -6994 6559 -6942
rect 6611 -6994 6639 -6942
rect 6691 -6994 6719 -6942
rect 6771 -6994 6799 -6942
rect 6851 -6994 6879 -6942
rect 6931 -6994 6959 -6942
rect 7011 -6994 7039 -6942
rect 7091 -6994 7119 -6942
rect 7171 -6994 7199 -6942
rect 7251 -6994 7279 -6942
rect 7331 -6994 7359 -6942
rect 7411 -6994 7439 -6942
rect 7491 -6994 7519 -6942
rect 7571 -6994 7599 -6942
rect 7651 -6994 7679 -6942
rect 7731 -6994 7759 -6942
rect 7811 -6994 7839 -6942
rect 7891 -6994 7919 -6942
rect 7971 -6994 7999 -6942
rect 8051 -6994 8079 -6942
rect 8131 -6994 8159 -6942
rect 8211 -6994 8239 -6942
rect 8291 -6994 8319 -6942
rect 8371 -6994 8399 -6942
rect 8451 -6994 8479 -6942
rect 8531 -6994 8559 -6942
rect 8611 -6994 8639 -6942
rect 8691 -6994 8719 -6942
rect 8771 -6994 8799 -6942
rect 8851 -6994 8879 -6942
rect 8931 -6994 8959 -6942
rect 9011 -6994 9039 -6942
rect 9091 -6994 9119 -6942
rect 9171 -6994 9199 -6942
rect 9251 -6994 9279 -6942
rect 9331 -6994 9359 -6942
rect 9411 -6994 9439 -6942
rect 9491 -6994 9519 -6942
rect 9571 -6994 9599 -6942
rect 9651 -6994 9679 -6942
rect 9731 -6994 9759 -6942
rect 9811 -6994 9839 -6942
rect 9891 -6994 9919 -6942
rect 9971 -6994 9999 -6942
rect 10051 -6994 10079 -6942
rect 10131 -6994 10159 -6942
rect 10211 -6994 10239 -6942
rect 10291 -6994 10319 -6942
rect 10371 -6994 10399 -6942
rect 10451 -6994 10479 -6942
rect 10531 -6994 10559 -6942
rect 10611 -6994 10639 -6942
rect 10691 -6994 10719 -6942
rect 10771 -6994 10799 -6942
rect 10851 -6994 10875 -6942
rect 11054 -6960 11068 -6908
rect 11120 -6960 11149 -6908
rect 11201 -6960 11230 -6908
rect 11282 -6960 11311 -6908
rect 11363 -6960 11392 -6908
rect 11444 -6960 11473 -6908
rect 11525 -6960 11554 -6908
rect 11606 -6960 11621 -6908
rect 5745 -7022 10875 -6994
rect 4060 -7063 5610 -7035
rect 4060 -7115 4094 -7063
rect 4146 -7115 4175 -7063
rect 4227 -7115 4256 -7063
rect 4308 -7115 4337 -7063
rect 4389 -7115 4418 -7063
rect 4470 -7115 4499 -7063
rect 4551 -7115 4580 -7063
rect 4632 -7115 4662 -7063
rect 4714 -7115 4743 -7063
rect 4795 -7115 4824 -7063
rect 4876 -7115 4905 -7063
rect 4957 -7115 4986 -7063
rect 5038 -7115 5067 -7063
rect 5119 -7115 5148 -7063
rect 5200 -7115 5230 -7063
rect 5282 -7115 5311 -7063
rect 5363 -7115 5392 -7063
rect 5444 -7115 5610 -7063
rect 5745 -7074 5759 -7022
rect 5811 -7074 5839 -7022
rect 5891 -7074 5919 -7022
rect 5971 -7074 5999 -7022
rect 6051 -7074 6079 -7022
rect 6131 -7074 6159 -7022
rect 6211 -7074 6239 -7022
rect 6291 -7074 6319 -7022
rect 6371 -7074 6399 -7022
rect 6451 -7074 6479 -7022
rect 6531 -7074 6559 -7022
rect 6611 -7074 6639 -7022
rect 6691 -7074 6719 -7022
rect 6771 -7074 6799 -7022
rect 6851 -7074 6879 -7022
rect 6931 -7074 6959 -7022
rect 7011 -7074 7039 -7022
rect 7091 -7074 7119 -7022
rect 7171 -7074 7199 -7022
rect 7251 -7074 7279 -7022
rect 7331 -7074 7359 -7022
rect 7411 -7074 7439 -7022
rect 7491 -7074 7519 -7022
rect 7571 -7074 7599 -7022
rect 7651 -7074 7679 -7022
rect 7731 -7074 7759 -7022
rect 7811 -7074 7839 -7022
rect 7891 -7074 7919 -7022
rect 7971 -7074 7999 -7022
rect 8051 -7074 8079 -7022
rect 8131 -7074 8159 -7022
rect 8211 -7074 8239 -7022
rect 8291 -7074 8319 -7022
rect 8371 -7074 8399 -7022
rect 8451 -7074 8479 -7022
rect 8531 -7074 8559 -7022
rect 8611 -7074 8639 -7022
rect 8691 -7074 8719 -7022
rect 8771 -7074 8799 -7022
rect 8851 -7074 8879 -7022
rect 8931 -7074 8959 -7022
rect 9011 -7074 9039 -7022
rect 9091 -7074 9119 -7022
rect 9171 -7074 9199 -7022
rect 9251 -7074 9279 -7022
rect 9331 -7074 9359 -7022
rect 9411 -7074 9439 -7022
rect 9491 -7074 9519 -7022
rect 9571 -7074 9599 -7022
rect 9651 -7074 9679 -7022
rect 9731 -7074 9759 -7022
rect 9811 -7074 9839 -7022
rect 9891 -7074 9919 -7022
rect 9971 -7074 9999 -7022
rect 10051 -7074 10079 -7022
rect 10131 -7074 10159 -7022
rect 10211 -7074 10239 -7022
rect 10291 -7074 10319 -7022
rect 10371 -7074 10399 -7022
rect 10451 -7074 10479 -7022
rect 10531 -7074 10559 -7022
rect 10611 -7074 10639 -7022
rect 10691 -7074 10719 -7022
rect 10771 -7074 10799 -7022
rect 10851 -7074 10875 -7022
rect 5745 -7088 10875 -7074
rect 4060 -7125 5610 -7115
rect 4060 -7159 4098 -7125
rect 4132 -7159 4170 -7125
rect 4204 -7159 4242 -7125
rect 4276 -7159 4314 -7125
rect 4348 -7159 4386 -7125
rect 4420 -7159 4458 -7125
rect 4492 -7159 4530 -7125
rect 4564 -7159 4602 -7125
rect 4636 -7159 4674 -7125
rect 4708 -7159 4746 -7125
rect 4780 -7159 4818 -7125
rect 4852 -7159 4890 -7125
rect 4924 -7159 4962 -7125
rect 4996 -7159 5034 -7125
rect 5068 -7159 5106 -7125
rect 5140 -7159 5178 -7125
rect 5212 -7159 5250 -7125
rect 5284 -7159 5322 -7125
rect 5356 -7159 5394 -7125
rect 5428 -7159 5466 -7125
rect 5500 -7159 5538 -7125
rect 5572 -7159 5610 -7125
rect 4060 -7167 5610 -7159
rect 4060 -7219 4094 -7167
rect 4146 -7199 4175 -7167
rect 4227 -7199 4256 -7167
rect 4308 -7199 4337 -7167
rect 4389 -7199 4418 -7167
rect 4470 -7199 4499 -7167
rect 4551 -7199 4580 -7167
rect 4632 -7199 4662 -7167
rect 4146 -7219 4170 -7199
rect 4227 -7219 4242 -7199
rect 4308 -7219 4314 -7199
rect 4492 -7219 4499 -7199
rect 4564 -7219 4580 -7199
rect 4636 -7219 4662 -7199
rect 4714 -7219 4743 -7167
rect 4795 -7199 4824 -7167
rect 4876 -7199 4905 -7167
rect 4957 -7199 4986 -7167
rect 5038 -7199 5067 -7167
rect 5119 -7199 5148 -7167
rect 5200 -7199 5230 -7167
rect 5282 -7199 5311 -7167
rect 4795 -7219 4818 -7199
rect 4876 -7219 4890 -7199
rect 4957 -7219 4962 -7199
rect 5140 -7219 5148 -7199
rect 5212 -7219 5230 -7199
rect 5284 -7219 5311 -7199
rect 5363 -7219 5392 -7167
rect 5444 -7199 5610 -7167
rect 5444 -7219 5466 -7199
rect 4060 -7233 4098 -7219
rect 4132 -7233 4170 -7219
rect 4204 -7233 4242 -7219
rect 4276 -7233 4314 -7219
rect 4348 -7233 4386 -7219
rect 4420 -7233 4458 -7219
rect 4492 -7233 4530 -7219
rect 4564 -7233 4602 -7219
rect 4636 -7233 4674 -7219
rect 4708 -7233 4746 -7219
rect 4780 -7233 4818 -7219
rect 4852 -7233 4890 -7219
rect 4924 -7233 4962 -7219
rect 4996 -7233 5034 -7219
rect 5068 -7233 5106 -7219
rect 5140 -7233 5178 -7219
rect 5212 -7233 5250 -7219
rect 5284 -7233 5322 -7219
rect 5356 -7233 5394 -7219
rect 5428 -7233 5466 -7219
rect 5500 -7233 5538 -7199
rect 5572 -7233 5610 -7199
rect 9794 -7189 10371 -7088
rect 6106 -7215 6152 -7203
rect 6106 -7223 6112 -7215
rect 6146 -7223 6152 -7215
rect 6224 -7215 6270 -7203
rect 6224 -7223 6230 -7215
rect 6264 -7223 6270 -7215
rect 6342 -7215 6388 -7203
rect 6342 -7223 6348 -7215
rect 6382 -7223 6388 -7215
rect 6460 -7215 6506 -7203
rect 6460 -7223 6466 -7215
rect 6500 -7223 6506 -7215
rect 6578 -7215 6624 -7203
rect 6578 -7223 6584 -7215
rect 6618 -7223 6624 -7215
rect 6696 -7215 6742 -7203
rect 6696 -7223 6702 -7215
rect 6736 -7223 6742 -7215
rect 6814 -7215 6860 -7203
rect 6814 -7223 6820 -7215
rect 6854 -7223 6860 -7215
rect 6932 -7215 6978 -7203
rect 6932 -7223 6938 -7215
rect 6972 -7223 6978 -7215
rect 7050 -7215 7096 -7203
rect 7050 -7223 7056 -7215
rect 7090 -7223 7096 -7215
rect 7168 -7215 7214 -7203
rect 7168 -7223 7174 -7215
rect 7208 -7223 7214 -7215
rect 7286 -7215 7332 -7203
rect 7286 -7223 7292 -7215
rect 7326 -7223 7332 -7215
rect 7404 -7215 7450 -7203
rect 7404 -7223 7410 -7215
rect 7444 -7223 7450 -7215
rect 7522 -7215 7568 -7203
rect 7522 -7223 7528 -7215
rect 7562 -7223 7568 -7215
rect 7640 -7215 7686 -7203
rect 7640 -7223 7646 -7215
rect 7680 -7223 7686 -7215
rect 7868 -7215 7914 -7203
rect 7868 -7223 7874 -7215
rect 7908 -7223 7914 -7215
rect 7986 -7215 8032 -7203
rect 7986 -7223 7992 -7215
rect 8026 -7223 8032 -7215
rect 8104 -7215 8150 -7203
rect 8104 -7223 8110 -7215
rect 8144 -7223 8150 -7215
rect 8222 -7215 8268 -7203
rect 8222 -7223 8228 -7215
rect 8262 -7223 8268 -7215
rect 8340 -7215 8386 -7203
rect 8340 -7223 8346 -7215
rect 8380 -7223 8386 -7215
rect 8458 -7215 8504 -7203
rect 8458 -7223 8464 -7215
rect 8498 -7223 8504 -7215
rect 8576 -7215 8622 -7203
rect 8576 -7223 8582 -7215
rect 8616 -7223 8622 -7215
rect 8694 -7215 8740 -7203
rect 8694 -7223 8700 -7215
rect 8734 -7223 8740 -7215
rect 8812 -7215 8858 -7203
rect 8812 -7223 8818 -7215
rect 8852 -7223 8858 -7215
rect 8930 -7215 8976 -7203
rect 8930 -7223 8936 -7215
rect 8970 -7223 8976 -7215
rect 9048 -7215 9094 -7203
rect 9048 -7223 9054 -7215
rect 9088 -7223 9094 -7215
rect 9166 -7215 9212 -7203
rect 9166 -7223 9172 -7215
rect 9206 -7223 9212 -7215
rect 9284 -7215 9330 -7203
rect 9284 -7223 9290 -7215
rect 9324 -7223 9330 -7215
rect 9402 -7215 9448 -7203
rect 9402 -7223 9408 -7215
rect 9442 -7223 9448 -7215
rect 9520 -7215 9566 -7203
rect 9520 -7223 9526 -7215
rect 9560 -7223 9566 -7215
rect 9638 -7215 9684 -7203
rect 9638 -7223 9644 -7215
rect 9678 -7223 9684 -7215
rect 9794 -7223 9834 -7189
rect 9868 -7206 9906 -7189
rect 9940 -7206 9978 -7189
rect 10012 -7206 10050 -7189
rect 10084 -7206 10122 -7189
rect 10156 -7206 10194 -7189
rect 10228 -7206 10266 -7189
rect 10300 -7206 10371 -7189
rect 9891 -7223 9906 -7206
rect 9971 -7223 9978 -7206
rect 10156 -7223 10159 -7206
rect 10228 -7223 10239 -7206
rect 10300 -7223 10319 -7206
rect 4060 -7271 5610 -7233
rect 4060 -7323 4094 -7271
rect 4146 -7273 4175 -7271
rect 4227 -7273 4256 -7271
rect 4308 -7273 4337 -7271
rect 4389 -7273 4418 -7271
rect 4470 -7273 4499 -7271
rect 4551 -7273 4580 -7271
rect 4632 -7273 4662 -7271
rect 4146 -7307 4170 -7273
rect 4227 -7307 4242 -7273
rect 4308 -7307 4314 -7273
rect 4492 -7307 4499 -7273
rect 4564 -7307 4580 -7273
rect 4636 -7307 4662 -7273
rect 4146 -7323 4175 -7307
rect 4227 -7323 4256 -7307
rect 4308 -7323 4337 -7307
rect 4389 -7323 4418 -7307
rect 4470 -7323 4499 -7307
rect 4551 -7323 4580 -7307
rect 4632 -7323 4662 -7307
rect 4714 -7323 4743 -7271
rect 4795 -7273 4824 -7271
rect 4876 -7273 4905 -7271
rect 4957 -7273 4986 -7271
rect 5038 -7273 5067 -7271
rect 5119 -7273 5148 -7271
rect 5200 -7273 5230 -7271
rect 5282 -7273 5311 -7271
rect 4795 -7307 4818 -7273
rect 4876 -7307 4890 -7273
rect 4957 -7307 4962 -7273
rect 5140 -7307 5148 -7273
rect 5212 -7307 5230 -7273
rect 5284 -7307 5311 -7273
rect 4795 -7323 4824 -7307
rect 4876 -7323 4905 -7307
rect 4957 -7323 4986 -7307
rect 5038 -7323 5067 -7307
rect 5119 -7323 5148 -7307
rect 5200 -7323 5230 -7307
rect 5282 -7323 5311 -7307
rect 5363 -7323 5392 -7271
rect 5444 -7273 5610 -7271
rect 5444 -7307 5466 -7273
rect 5500 -7307 5538 -7273
rect 5572 -7307 5610 -7273
rect 5444 -7323 5610 -7307
rect 4060 -7347 5610 -7323
rect 4060 -7375 4098 -7347
rect 4132 -7375 4170 -7347
rect 4204 -7375 4242 -7347
rect 4276 -7375 4314 -7347
rect 4348 -7375 4386 -7347
rect 4420 -7375 4458 -7347
rect 4492 -7375 4530 -7347
rect 4564 -7375 4602 -7347
rect 4636 -7375 4674 -7347
rect 4708 -7375 4746 -7347
rect 4780 -7375 4818 -7347
rect 4852 -7375 4890 -7347
rect 4924 -7375 4962 -7347
rect 4996 -7375 5034 -7347
rect 5068 -7375 5106 -7347
rect 5140 -7375 5178 -7347
rect 5212 -7375 5250 -7347
rect 5284 -7375 5322 -7347
rect 5356 -7375 5394 -7347
rect 5428 -7375 5466 -7347
rect 4060 -7427 4094 -7375
rect 4146 -7381 4170 -7375
rect 4227 -7381 4242 -7375
rect 4308 -7381 4314 -7375
rect 4492 -7381 4499 -7375
rect 4564 -7381 4580 -7375
rect 4636 -7381 4662 -7375
rect 4146 -7421 4175 -7381
rect 4227 -7421 4256 -7381
rect 4308 -7421 4337 -7381
rect 4389 -7421 4418 -7381
rect 4470 -7421 4499 -7381
rect 4551 -7421 4580 -7381
rect 4632 -7421 4662 -7381
rect 4146 -7427 4170 -7421
rect 4227 -7427 4242 -7421
rect 4308 -7427 4314 -7421
rect 4492 -7427 4499 -7421
rect 4564 -7427 4580 -7421
rect 4636 -7427 4662 -7421
rect 4714 -7427 4743 -7375
rect 4795 -7381 4818 -7375
rect 4876 -7381 4890 -7375
rect 4957 -7381 4962 -7375
rect 5140 -7381 5148 -7375
rect 5212 -7381 5230 -7375
rect 5284 -7381 5311 -7375
rect 4795 -7421 4824 -7381
rect 4876 -7421 4905 -7381
rect 4957 -7421 4986 -7381
rect 5038 -7421 5067 -7381
rect 5119 -7421 5148 -7381
rect 5200 -7421 5230 -7381
rect 5282 -7421 5311 -7381
rect 4795 -7427 4818 -7421
rect 4876 -7427 4890 -7421
rect 4957 -7427 4962 -7421
rect 5140 -7427 5148 -7421
rect 5212 -7427 5230 -7421
rect 5284 -7427 5311 -7421
rect 5363 -7427 5392 -7375
rect 5444 -7381 5466 -7375
rect 5500 -7381 5538 -7347
rect 5572 -7381 5610 -7347
rect 5444 -7421 5610 -7381
rect 5444 -7427 5466 -7421
rect 4060 -7455 4098 -7427
rect 4132 -7455 4170 -7427
rect 4204 -7455 4242 -7427
rect 4276 -7455 4314 -7427
rect 4348 -7455 4386 -7427
rect 4420 -7455 4458 -7427
rect 4492 -7455 4530 -7427
rect 4564 -7455 4602 -7427
rect 4636 -7455 4674 -7427
rect 4708 -7455 4746 -7427
rect 4780 -7455 4818 -7427
rect 4852 -7455 4890 -7427
rect 4924 -7455 4962 -7427
rect 4996 -7455 5034 -7427
rect 5068 -7455 5106 -7427
rect 5140 -7455 5178 -7427
rect 5212 -7455 5250 -7427
rect 5284 -7455 5322 -7427
rect 5356 -7455 5394 -7427
rect 5428 -7455 5466 -7427
rect 5500 -7455 5538 -7421
rect 5572 -7455 5610 -7421
rect 4060 -7479 5610 -7455
rect 4060 -7531 4094 -7479
rect 4146 -7495 4175 -7479
rect 4227 -7495 4256 -7479
rect 4308 -7495 4337 -7479
rect 4389 -7495 4418 -7479
rect 4470 -7495 4499 -7479
rect 4551 -7495 4580 -7479
rect 4632 -7495 4662 -7479
rect 4146 -7529 4170 -7495
rect 4227 -7529 4242 -7495
rect 4308 -7529 4314 -7495
rect 4492 -7529 4499 -7495
rect 4564 -7529 4580 -7495
rect 4636 -7529 4662 -7495
rect 4146 -7531 4175 -7529
rect 4227 -7531 4256 -7529
rect 4308 -7531 4337 -7529
rect 4389 -7531 4418 -7529
rect 4470 -7531 4499 -7529
rect 4551 -7531 4580 -7529
rect 4632 -7531 4662 -7529
rect 4714 -7531 4743 -7479
rect 4795 -7495 4824 -7479
rect 4876 -7495 4905 -7479
rect 4957 -7495 4986 -7479
rect 5038 -7495 5067 -7479
rect 5119 -7495 5148 -7479
rect 5200 -7495 5230 -7479
rect 5282 -7495 5311 -7479
rect 4795 -7529 4818 -7495
rect 4876 -7529 4890 -7495
rect 4957 -7529 4962 -7495
rect 5140 -7529 5148 -7495
rect 5212 -7529 5230 -7495
rect 5284 -7529 5311 -7495
rect 4795 -7531 4824 -7529
rect 4876 -7531 4905 -7529
rect 4957 -7531 4986 -7529
rect 5038 -7531 5067 -7529
rect 5119 -7531 5148 -7529
rect 5200 -7531 5230 -7529
rect 5282 -7531 5311 -7529
rect 5363 -7531 5392 -7479
rect 5444 -7495 5610 -7479
rect 5444 -7529 5466 -7495
rect 5500 -7529 5538 -7495
rect 5572 -7529 5610 -7495
rect 5444 -7531 5610 -7529
rect 4060 -7569 5610 -7531
rect 4060 -7583 4098 -7569
rect 4132 -7583 4170 -7569
rect 4204 -7583 4242 -7569
rect 4276 -7583 4314 -7569
rect 4348 -7583 4386 -7569
rect 4420 -7583 4458 -7569
rect 4492 -7583 4530 -7569
rect 4564 -7583 4602 -7569
rect 4636 -7583 4674 -7569
rect 4708 -7583 4746 -7569
rect 4780 -7583 4818 -7569
rect 4852 -7583 4890 -7569
rect 4924 -7583 4962 -7569
rect 4996 -7583 5034 -7569
rect 5068 -7583 5106 -7569
rect 5140 -7583 5178 -7569
rect 5212 -7583 5250 -7569
rect 5284 -7583 5322 -7569
rect 5356 -7583 5394 -7569
rect 5428 -7583 5466 -7569
rect 4060 -7635 4094 -7583
rect 4146 -7603 4170 -7583
rect 4227 -7603 4242 -7583
rect 4308 -7603 4314 -7583
rect 4492 -7603 4499 -7583
rect 4564 -7603 4580 -7583
rect 4636 -7603 4662 -7583
rect 4146 -7635 4175 -7603
rect 4227 -7635 4256 -7603
rect 4308 -7635 4337 -7603
rect 4389 -7635 4418 -7603
rect 4470 -7635 4499 -7603
rect 4551 -7635 4580 -7603
rect 4632 -7635 4662 -7603
rect 4714 -7635 4743 -7583
rect 4795 -7603 4818 -7583
rect 4876 -7603 4890 -7583
rect 4957 -7603 4962 -7583
rect 5140 -7603 5148 -7583
rect 5212 -7603 5230 -7583
rect 5284 -7603 5311 -7583
rect 4795 -7635 4824 -7603
rect 4876 -7635 4905 -7603
rect 4957 -7635 4986 -7603
rect 5038 -7635 5067 -7603
rect 5119 -7635 5148 -7603
rect 5200 -7635 5230 -7603
rect 5282 -7635 5311 -7603
rect 5363 -7635 5392 -7583
rect 5444 -7603 5466 -7583
rect 5500 -7603 5538 -7569
rect 5572 -7603 5610 -7569
rect 5444 -7635 5610 -7603
rect 4060 -7643 5610 -7635
rect 4060 -7677 4098 -7643
rect 4132 -7677 4170 -7643
rect 4204 -7677 4242 -7643
rect 4276 -7677 4314 -7643
rect 4348 -7677 4386 -7643
rect 4420 -7677 4458 -7643
rect 4492 -7677 4530 -7643
rect 4564 -7677 4602 -7643
rect 4636 -7677 4674 -7643
rect 4708 -7677 4746 -7643
rect 4780 -7677 4818 -7643
rect 4852 -7677 4890 -7643
rect 4924 -7677 4962 -7643
rect 4996 -7677 5034 -7643
rect 5068 -7677 5106 -7643
rect 5140 -7677 5178 -7643
rect 5212 -7677 5250 -7643
rect 5284 -7677 5322 -7643
rect 5356 -7677 5394 -7643
rect 5428 -7677 5466 -7643
rect 5500 -7677 5538 -7643
rect 5572 -7677 5610 -7643
rect 4060 -7687 5610 -7677
rect 4060 -7739 4094 -7687
rect 4146 -7717 4175 -7687
rect 4227 -7717 4256 -7687
rect 4308 -7717 4337 -7687
rect 4389 -7717 4418 -7687
rect 4470 -7717 4499 -7687
rect 4551 -7717 4580 -7687
rect 4632 -7717 4662 -7687
rect 4146 -7739 4170 -7717
rect 4227 -7739 4242 -7717
rect 4308 -7739 4314 -7717
rect 4492 -7739 4499 -7717
rect 4564 -7739 4580 -7717
rect 4636 -7739 4662 -7717
rect 4714 -7739 4743 -7687
rect 4795 -7717 4824 -7687
rect 4876 -7717 4905 -7687
rect 4957 -7717 4986 -7687
rect 5038 -7717 5067 -7687
rect 5119 -7717 5148 -7687
rect 5200 -7717 5230 -7687
rect 5282 -7717 5311 -7687
rect 4795 -7739 4818 -7717
rect 4876 -7739 4890 -7717
rect 4957 -7739 4962 -7717
rect 5140 -7739 5148 -7717
rect 5212 -7739 5230 -7717
rect 5284 -7739 5311 -7717
rect 5363 -7739 5392 -7687
rect 5444 -7717 5610 -7687
rect 5444 -7739 5466 -7717
rect 4060 -7751 4098 -7739
rect 4132 -7751 4170 -7739
rect 4204 -7751 4242 -7739
rect 4276 -7751 4314 -7739
rect 4348 -7751 4386 -7739
rect 4420 -7751 4458 -7739
rect 4492 -7751 4530 -7739
rect 4564 -7751 4602 -7739
rect 4636 -7751 4674 -7739
rect 4708 -7751 4746 -7739
rect 4780 -7751 4818 -7739
rect 4852 -7751 4890 -7739
rect 4924 -7751 4962 -7739
rect 4996 -7751 5034 -7739
rect 5068 -7751 5106 -7739
rect 5140 -7751 5178 -7739
rect 5212 -7751 5250 -7739
rect 5284 -7751 5322 -7739
rect 5356 -7751 5394 -7739
rect 5428 -7751 5466 -7739
rect 5500 -7751 5538 -7717
rect 5572 -7751 5610 -7717
rect 4060 -7791 5610 -7751
rect 5857 -7783 5867 -7223
rect 5919 -7783 5929 -7223
rect 5975 -7783 5985 -7223
rect 6037 -7783 6047 -7223
rect 6093 -7783 6103 -7223
rect 6155 -7783 6165 -7223
rect 6211 -7783 6221 -7223
rect 6273 -7783 6283 -7223
rect 6329 -7783 6339 -7223
rect 6391 -7783 6401 -7223
rect 6447 -7783 6457 -7223
rect 6509 -7783 6519 -7223
rect 6565 -7783 6575 -7223
rect 6627 -7783 6637 -7223
rect 6683 -7783 6693 -7223
rect 6745 -7783 6755 -7223
rect 6801 -7783 6811 -7223
rect 6863 -7783 6873 -7223
rect 6919 -7783 6929 -7223
rect 6981 -7783 6991 -7223
rect 7037 -7783 7047 -7223
rect 7099 -7783 7109 -7223
rect 7155 -7783 7165 -7223
rect 7217 -7783 7227 -7223
rect 7273 -7783 7283 -7223
rect 7335 -7783 7345 -7223
rect 7391 -7783 7401 -7223
rect 7453 -7783 7463 -7223
rect 7509 -7783 7519 -7223
rect 7571 -7783 7581 -7223
rect 7627 -7783 7637 -7223
rect 7689 -7783 7699 -7223
rect 7855 -7783 7865 -7223
rect 7917 -7783 7927 -7223
rect 7973 -7783 7983 -7223
rect 8035 -7783 8045 -7223
rect 8091 -7783 8101 -7223
rect 8153 -7783 8163 -7223
rect 8209 -7783 8219 -7223
rect 8271 -7783 8281 -7223
rect 8327 -7783 8337 -7223
rect 8389 -7783 8399 -7223
rect 8445 -7783 8455 -7223
rect 8507 -7783 8517 -7223
rect 8563 -7783 8573 -7223
rect 8625 -7783 8635 -7223
rect 8681 -7783 8691 -7223
rect 8743 -7783 8753 -7223
rect 8799 -7783 8809 -7223
rect 8861 -7783 8871 -7223
rect 8917 -7783 8927 -7223
rect 8979 -7783 8989 -7223
rect 9035 -7783 9045 -7223
rect 9097 -7783 9107 -7223
rect 9153 -7783 9163 -7223
rect 9215 -7783 9225 -7223
rect 9271 -7783 9281 -7223
rect 9333 -7783 9343 -7223
rect 9389 -7783 9399 -7223
rect 9451 -7783 9461 -7223
rect 9507 -7783 9517 -7223
rect 9569 -7783 9579 -7223
rect 9625 -7783 9635 -7223
rect 9687 -7783 9697 -7223
rect 9794 -7246 9839 -7223
rect 9796 -7258 9839 -7246
rect 9891 -7258 9919 -7223
rect 9971 -7258 9999 -7223
rect 10051 -7258 10079 -7223
rect 10131 -7258 10159 -7223
rect 10211 -7258 10239 -7223
rect 10291 -7258 10319 -7223
rect 9796 -7263 10371 -7258
rect 9796 -7297 9834 -7263
rect 9868 -7285 9906 -7263
rect 9940 -7285 9978 -7263
rect 10012 -7285 10050 -7263
rect 10084 -7285 10122 -7263
rect 10156 -7285 10194 -7263
rect 10228 -7285 10266 -7263
rect 10300 -7285 10371 -7263
rect 9891 -7297 9906 -7285
rect 9971 -7297 9978 -7285
rect 10156 -7297 10159 -7285
rect 10228 -7297 10239 -7285
rect 10300 -7297 10319 -7285
rect 9796 -7337 9839 -7297
rect 9891 -7337 9919 -7297
rect 9971 -7337 9999 -7297
rect 10051 -7337 10079 -7297
rect 10131 -7337 10159 -7297
rect 10211 -7337 10239 -7297
rect 10291 -7337 10319 -7297
rect 9796 -7371 9834 -7337
rect 9868 -7354 9906 -7337
rect 9940 -7354 9978 -7337
rect 10012 -7354 10050 -7337
rect 10084 -7354 10122 -7337
rect 10156 -7354 10194 -7337
rect 10228 -7354 10266 -7337
rect 10300 -7354 10371 -7337
rect 9891 -7371 9906 -7354
rect 9971 -7371 9978 -7354
rect 10156 -7371 10159 -7354
rect 10228 -7371 10239 -7354
rect 10300 -7371 10319 -7354
rect 9796 -7406 9839 -7371
rect 9891 -7406 9919 -7371
rect 9971 -7406 9999 -7371
rect 10051 -7406 10079 -7371
rect 10131 -7406 10159 -7371
rect 10211 -7406 10239 -7371
rect 10291 -7406 10319 -7371
rect 9796 -7411 10371 -7406
rect 9796 -7445 9834 -7411
rect 9868 -7433 9906 -7411
rect 9940 -7433 9978 -7411
rect 10012 -7433 10050 -7411
rect 10084 -7433 10122 -7411
rect 10156 -7433 10194 -7411
rect 10228 -7433 10266 -7411
rect 10300 -7433 10371 -7411
rect 9891 -7445 9906 -7433
rect 9971 -7445 9978 -7433
rect 10156 -7445 10159 -7433
rect 10228 -7445 10239 -7433
rect 10300 -7445 10319 -7433
rect 9796 -7485 9839 -7445
rect 9891 -7485 9919 -7445
rect 9971 -7485 9999 -7445
rect 10051 -7485 10079 -7445
rect 10131 -7485 10159 -7445
rect 10211 -7485 10239 -7445
rect 10291 -7485 10319 -7445
rect 9796 -7519 9834 -7485
rect 9868 -7519 9906 -7485
rect 9940 -7519 9978 -7485
rect 10012 -7519 10050 -7485
rect 10084 -7519 10122 -7485
rect 10156 -7519 10194 -7485
rect 10228 -7519 10266 -7485
rect 10300 -7519 10371 -7485
rect 9796 -7559 10371 -7519
rect 9796 -7593 9834 -7559
rect 9868 -7593 9906 -7559
rect 9940 -7593 9978 -7559
rect 10012 -7593 10050 -7559
rect 10084 -7593 10122 -7559
rect 10156 -7593 10194 -7559
rect 10228 -7593 10266 -7559
rect 10300 -7582 10371 -7559
rect 10415 -7191 10461 -7179
rect 10415 -7225 10421 -7191
rect 10455 -7225 10461 -7191
rect 10415 -7264 10461 -7225
rect 10415 -7298 10421 -7264
rect 10455 -7298 10461 -7264
rect 10415 -7337 10461 -7298
rect 10415 -7371 10421 -7337
rect 10455 -7371 10461 -7337
rect 10415 -7410 10461 -7371
rect 10731 -7191 10777 -7179
rect 10731 -7225 10737 -7191
rect 10771 -7225 10777 -7191
rect 10731 -7264 10777 -7225
rect 10731 -7298 10737 -7264
rect 10771 -7298 10777 -7264
rect 10731 -7337 10777 -7298
rect 10731 -7371 10737 -7337
rect 10771 -7371 10777 -7337
rect 11047 -7191 11093 -7179
rect 11047 -7225 11053 -7191
rect 11087 -7225 11093 -7191
rect 11047 -7264 11093 -7225
rect 11047 -7298 11053 -7264
rect 11087 -7298 11093 -7264
rect 11047 -7337 11093 -7298
rect 10415 -7444 10421 -7410
rect 10455 -7444 10461 -7410
rect 10415 -7483 10461 -7444
rect 10415 -7517 10421 -7483
rect 10455 -7517 10461 -7483
rect 10503 -7515 10513 -7395
rect 10565 -7515 10575 -7395
rect 10617 -7515 10627 -7395
rect 10679 -7515 10689 -7395
rect 10731 -7410 10777 -7371
rect 10845 -7377 10891 -7365
rect 10845 -7395 10851 -7377
rect 10731 -7444 10737 -7410
rect 10771 -7444 10777 -7410
rect 10731 -7483 10777 -7444
rect 10415 -7556 10461 -7517
rect 10300 -7593 10359 -7582
rect 9796 -7633 10359 -7593
rect 9796 -7667 9834 -7633
rect 9868 -7667 9906 -7633
rect 9940 -7667 9978 -7633
rect 10012 -7667 10050 -7633
rect 10084 -7667 10122 -7633
rect 10156 -7667 10194 -7633
rect 10228 -7667 10266 -7633
rect 10300 -7667 10359 -7633
rect 9796 -7689 10359 -7667
rect 10415 -7590 10421 -7556
rect 10455 -7590 10461 -7556
rect 10415 -7649 10461 -7590
rect 10731 -7517 10737 -7483
rect 10771 -7517 10777 -7483
rect 10819 -7515 10829 -7395
rect 10885 -7503 10891 -7377
rect 10881 -7515 10891 -7503
rect 10933 -7377 10979 -7365
rect 10933 -7503 10939 -7377
rect 10973 -7395 10979 -7377
rect 11047 -7371 11053 -7337
rect 11087 -7371 11093 -7337
rect 11363 -7191 11409 -7179
rect 11363 -7225 11369 -7191
rect 11403 -7225 11409 -7191
rect 11363 -7264 11409 -7225
rect 11363 -7298 11369 -7264
rect 11403 -7298 11409 -7264
rect 11363 -7337 11409 -7298
rect 10933 -7515 10943 -7503
rect 10995 -7515 11005 -7395
rect 11047 -7410 11093 -7371
rect 11161 -7377 11207 -7365
rect 11161 -7395 11167 -7377
rect 11047 -7444 11053 -7410
rect 11087 -7444 11093 -7410
rect 11047 -7483 11093 -7444
rect 10731 -7556 10777 -7517
rect 10731 -7590 10737 -7556
rect 10771 -7590 10777 -7556
rect 10731 -7649 10777 -7590
rect 11047 -7517 11053 -7483
rect 11087 -7517 11093 -7483
rect 11135 -7515 11145 -7395
rect 11201 -7503 11207 -7377
rect 11197 -7515 11207 -7503
rect 11249 -7377 11295 -7365
rect 11249 -7503 11255 -7377
rect 11289 -7395 11295 -7377
rect 11363 -7371 11369 -7337
rect 11403 -7371 11409 -7337
rect 11679 -7191 11725 -7179
rect 11679 -7225 11685 -7191
rect 11719 -7225 11725 -7191
rect 11679 -7264 11725 -7225
rect 11679 -7298 11685 -7264
rect 11719 -7298 11725 -7264
rect 11679 -7337 11725 -7298
rect 11249 -7515 11259 -7503
rect 11311 -7515 11321 -7395
rect 11363 -7410 11409 -7371
rect 11477 -7377 11523 -7365
rect 11477 -7395 11483 -7377
rect 11363 -7444 11369 -7410
rect 11403 -7444 11409 -7410
rect 11363 -7483 11409 -7444
rect 11047 -7556 11093 -7517
rect 11047 -7590 11053 -7556
rect 11087 -7590 11093 -7556
rect 11047 -7649 11093 -7590
rect 11363 -7517 11369 -7483
rect 11403 -7517 11409 -7483
rect 11451 -7515 11461 -7395
rect 11517 -7503 11523 -7377
rect 11513 -7515 11523 -7503
rect 11565 -7377 11611 -7365
rect 11565 -7503 11571 -7377
rect 11605 -7395 11611 -7377
rect 11679 -7371 11685 -7337
rect 11719 -7371 11725 -7337
rect 11995 -7191 12041 -7179
rect 11995 -7225 12001 -7191
rect 12035 -7225 12041 -7191
rect 11995 -7264 12041 -7225
rect 11995 -7298 12001 -7264
rect 12035 -7298 12041 -7264
rect 11995 -7337 12041 -7298
rect 11565 -7515 11575 -7503
rect 11627 -7515 11637 -7395
rect 11679 -7410 11725 -7371
rect 11793 -7377 11839 -7365
rect 11793 -7395 11799 -7377
rect 11679 -7444 11685 -7410
rect 11719 -7444 11725 -7410
rect 11679 -7483 11725 -7444
rect 11363 -7556 11409 -7517
rect 11363 -7590 11369 -7556
rect 11403 -7590 11409 -7556
rect 11363 -7649 11409 -7590
rect 11679 -7517 11685 -7483
rect 11719 -7517 11725 -7483
rect 11767 -7515 11777 -7395
rect 11833 -7503 11839 -7377
rect 11829 -7515 11839 -7503
rect 11881 -7377 11927 -7365
rect 11881 -7503 11887 -7377
rect 11921 -7395 11927 -7377
rect 11995 -7371 12001 -7337
rect 12035 -7371 12041 -7337
rect 12311 -7191 12357 -7179
rect 12311 -7225 12317 -7191
rect 12351 -7225 12357 -7191
rect 12528 -7215 12574 -7203
rect 12528 -7219 12534 -7215
rect 12568 -7219 12574 -7215
rect 12676 -7215 12722 -7203
rect 12676 -7219 12682 -7215
rect 12716 -7219 12722 -7215
rect 12824 -7215 12870 -7203
rect 12824 -7219 12830 -7215
rect 12864 -7219 12870 -7215
rect 12972 -7215 13018 -7203
rect 12972 -7219 12978 -7215
rect 13012 -7219 13018 -7215
rect 13120 -7215 13166 -7203
rect 13120 -7219 13126 -7215
rect 13160 -7219 13166 -7215
rect 13268 -7215 13314 -7203
rect 13268 -7219 13274 -7215
rect 13308 -7219 13314 -7215
rect 13416 -7215 13462 -7203
rect 13416 -7219 13422 -7215
rect 13456 -7219 13462 -7215
rect 13564 -7215 13610 -7203
rect 13564 -7219 13570 -7215
rect 13604 -7219 13610 -7215
rect 13712 -7215 13758 -7203
rect 13712 -7219 13718 -7215
rect 13752 -7219 13758 -7215
rect 13860 -7215 13906 -7203
rect 13860 -7219 13866 -7215
rect 13900 -7219 13906 -7215
rect 14008 -7215 14054 -7203
rect 14008 -7219 14014 -7215
rect 14048 -7219 14054 -7215
rect 14156 -7215 14202 -7203
rect 14156 -7219 14162 -7215
rect 14196 -7219 14202 -7215
rect 14304 -7215 14350 -7203
rect 14304 -7219 14310 -7215
rect 14344 -7219 14350 -7215
rect 14452 -7215 14498 -7203
rect 14452 -7219 14458 -7215
rect 14492 -7219 14498 -7215
rect 14600 -7215 14646 -7203
rect 14600 -7219 14606 -7215
rect 14640 -7219 14646 -7215
rect 14748 -7215 14794 -7203
rect 14748 -7219 14754 -7215
rect 14788 -7219 14794 -7215
rect 14896 -7215 14942 -7203
rect 14896 -7219 14902 -7215
rect 14936 -7219 14942 -7215
rect 15044 -7215 15090 -7203
rect 15044 -7219 15050 -7215
rect 15084 -7219 15090 -7215
rect 15192 -7215 15238 -7203
rect 15192 -7219 15198 -7215
rect 15232 -7219 15238 -7215
rect 15340 -7215 15386 -7203
rect 15340 -7219 15346 -7215
rect 15380 -7219 15386 -7215
rect 15488 -7215 15534 -7203
rect 15488 -7219 15494 -7215
rect 15528 -7219 15534 -7215
rect 15636 -7215 15682 -7203
rect 15636 -7219 15642 -7215
rect 15676 -7219 15682 -7215
rect 15784 -7215 15830 -7203
rect 15784 -7219 15790 -7215
rect 15824 -7219 15830 -7215
rect 15932 -7215 15978 -7203
rect 15932 -7219 15938 -7215
rect 15972 -7219 15978 -7215
rect 16080 -7215 16126 -7203
rect 16080 -7219 16086 -7215
rect 16120 -7219 16126 -7215
rect 16228 -7215 16274 -7203
rect 16228 -7219 16234 -7215
rect 16268 -7219 16274 -7215
rect 16376 -7215 16422 -7203
rect 16376 -7219 16382 -7215
rect 16416 -7219 16422 -7215
rect 16524 -7215 16570 -7203
rect 16524 -7219 16530 -7215
rect 16564 -7219 16570 -7215
rect 16672 -7215 16718 -7203
rect 16672 -7219 16678 -7215
rect 16712 -7219 16718 -7215
rect 16820 -7215 16866 -7203
rect 16820 -7219 16826 -7215
rect 16860 -7219 16866 -7215
rect 16968 -7215 17014 -7203
rect 16968 -7219 16974 -7215
rect 17008 -7219 17014 -7215
rect 17116 -7215 17162 -7203
rect 17116 -7219 17122 -7215
rect 17156 -7219 17162 -7215
rect 17264 -7215 17310 -7203
rect 17264 -7219 17270 -7215
rect 17304 -7219 17310 -7215
rect 17412 -7215 17458 -7203
rect 17412 -7219 17418 -7215
rect 17452 -7219 17458 -7215
rect 17560 -7215 17606 -7203
rect 17560 -7219 17566 -7215
rect 17600 -7219 17606 -7215
rect 17708 -7215 17754 -7203
rect 17708 -7219 17714 -7215
rect 17748 -7219 17754 -7215
rect 17856 -7215 17902 -7203
rect 17856 -7219 17862 -7215
rect 17896 -7219 17902 -7215
rect 18004 -7215 18050 -7203
rect 18004 -7219 18010 -7215
rect 18044 -7219 18050 -7215
rect 18152 -7215 18198 -7203
rect 18152 -7219 18158 -7215
rect 18192 -7219 18198 -7215
rect 18300 -7215 18346 -7203
rect 18300 -7219 18306 -7215
rect 18340 -7219 18346 -7215
rect 18448 -7215 18494 -7203
rect 18448 -7219 18454 -7215
rect 18488 -7219 18494 -7215
rect 18596 -7215 18642 -7203
rect 18596 -7219 18602 -7215
rect 18636 -7219 18642 -7215
rect 18744 -7215 18790 -7203
rect 18744 -7219 18750 -7215
rect 18784 -7219 18790 -7215
rect 18892 -7215 18938 -7203
rect 18892 -7219 18898 -7215
rect 18932 -7219 18938 -7215
rect 19040 -7215 19086 -7203
rect 19040 -7219 19046 -7215
rect 19080 -7219 19086 -7215
rect 19188 -7215 19234 -7203
rect 19188 -7219 19194 -7215
rect 19228 -7219 19234 -7215
rect 19336 -7215 19382 -7203
rect 19336 -7219 19342 -7215
rect 19376 -7219 19382 -7215
rect 19484 -7215 19530 -7203
rect 19484 -7219 19490 -7215
rect 19524 -7219 19530 -7215
rect 19632 -7215 19678 -7203
rect 19632 -7219 19638 -7215
rect 19672 -7219 19678 -7215
rect 19780 -7215 19826 -7203
rect 19780 -7219 19786 -7215
rect 19820 -7219 19826 -7215
rect 19928 -7215 19974 -7203
rect 19928 -7219 19934 -7215
rect 19968 -7219 19974 -7215
rect 20076 -7215 20122 -7203
rect 20076 -7219 20082 -7215
rect 20116 -7219 20122 -7215
rect 20224 -7215 20270 -7203
rect 20224 -7219 20230 -7215
rect 20264 -7219 20270 -7215
rect 20372 -7215 20418 -7203
rect 20372 -7219 20378 -7215
rect 20412 -7219 20418 -7215
rect 20520 -7215 20566 -7203
rect 20520 -7219 20526 -7215
rect 20560 -7219 20566 -7215
rect 20668 -7215 20714 -7203
rect 20668 -7219 20674 -7215
rect 20708 -7219 20714 -7215
rect 20816 -7215 20862 -7203
rect 20816 -7219 20822 -7215
rect 20856 -7219 20862 -7215
rect 20964 -7215 21010 -7203
rect 20964 -7219 20970 -7215
rect 21004 -7219 21010 -7215
rect 21112 -7215 21158 -7203
rect 21112 -7219 21118 -7215
rect 21152 -7219 21158 -7215
rect 21260 -7215 21306 -7203
rect 21260 -7219 21266 -7215
rect 21300 -7219 21306 -7215
rect 21408 -7215 21454 -7203
rect 21408 -7219 21414 -7215
rect 21448 -7219 21454 -7215
rect 21556 -7215 21602 -7203
rect 21556 -7219 21562 -7215
rect 21596 -7219 21602 -7215
rect 21704 -7215 21750 -7203
rect 21704 -7219 21710 -7215
rect 21744 -7219 21750 -7215
rect 21852 -7215 21898 -7203
rect 21852 -7219 21858 -7215
rect 21892 -7219 21898 -7215
rect 22000 -7215 22046 -7203
rect 22000 -7219 22006 -7215
rect 22040 -7219 22046 -7215
rect 22148 -7215 22194 -7203
rect 22148 -7219 22154 -7215
rect 22188 -7219 22194 -7215
rect 22296 -7215 22342 -7203
rect 22296 -7219 22302 -7215
rect 22336 -7219 22342 -7215
rect 22444 -7215 22490 -7203
rect 22444 -7219 22450 -7215
rect 22484 -7219 22490 -7215
rect 22592 -7215 22638 -7203
rect 22592 -7219 22598 -7215
rect 22632 -7219 22638 -7215
rect 22740 -7215 22786 -7203
rect 22740 -7219 22746 -7215
rect 22780 -7219 22786 -7215
rect 22888 -7215 22934 -7203
rect 22888 -7219 22894 -7215
rect 22928 -7219 22934 -7215
rect 23036 -7215 23082 -7203
rect 23036 -7219 23042 -7215
rect 23076 -7219 23082 -7215
rect 23184 -7215 23230 -7203
rect 23184 -7219 23190 -7215
rect 23224 -7219 23230 -7215
rect 23332 -7215 23378 -7203
rect 23332 -7219 23338 -7215
rect 23372 -7219 23378 -7215
rect 23628 -7215 23674 -7203
rect 23628 -7219 23634 -7215
rect 23668 -7219 23674 -7215
rect 12311 -7264 12357 -7225
rect 12311 -7298 12317 -7264
rect 12351 -7298 12357 -7264
rect 12311 -7337 12357 -7298
rect 11881 -7515 11891 -7503
rect 11943 -7515 11953 -7395
rect 11995 -7410 12041 -7371
rect 12109 -7377 12155 -7365
rect 12109 -7395 12115 -7377
rect 11995 -7444 12001 -7410
rect 12035 -7444 12041 -7410
rect 11995 -7483 12041 -7444
rect 11679 -7556 11725 -7517
rect 11679 -7590 11685 -7556
rect 11719 -7590 11725 -7556
rect 11679 -7649 11725 -7590
rect 11995 -7517 12001 -7483
rect 12035 -7517 12041 -7483
rect 12083 -7515 12093 -7395
rect 12149 -7503 12155 -7377
rect 12145 -7515 12155 -7503
rect 12197 -7377 12243 -7365
rect 12197 -7503 12203 -7377
rect 12237 -7395 12243 -7377
rect 12311 -7371 12317 -7337
rect 12351 -7371 12357 -7337
rect 12197 -7515 12207 -7503
rect 12259 -7515 12269 -7395
rect 12311 -7410 12357 -7371
rect 12311 -7444 12317 -7410
rect 12351 -7444 12357 -7410
rect 12311 -7483 12357 -7444
rect 11995 -7556 12041 -7517
rect 11995 -7590 12001 -7556
rect 12035 -7590 12041 -7556
rect 11995 -7649 12041 -7590
rect 12311 -7517 12317 -7483
rect 12351 -7517 12357 -7483
rect 12311 -7556 12357 -7517
rect 12311 -7590 12317 -7556
rect 12351 -7590 12357 -7556
rect 12311 -7649 12357 -7590
rect 10415 -7655 12365 -7649
rect 10415 -7689 10421 -7655
rect 10455 -7689 10494 -7655
rect 10528 -7689 10567 -7655
rect 10601 -7689 10640 -7655
rect 10674 -7689 10713 -7655
rect 10747 -7689 10786 -7655
rect 10820 -7689 10859 -7655
rect 10893 -7689 10932 -7655
rect 10966 -7689 11005 -7655
rect 11039 -7689 11078 -7655
rect 11112 -7689 11151 -7655
rect 11185 -7689 11224 -7655
rect 11258 -7689 11297 -7655
rect 11331 -7689 11370 -7655
rect 11404 -7689 11443 -7655
rect 11477 -7689 11516 -7655
rect 11550 -7689 11589 -7655
rect 11623 -7689 11662 -7655
rect 11696 -7689 11735 -7655
rect 11769 -7689 11808 -7655
rect 11842 -7689 11881 -7655
rect 11915 -7689 11954 -7655
rect 11988 -7689 12027 -7655
rect 12061 -7689 12100 -7655
rect 12134 -7689 12173 -7655
rect 12207 -7689 12246 -7655
rect 12280 -7689 12319 -7655
rect 12353 -7689 12365 -7655
rect 9796 -7695 12365 -7689
rect 9796 -7707 12342 -7695
rect 9796 -7741 9834 -7707
rect 9868 -7741 9906 -7707
rect 9940 -7741 9978 -7707
rect 10012 -7741 10050 -7707
rect 10084 -7741 10122 -7707
rect 10156 -7741 10194 -7707
rect 10228 -7741 10266 -7707
rect 10300 -7741 12342 -7707
rect 9796 -7781 12342 -7741
rect 4060 -7843 4094 -7791
rect 4146 -7825 4170 -7791
rect 4227 -7825 4242 -7791
rect 4308 -7825 4314 -7791
rect 4492 -7825 4499 -7791
rect 4564 -7825 4580 -7791
rect 4636 -7825 4662 -7791
rect 4146 -7843 4175 -7825
rect 4227 -7843 4256 -7825
rect 4308 -7843 4337 -7825
rect 4389 -7843 4418 -7825
rect 4470 -7843 4499 -7825
rect 4551 -7843 4580 -7825
rect 4632 -7843 4662 -7825
rect 4714 -7843 4743 -7791
rect 4795 -7825 4818 -7791
rect 4876 -7825 4890 -7791
rect 4957 -7825 4962 -7791
rect 5140 -7825 5148 -7791
rect 5212 -7825 5230 -7791
rect 5284 -7825 5311 -7791
rect 4795 -7843 4824 -7825
rect 4876 -7843 4905 -7825
rect 4957 -7843 4986 -7825
rect 5038 -7843 5067 -7825
rect 5119 -7843 5148 -7825
rect 5200 -7843 5230 -7825
rect 5282 -7843 5311 -7825
rect 5363 -7843 5392 -7791
rect 5444 -7825 5466 -7791
rect 5500 -7825 5538 -7791
rect 5572 -7825 5610 -7791
rect 6106 -7791 6112 -7783
rect 6146 -7791 6152 -7783
rect 6106 -7803 6152 -7791
rect 6224 -7791 6230 -7783
rect 6264 -7791 6270 -7783
rect 6224 -7803 6270 -7791
rect 6342 -7791 6348 -7783
rect 6382 -7791 6388 -7783
rect 6342 -7803 6388 -7791
rect 6460 -7791 6466 -7783
rect 6500 -7791 6506 -7783
rect 6460 -7803 6506 -7791
rect 6578 -7791 6584 -7783
rect 6618 -7791 6624 -7783
rect 6578 -7803 6624 -7791
rect 6696 -7791 6702 -7783
rect 6736 -7791 6742 -7783
rect 6696 -7803 6742 -7791
rect 6814 -7791 6820 -7783
rect 6854 -7791 6860 -7783
rect 6814 -7803 6860 -7791
rect 6932 -7791 6938 -7783
rect 6972 -7791 6978 -7783
rect 6932 -7803 6978 -7791
rect 7050 -7791 7056 -7783
rect 7090 -7791 7096 -7783
rect 7050 -7803 7096 -7791
rect 7168 -7791 7174 -7783
rect 7208 -7791 7214 -7783
rect 7168 -7803 7214 -7791
rect 7286 -7791 7292 -7783
rect 7326 -7791 7332 -7783
rect 7286 -7803 7332 -7791
rect 7404 -7791 7410 -7783
rect 7444 -7791 7450 -7783
rect 7404 -7803 7450 -7791
rect 7522 -7791 7528 -7783
rect 7562 -7791 7568 -7783
rect 7522 -7803 7568 -7791
rect 7640 -7791 7646 -7783
rect 7680 -7791 7686 -7783
rect 7640 -7803 7686 -7791
rect 7868 -7791 7874 -7783
rect 7908 -7791 7914 -7783
rect 7868 -7803 7914 -7791
rect 7986 -7791 7992 -7783
rect 8026 -7791 8032 -7783
rect 7986 -7803 8032 -7791
rect 8104 -7791 8110 -7783
rect 8144 -7791 8150 -7783
rect 8104 -7803 8150 -7791
rect 8222 -7791 8228 -7783
rect 8262 -7791 8268 -7783
rect 8222 -7803 8268 -7791
rect 8340 -7791 8346 -7783
rect 8380 -7791 8386 -7783
rect 8340 -7803 8386 -7791
rect 8458 -7791 8464 -7783
rect 8498 -7791 8504 -7783
rect 8458 -7803 8504 -7791
rect 8576 -7791 8582 -7783
rect 8616 -7791 8622 -7783
rect 8576 -7803 8622 -7791
rect 8694 -7791 8700 -7783
rect 8734 -7791 8740 -7783
rect 8694 -7803 8740 -7791
rect 8812 -7791 8818 -7783
rect 8852 -7791 8858 -7783
rect 8812 -7803 8858 -7791
rect 8930 -7791 8936 -7783
rect 8970 -7791 8976 -7783
rect 8930 -7803 8976 -7791
rect 9048 -7791 9054 -7783
rect 9088 -7791 9094 -7783
rect 9048 -7803 9094 -7791
rect 9166 -7791 9172 -7783
rect 9206 -7791 9212 -7783
rect 9166 -7803 9212 -7791
rect 9284 -7791 9290 -7783
rect 9324 -7791 9330 -7783
rect 9284 -7803 9330 -7791
rect 9402 -7791 9408 -7783
rect 9442 -7791 9448 -7783
rect 9402 -7803 9448 -7791
rect 9520 -7791 9526 -7783
rect 9560 -7791 9566 -7783
rect 9520 -7803 9566 -7791
rect 9638 -7791 9644 -7783
rect 9678 -7791 9684 -7783
rect 9638 -7803 9684 -7791
rect 5444 -7843 5610 -7825
rect 9796 -7815 9834 -7781
rect 9868 -7815 9906 -7781
rect 9940 -7815 9978 -7781
rect 10012 -7815 10050 -7781
rect 10084 -7815 10122 -7781
rect 10156 -7815 10194 -7781
rect 10228 -7815 10266 -7781
rect 10300 -7815 10338 -7781
rect 10372 -7815 10410 -7781
rect 10444 -7815 10482 -7781
rect 10516 -7815 10554 -7781
rect 10588 -7815 12342 -7781
rect 4060 -7865 5610 -7843
rect 4060 -7895 4098 -7865
rect 4132 -7895 4170 -7865
rect 4204 -7895 4242 -7865
rect 4276 -7895 4314 -7865
rect 4348 -7895 4386 -7865
rect 4420 -7895 4458 -7865
rect 4492 -7895 4530 -7865
rect 4564 -7895 4602 -7865
rect 4636 -7895 4674 -7865
rect 4708 -7895 4746 -7865
rect 4780 -7895 4818 -7865
rect 4852 -7895 4890 -7865
rect 4924 -7895 4962 -7865
rect 4996 -7895 5034 -7865
rect 5068 -7895 5106 -7865
rect 5140 -7895 5178 -7865
rect 5212 -7895 5250 -7865
rect 5284 -7895 5322 -7865
rect 5356 -7895 5394 -7865
rect 5428 -7895 5466 -7865
rect 4060 -7947 4094 -7895
rect 4146 -7899 4170 -7895
rect 4227 -7899 4242 -7895
rect 4308 -7899 4314 -7895
rect 4492 -7899 4499 -7895
rect 4564 -7899 4580 -7895
rect 4636 -7899 4662 -7895
rect 4146 -7939 4175 -7899
rect 4227 -7939 4256 -7899
rect 4308 -7939 4337 -7899
rect 4389 -7939 4418 -7899
rect 4470 -7939 4499 -7899
rect 4551 -7939 4580 -7899
rect 4632 -7939 4662 -7899
rect 4146 -7947 4170 -7939
rect 4227 -7947 4242 -7939
rect 4308 -7947 4314 -7939
rect 4492 -7947 4499 -7939
rect 4564 -7947 4580 -7939
rect 4636 -7947 4662 -7939
rect 4714 -7947 4743 -7895
rect 4795 -7899 4818 -7895
rect 4876 -7899 4890 -7895
rect 4957 -7899 4962 -7895
rect 5140 -7899 5148 -7895
rect 5212 -7899 5230 -7895
rect 5284 -7899 5311 -7895
rect 4795 -7939 4824 -7899
rect 4876 -7939 4905 -7899
rect 4957 -7939 4986 -7899
rect 5038 -7939 5067 -7899
rect 5119 -7939 5148 -7899
rect 5200 -7939 5230 -7899
rect 5282 -7939 5311 -7899
rect 4795 -7947 4818 -7939
rect 4876 -7947 4890 -7939
rect 4957 -7947 4962 -7939
rect 5140 -7947 5148 -7939
rect 5212 -7947 5230 -7939
rect 5284 -7947 5311 -7939
rect 5363 -7947 5392 -7895
rect 5444 -7899 5466 -7895
rect 5500 -7899 5538 -7865
rect 5572 -7899 5610 -7865
rect 5444 -7939 5610 -7899
rect 5444 -7947 5466 -7939
rect 4060 -7973 4098 -7947
rect 4132 -7973 4170 -7947
rect 4204 -7973 4242 -7947
rect 4276 -7973 4314 -7947
rect 4348 -7973 4386 -7947
rect 4420 -7973 4458 -7947
rect 4492 -7973 4530 -7947
rect 4564 -7973 4602 -7947
rect 4636 -7973 4674 -7947
rect 4708 -7973 4746 -7947
rect 4780 -7973 4818 -7947
rect 4852 -7973 4890 -7947
rect 4924 -7973 4962 -7947
rect 4996 -7973 5034 -7947
rect 5068 -7973 5106 -7947
rect 5140 -7973 5178 -7947
rect 5212 -7973 5250 -7947
rect 5284 -7973 5322 -7947
rect 5356 -7973 5394 -7947
rect 5428 -7973 5466 -7947
rect 5500 -7973 5538 -7939
rect 5572 -7973 5610 -7939
rect 4060 -7999 5610 -7973
rect 5913 -7989 5923 -7835
rect 5981 -7989 5991 -7835
rect 6031 -7989 6041 -7835
rect 6099 -7989 6109 -7835
rect 6149 -7989 6159 -7835
rect 6217 -7989 6227 -7835
rect 6267 -7989 6277 -7835
rect 6335 -7989 6345 -7835
rect 6385 -7989 6395 -7835
rect 6453 -7989 6463 -7835
rect 6503 -7989 6513 -7835
rect 6571 -7989 6581 -7835
rect 6621 -7989 6631 -7835
rect 6689 -7989 6699 -7835
rect 6739 -7989 6749 -7835
rect 6807 -7989 6817 -7835
rect 6857 -7989 6867 -7835
rect 6925 -7989 6935 -7835
rect 6975 -7989 6985 -7835
rect 7043 -7989 7053 -7835
rect 7093 -7989 7103 -7835
rect 7161 -7989 7171 -7835
rect 7211 -7989 7221 -7835
rect 7279 -7989 7289 -7835
rect 7329 -7989 7339 -7835
rect 7397 -7989 7407 -7835
rect 7447 -7989 7457 -7835
rect 7515 -7989 7525 -7835
rect 7565 -7989 7575 -7835
rect 7633 -7989 7643 -7835
rect 7911 -7989 7921 -7835
rect 7979 -7989 7989 -7835
rect 8029 -7989 8039 -7835
rect 8097 -7989 8107 -7835
rect 8147 -7989 8157 -7835
rect 8215 -7989 8225 -7835
rect 8265 -7989 8275 -7835
rect 8333 -7989 8343 -7835
rect 8383 -7989 8393 -7835
rect 8451 -7989 8461 -7835
rect 8501 -7989 8511 -7835
rect 8569 -7989 8579 -7835
rect 8619 -7989 8629 -7835
rect 8687 -7989 8697 -7835
rect 8737 -7989 8747 -7835
rect 8805 -7989 8815 -7835
rect 8855 -7989 8865 -7835
rect 8923 -7989 8933 -7835
rect 8973 -7989 8983 -7835
rect 9041 -7989 9051 -7835
rect 9091 -7989 9101 -7835
rect 9159 -7989 9169 -7835
rect 9209 -7989 9219 -7835
rect 9277 -7989 9287 -7835
rect 9327 -7989 9337 -7835
rect 9395 -7989 9405 -7835
rect 9445 -7989 9455 -7835
rect 9513 -7989 9523 -7835
rect 9563 -7989 9573 -7835
rect 9631 -7989 9641 -7835
rect 9796 -7855 12342 -7815
rect 9796 -7889 9834 -7855
rect 9868 -7889 9906 -7855
rect 9940 -7889 9978 -7855
rect 10012 -7889 10050 -7855
rect 10084 -7889 10122 -7855
rect 10156 -7889 10194 -7855
rect 10228 -7889 10266 -7855
rect 10300 -7889 10338 -7855
rect 10372 -7889 10410 -7855
rect 10444 -7889 10482 -7855
rect 10516 -7889 10554 -7855
rect 10588 -7889 12342 -7855
rect 9796 -7905 12342 -7889
rect 9796 -7929 10482 -7905
rect 9796 -7963 9834 -7929
rect 9868 -7963 9906 -7929
rect 9940 -7963 9978 -7929
rect 10012 -7963 10050 -7929
rect 10084 -7963 10122 -7929
rect 10156 -7963 10194 -7929
rect 10228 -7963 10266 -7929
rect 10300 -7963 10338 -7929
rect 10372 -7963 10410 -7929
rect 10444 -7963 10482 -7929
rect 4060 -8051 4094 -7999
rect 4146 -8013 4175 -7999
rect 4227 -8013 4256 -7999
rect 4308 -8013 4337 -7999
rect 4389 -8013 4418 -7999
rect 4470 -8013 4499 -7999
rect 4551 -8013 4580 -7999
rect 4632 -8013 4662 -7999
rect 4146 -8047 4170 -8013
rect 4227 -8047 4242 -8013
rect 4308 -8047 4314 -8013
rect 4492 -8047 4499 -8013
rect 4564 -8047 4580 -8013
rect 4636 -8047 4662 -8013
rect 4146 -8051 4175 -8047
rect 4227 -8051 4256 -8047
rect 4308 -8051 4337 -8047
rect 4389 -8051 4418 -8047
rect 4470 -8051 4499 -8047
rect 4551 -8051 4580 -8047
rect 4632 -8051 4662 -8047
rect 4714 -8051 4743 -7999
rect 4795 -8013 4824 -7999
rect 4876 -8013 4905 -7999
rect 4957 -8013 4986 -7999
rect 5038 -8013 5067 -7999
rect 5119 -8013 5148 -7999
rect 5200 -8013 5230 -7999
rect 5282 -8013 5311 -7999
rect 4795 -8047 4818 -8013
rect 4876 -8047 4890 -8013
rect 4957 -8047 4962 -8013
rect 5140 -8047 5148 -8013
rect 5212 -8047 5230 -8013
rect 5284 -8047 5311 -8013
rect 4795 -8051 4824 -8047
rect 4876 -8051 4905 -8047
rect 4957 -8051 4986 -8047
rect 5038 -8051 5067 -8047
rect 5119 -8051 5148 -8047
rect 5200 -8051 5230 -8047
rect 5282 -8051 5311 -8047
rect 5363 -8051 5392 -7999
rect 5444 -8013 5610 -7999
rect 5444 -8047 5466 -8013
rect 5500 -8047 5538 -8013
rect 5572 -8047 5610 -8013
rect 9796 -8003 10482 -7963
rect 5870 -8033 5916 -8021
rect 5870 -8041 5876 -8033
rect 5910 -8041 5916 -8033
rect 5988 -8033 6034 -8021
rect 5988 -8041 5994 -8033
rect 6028 -8041 6034 -8033
rect 6106 -8033 6152 -8021
rect 6106 -8041 6112 -8033
rect 6146 -8041 6152 -8033
rect 6224 -8033 6270 -8021
rect 6224 -8041 6230 -8033
rect 6264 -8041 6270 -8033
rect 6342 -8033 6388 -8021
rect 6342 -8041 6348 -8033
rect 6382 -8041 6388 -8033
rect 6460 -8033 6506 -8021
rect 6460 -8041 6466 -8033
rect 6500 -8041 6506 -8033
rect 6578 -8033 6624 -8021
rect 6578 -8041 6584 -8033
rect 6618 -8041 6624 -8033
rect 6696 -8033 6742 -8021
rect 6696 -8041 6702 -8033
rect 6736 -8041 6742 -8033
rect 6814 -8033 6860 -8021
rect 6814 -8041 6820 -8033
rect 6854 -8041 6860 -8033
rect 6932 -8033 6978 -8021
rect 6932 -8041 6938 -8033
rect 6972 -8041 6978 -8033
rect 7050 -8033 7096 -8021
rect 7050 -8041 7056 -8033
rect 7090 -8041 7096 -8033
rect 7168 -8033 7214 -8021
rect 7168 -8041 7174 -8033
rect 7208 -8041 7214 -8033
rect 7286 -8033 7332 -8021
rect 7286 -8041 7292 -8033
rect 7326 -8041 7332 -8033
rect 7404 -8033 7450 -8021
rect 7404 -8041 7410 -8033
rect 7444 -8041 7450 -8033
rect 7522 -8033 7568 -8021
rect 7522 -8041 7528 -8033
rect 7562 -8041 7568 -8033
rect 7640 -8033 7686 -8021
rect 7640 -8041 7646 -8033
rect 7680 -8041 7686 -8033
rect 7868 -8033 7914 -8021
rect 7868 -8041 7874 -8033
rect 7908 -8041 7914 -8033
rect 7986 -8033 8032 -8021
rect 7986 -8041 7992 -8033
rect 8026 -8041 8032 -8033
rect 8104 -8033 8150 -8021
rect 8104 -8041 8110 -8033
rect 8144 -8041 8150 -8033
rect 8222 -8033 8268 -8021
rect 8222 -8041 8228 -8033
rect 8262 -8041 8268 -8033
rect 8340 -8033 8386 -8021
rect 8340 -8041 8346 -8033
rect 8380 -8041 8386 -8033
rect 8458 -8033 8504 -8021
rect 8458 -8041 8464 -8033
rect 8498 -8041 8504 -8033
rect 8576 -8033 8622 -8021
rect 8576 -8041 8582 -8033
rect 8616 -8041 8622 -8033
rect 8694 -8033 8740 -8021
rect 8694 -8041 8700 -8033
rect 8734 -8041 8740 -8033
rect 8812 -8033 8858 -8021
rect 8812 -8041 8818 -8033
rect 8852 -8041 8858 -8033
rect 8930 -8033 8976 -8021
rect 8930 -8041 8936 -8033
rect 8970 -8041 8976 -8033
rect 9048 -8033 9094 -8021
rect 9048 -8041 9054 -8033
rect 9088 -8041 9094 -8033
rect 9166 -8033 9212 -8021
rect 9166 -8041 9172 -8033
rect 9206 -8041 9212 -8033
rect 9284 -8033 9330 -8021
rect 9284 -8041 9290 -8033
rect 9324 -8041 9330 -8033
rect 9402 -8033 9448 -8021
rect 9402 -8041 9408 -8033
rect 9442 -8041 9448 -8033
rect 9520 -8033 9566 -8021
rect 9520 -8041 9526 -8033
rect 9560 -8041 9566 -8033
rect 9638 -8033 9684 -8021
rect 9638 -8041 9644 -8033
rect 9678 -8041 9684 -8033
rect 9796 -8037 9834 -8003
rect 9868 -8037 9906 -8003
rect 9940 -8037 9978 -8003
rect 10012 -8037 10050 -8003
rect 10084 -8037 10122 -8003
rect 10156 -8037 10194 -8003
rect 10228 -8037 10266 -8003
rect 10300 -8037 10338 -8003
rect 10372 -8037 10410 -8003
rect 10444 -8037 10482 -8003
rect 5444 -8051 5610 -8047
rect 4060 -8087 5610 -8051
rect 4060 -8103 4098 -8087
rect 4132 -8103 4170 -8087
rect 4204 -8103 4242 -8087
rect 4276 -8103 4314 -8087
rect 4348 -8103 4386 -8087
rect 4420 -8103 4458 -8087
rect 4492 -8103 4530 -8087
rect 4564 -8103 4602 -8087
rect 4636 -8103 4674 -8087
rect 4708 -8103 4746 -8087
rect 4780 -8103 4818 -8087
rect 4852 -8103 4890 -8087
rect 4924 -8103 4962 -8087
rect 4996 -8103 5034 -8087
rect 5068 -8103 5106 -8087
rect 5140 -8103 5178 -8087
rect 5212 -8103 5250 -8087
rect 5284 -8103 5322 -8087
rect 5356 -8103 5394 -8087
rect 5428 -8103 5466 -8087
rect 4060 -8155 4094 -8103
rect 4146 -8121 4170 -8103
rect 4227 -8121 4242 -8103
rect 4308 -8121 4314 -8103
rect 4492 -8121 4499 -8103
rect 4564 -8121 4580 -8103
rect 4636 -8121 4662 -8103
rect 4146 -8155 4175 -8121
rect 4227 -8155 4256 -8121
rect 4308 -8155 4337 -8121
rect 4389 -8155 4418 -8121
rect 4470 -8155 4499 -8121
rect 4551 -8155 4580 -8121
rect 4632 -8155 4662 -8121
rect 4714 -8155 4743 -8103
rect 4795 -8121 4818 -8103
rect 4876 -8121 4890 -8103
rect 4957 -8121 4962 -8103
rect 5140 -8121 5148 -8103
rect 5212 -8121 5230 -8103
rect 5284 -8121 5311 -8103
rect 4795 -8155 4824 -8121
rect 4876 -8155 4905 -8121
rect 4957 -8155 4986 -8121
rect 5038 -8155 5067 -8121
rect 5119 -8155 5148 -8121
rect 5200 -8155 5230 -8121
rect 5282 -8155 5311 -8121
rect 5363 -8155 5392 -8103
rect 5444 -8121 5466 -8103
rect 5500 -8121 5538 -8087
rect 5572 -8121 5610 -8087
rect 5444 -8155 5610 -8121
rect 4060 -8161 5610 -8155
rect 4060 -8195 4098 -8161
rect 4132 -8195 4170 -8161
rect 4204 -8195 4242 -8161
rect 4276 -8195 4314 -8161
rect 4348 -8195 4386 -8161
rect 4420 -8195 4458 -8161
rect 4492 -8195 4530 -8161
rect 4564 -8195 4602 -8161
rect 4636 -8195 4674 -8161
rect 4708 -8195 4746 -8161
rect 4780 -8195 4818 -8161
rect 4852 -8195 4890 -8161
rect 4924 -8195 4962 -8161
rect 4996 -8195 5034 -8161
rect 5068 -8195 5106 -8161
rect 5140 -8195 5178 -8161
rect 5212 -8195 5250 -8161
rect 5284 -8195 5322 -8161
rect 5356 -8195 5394 -8161
rect 5428 -8195 5466 -8161
rect 5500 -8195 5538 -8161
rect 5572 -8195 5610 -8161
rect 4060 -8207 5610 -8195
rect 4060 -8259 4094 -8207
rect 4146 -8235 4175 -8207
rect 4227 -8235 4256 -8207
rect 4308 -8235 4337 -8207
rect 4389 -8235 4418 -8207
rect 4470 -8235 4499 -8207
rect 4551 -8235 4580 -8207
rect 4632 -8235 4662 -8207
rect 4146 -8259 4170 -8235
rect 4227 -8259 4242 -8235
rect 4308 -8259 4314 -8235
rect 4492 -8259 4499 -8235
rect 4564 -8259 4580 -8235
rect 4636 -8259 4662 -8235
rect 4714 -8259 4743 -8207
rect 4795 -8235 4824 -8207
rect 4876 -8235 4905 -8207
rect 4957 -8235 4986 -8207
rect 5038 -8235 5067 -8207
rect 5119 -8235 5148 -8207
rect 5200 -8235 5230 -8207
rect 5282 -8235 5311 -8207
rect 4795 -8259 4818 -8235
rect 4876 -8259 4890 -8235
rect 4957 -8259 4962 -8235
rect 5140 -8259 5148 -8235
rect 5212 -8259 5230 -8235
rect 5284 -8259 5311 -8235
rect 5363 -8259 5392 -8207
rect 5444 -8235 5610 -8207
rect 5444 -8259 5466 -8235
rect 4060 -8269 4098 -8259
rect 4132 -8269 4170 -8259
rect 4204 -8269 4242 -8259
rect 4276 -8269 4314 -8259
rect 4348 -8269 4386 -8259
rect 4420 -8269 4458 -8259
rect 4492 -8269 4530 -8259
rect 4564 -8269 4602 -8259
rect 4636 -8269 4674 -8259
rect 4708 -8269 4746 -8259
rect 4780 -8269 4818 -8259
rect 4852 -8269 4890 -8259
rect 4924 -8269 4962 -8259
rect 4996 -8269 5034 -8259
rect 5068 -8269 5106 -8259
rect 5140 -8269 5178 -8259
rect 5212 -8269 5250 -8259
rect 5284 -8269 5322 -8259
rect 5356 -8269 5394 -8259
rect 5428 -8269 5466 -8259
rect 5500 -8269 5538 -8235
rect 5572 -8269 5610 -8235
rect 4060 -8309 5610 -8269
rect 4060 -8311 4098 -8309
rect 4132 -8311 4170 -8309
rect 4204 -8311 4242 -8309
rect 4276 -8311 4314 -8309
rect 4348 -8311 4386 -8309
rect 4420 -8311 4458 -8309
rect 4492 -8311 4530 -8309
rect 4564 -8311 4602 -8309
rect 4636 -8311 4674 -8309
rect 4708 -8311 4746 -8309
rect 4780 -8311 4818 -8309
rect 4852 -8311 4890 -8309
rect 4924 -8311 4962 -8309
rect 4996 -8311 5034 -8309
rect 5068 -8311 5106 -8309
rect 5140 -8311 5178 -8309
rect 5212 -8311 5250 -8309
rect 5284 -8311 5322 -8309
rect 5356 -8311 5394 -8309
rect 5428 -8311 5466 -8309
rect 4060 -8363 4094 -8311
rect 4146 -8343 4170 -8311
rect 4227 -8343 4242 -8311
rect 4308 -8343 4314 -8311
rect 4492 -8343 4499 -8311
rect 4564 -8343 4580 -8311
rect 4636 -8343 4662 -8311
rect 4146 -8363 4175 -8343
rect 4227 -8363 4256 -8343
rect 4308 -8363 4337 -8343
rect 4389 -8363 4418 -8343
rect 4470 -8363 4499 -8343
rect 4551 -8363 4580 -8343
rect 4632 -8363 4662 -8343
rect 4714 -8363 4743 -8311
rect 4795 -8343 4818 -8311
rect 4876 -8343 4890 -8311
rect 4957 -8343 4962 -8311
rect 5140 -8343 5148 -8311
rect 5212 -8343 5230 -8311
rect 5284 -8343 5311 -8311
rect 4795 -8363 4824 -8343
rect 4876 -8363 4905 -8343
rect 4957 -8363 4986 -8343
rect 5038 -8363 5067 -8343
rect 5119 -8363 5148 -8343
rect 5200 -8363 5230 -8343
rect 5282 -8363 5311 -8343
rect 5363 -8363 5392 -8311
rect 5444 -8343 5466 -8311
rect 5500 -8343 5538 -8309
rect 5572 -8343 5610 -8309
rect 5444 -8363 5610 -8343
rect 4060 -8383 5610 -8363
rect 4060 -8415 4098 -8383
rect 4132 -8415 4170 -8383
rect 4204 -8415 4242 -8383
rect 4276 -8415 4314 -8383
rect 4348 -8415 4386 -8383
rect 4420 -8415 4458 -8383
rect 4492 -8415 4530 -8383
rect 4564 -8415 4602 -8383
rect 4636 -8415 4674 -8383
rect 4708 -8415 4746 -8383
rect 4780 -8415 4818 -8383
rect 4852 -8415 4890 -8383
rect 4924 -8415 4962 -8383
rect 4996 -8415 5034 -8383
rect 5068 -8415 5106 -8383
rect 5140 -8415 5178 -8383
rect 5212 -8415 5250 -8383
rect 5284 -8415 5322 -8383
rect 5356 -8415 5394 -8383
rect 5428 -8415 5466 -8383
rect 4060 -8467 4094 -8415
rect 4146 -8417 4170 -8415
rect 4227 -8417 4242 -8415
rect 4308 -8417 4314 -8415
rect 4492 -8417 4499 -8415
rect 4564 -8417 4580 -8415
rect 4636 -8417 4662 -8415
rect 4146 -8457 4175 -8417
rect 4227 -8457 4256 -8417
rect 4308 -8457 4337 -8417
rect 4389 -8457 4418 -8417
rect 4470 -8457 4499 -8417
rect 4551 -8457 4580 -8417
rect 4632 -8457 4662 -8417
rect 4146 -8467 4170 -8457
rect 4227 -8467 4242 -8457
rect 4308 -8467 4314 -8457
rect 4492 -8467 4499 -8457
rect 4564 -8467 4580 -8457
rect 4636 -8467 4662 -8457
rect 4714 -8467 4743 -8415
rect 4795 -8417 4818 -8415
rect 4876 -8417 4890 -8415
rect 4957 -8417 4962 -8415
rect 5140 -8417 5148 -8415
rect 5212 -8417 5230 -8415
rect 5284 -8417 5311 -8415
rect 4795 -8457 4824 -8417
rect 4876 -8457 4905 -8417
rect 4957 -8457 4986 -8417
rect 5038 -8457 5067 -8417
rect 5119 -8457 5148 -8417
rect 5200 -8457 5230 -8417
rect 5282 -8457 5311 -8417
rect 4795 -8467 4818 -8457
rect 4876 -8467 4890 -8457
rect 4957 -8467 4962 -8457
rect 5140 -8467 5148 -8457
rect 5212 -8467 5230 -8457
rect 5284 -8467 5311 -8457
rect 5363 -8467 5392 -8415
rect 5444 -8417 5466 -8415
rect 5500 -8417 5538 -8383
rect 5572 -8417 5610 -8383
rect 5444 -8457 5610 -8417
rect 5444 -8467 5466 -8457
rect 4060 -8491 4098 -8467
rect 4132 -8491 4170 -8467
rect 4204 -8491 4242 -8467
rect 4276 -8491 4314 -8467
rect 4348 -8491 4386 -8467
rect 4420 -8491 4458 -8467
rect 4492 -8491 4530 -8467
rect 4564 -8491 4602 -8467
rect 4636 -8491 4674 -8467
rect 4708 -8491 4746 -8467
rect 4780 -8491 4818 -8467
rect 4852 -8491 4890 -8467
rect 4924 -8491 4962 -8467
rect 4996 -8491 5034 -8467
rect 5068 -8491 5106 -8467
rect 5140 -8491 5178 -8467
rect 5212 -8491 5250 -8467
rect 5284 -8491 5322 -8467
rect 5356 -8491 5394 -8467
rect 5428 -8491 5466 -8467
rect 5500 -8491 5538 -8457
rect 5572 -8491 5610 -8457
rect 4060 -8519 5610 -8491
rect 4060 -8571 4094 -8519
rect 4146 -8531 4175 -8519
rect 4227 -8531 4256 -8519
rect 4308 -8531 4337 -8519
rect 4389 -8531 4418 -8519
rect 4470 -8531 4499 -8519
rect 4551 -8531 4580 -8519
rect 4632 -8531 4662 -8519
rect 4146 -8565 4170 -8531
rect 4227 -8565 4242 -8531
rect 4308 -8565 4314 -8531
rect 4492 -8565 4499 -8531
rect 4564 -8565 4580 -8531
rect 4636 -8565 4662 -8531
rect 4146 -8571 4175 -8565
rect 4227 -8571 4256 -8565
rect 4308 -8571 4337 -8565
rect 4389 -8571 4418 -8565
rect 4470 -8571 4499 -8565
rect 4551 -8571 4580 -8565
rect 4632 -8571 4662 -8565
rect 4714 -8571 4743 -8519
rect 4795 -8531 4824 -8519
rect 4876 -8531 4905 -8519
rect 4957 -8531 4986 -8519
rect 5038 -8531 5067 -8519
rect 5119 -8531 5148 -8519
rect 5200 -8531 5230 -8519
rect 5282 -8531 5311 -8519
rect 4795 -8565 4818 -8531
rect 4876 -8565 4890 -8531
rect 4957 -8565 4962 -8531
rect 5140 -8565 5148 -8531
rect 5212 -8565 5230 -8531
rect 5284 -8565 5311 -8531
rect 4795 -8571 4824 -8565
rect 4876 -8571 4905 -8565
rect 4957 -8571 4986 -8565
rect 5038 -8571 5067 -8565
rect 5119 -8571 5148 -8565
rect 5200 -8571 5230 -8565
rect 5282 -8571 5311 -8565
rect 5363 -8571 5392 -8519
rect 5444 -8531 5610 -8519
rect 5444 -8565 5466 -8531
rect 5500 -8565 5538 -8531
rect 5572 -8565 5610 -8531
rect 5444 -8571 5610 -8565
rect 4060 -8585 5610 -8571
rect 4083 -8606 5471 -8585
rect 5857 -8601 5867 -8041
rect 5919 -8601 5929 -8041
rect 5975 -8601 5985 -8041
rect 6037 -8601 6047 -8041
rect 6093 -8601 6103 -8041
rect 6155 -8601 6165 -8041
rect 6211 -8601 6221 -8041
rect 6273 -8601 6283 -8041
rect 6329 -8601 6339 -8041
rect 6391 -8601 6401 -8041
rect 6447 -8601 6457 -8041
rect 6509 -8601 6519 -8041
rect 6565 -8601 6575 -8041
rect 6627 -8601 6637 -8041
rect 6683 -8601 6693 -8041
rect 6745 -8601 6755 -8041
rect 6801 -8601 6811 -8041
rect 6863 -8601 6873 -8041
rect 6919 -8601 6929 -8041
rect 6981 -8601 6991 -8041
rect 7037 -8601 7047 -8041
rect 7099 -8601 7109 -8041
rect 7155 -8601 7165 -8041
rect 7217 -8601 7227 -8041
rect 7273 -8601 7283 -8041
rect 7335 -8601 7345 -8041
rect 7391 -8601 7401 -8041
rect 7453 -8601 7463 -8041
rect 7509 -8601 7519 -8041
rect 7571 -8601 7581 -8041
rect 7627 -8601 7637 -8041
rect 7689 -8601 7699 -8041
rect 7855 -8601 7865 -8041
rect 7917 -8601 7927 -8041
rect 7973 -8601 7983 -8041
rect 8035 -8601 8045 -8041
rect 8091 -8601 8101 -8041
rect 8153 -8601 8163 -8041
rect 8209 -8601 8219 -8041
rect 8271 -8601 8281 -8041
rect 8327 -8601 8337 -8041
rect 8389 -8601 8399 -8041
rect 8445 -8601 8455 -8041
rect 8507 -8601 8517 -8041
rect 8563 -8601 8573 -8041
rect 8625 -8601 8635 -8041
rect 8681 -8601 8691 -8041
rect 8743 -8601 8753 -8041
rect 8799 -8601 8809 -8041
rect 8861 -8601 8871 -8041
rect 8917 -8601 8927 -8041
rect 8979 -8601 8989 -8041
rect 9035 -8601 9045 -8041
rect 9097 -8601 9107 -8041
rect 9153 -8601 9163 -8041
rect 9215 -8601 9225 -8041
rect 9271 -8601 9281 -8041
rect 9333 -8601 9343 -8041
rect 9389 -8601 9399 -8041
rect 9451 -8601 9461 -8041
rect 9507 -8601 9517 -8041
rect 9569 -8601 9579 -8041
rect 9625 -8601 9635 -8041
rect 9687 -8601 9697 -8041
rect 9796 -8077 10482 -8037
rect 12515 -8059 12525 -7219
rect 12577 -8059 12587 -7219
rect 12663 -8059 12673 -7219
rect 12725 -8059 12735 -7219
rect 12811 -8059 12821 -7219
rect 12873 -8059 12883 -7219
rect 12959 -8059 12969 -7219
rect 13021 -8059 13031 -7219
rect 13107 -8059 13117 -7219
rect 13169 -8059 13179 -7219
rect 13255 -8059 13265 -7219
rect 13317 -8059 13327 -7219
rect 13403 -8059 13413 -7219
rect 13465 -8059 13475 -7219
rect 13551 -8059 13561 -7219
rect 13613 -8059 13623 -7219
rect 13699 -8059 13709 -7219
rect 13761 -8059 13771 -7219
rect 13847 -8059 13857 -7219
rect 13909 -8059 13919 -7219
rect 13995 -8059 14005 -7219
rect 14057 -8059 14067 -7219
rect 14143 -8059 14153 -7219
rect 14205 -8059 14215 -7219
rect 14291 -8059 14301 -7219
rect 14353 -8059 14363 -7219
rect 14439 -8059 14449 -7219
rect 14501 -8059 14511 -7219
rect 14587 -8059 14597 -7219
rect 14649 -8059 14659 -7219
rect 14735 -8059 14745 -7219
rect 14797 -8059 14807 -7219
rect 14883 -8059 14893 -7219
rect 14945 -8059 14955 -7219
rect 15031 -8059 15041 -7219
rect 15093 -8059 15103 -7219
rect 15179 -8059 15189 -7219
rect 15241 -8059 15251 -7219
rect 15327 -8059 15337 -7219
rect 15389 -8059 15399 -7219
rect 15475 -8059 15485 -7219
rect 15537 -8059 15547 -7219
rect 15623 -8059 15633 -7219
rect 15685 -8059 15695 -7219
rect 15771 -8059 15781 -7219
rect 15833 -8059 15843 -7219
rect 15919 -8059 15929 -7219
rect 15981 -8059 15991 -7219
rect 16067 -8059 16077 -7219
rect 16129 -8059 16139 -7219
rect 16215 -8059 16225 -7219
rect 16277 -8059 16287 -7219
rect 16363 -8059 16373 -7219
rect 16425 -8059 16435 -7219
rect 16511 -8059 16521 -7219
rect 16573 -8059 16583 -7219
rect 16659 -8059 16669 -7219
rect 16721 -8059 16731 -7219
rect 16807 -8059 16817 -7219
rect 16869 -8059 16879 -7219
rect 16955 -8059 16965 -7219
rect 17017 -8059 17027 -7219
rect 17103 -8059 17113 -7219
rect 17165 -8059 17175 -7219
rect 17251 -8059 17261 -7219
rect 17313 -8059 17323 -7219
rect 17399 -8059 17409 -7219
rect 17461 -8059 17471 -7219
rect 17547 -8059 17557 -7219
rect 17609 -8059 17619 -7219
rect 17695 -8059 17705 -7219
rect 17757 -8059 17767 -7219
rect 17843 -8059 17853 -7219
rect 17905 -8059 17915 -7219
rect 17991 -8059 18001 -7219
rect 18053 -8059 18063 -7219
rect 18139 -8059 18149 -7219
rect 18201 -8059 18211 -7219
rect 18287 -8059 18297 -7219
rect 18349 -8059 18359 -7219
rect 18435 -8059 18445 -7219
rect 18497 -8059 18507 -7219
rect 18583 -8059 18593 -7219
rect 18645 -8059 18655 -7219
rect 18731 -8059 18741 -7219
rect 18793 -8059 18803 -7219
rect 18879 -8059 18889 -7219
rect 18941 -8059 18951 -7219
rect 19027 -8059 19037 -7219
rect 19089 -8059 19099 -7219
rect 19175 -8059 19185 -7219
rect 19237 -8059 19247 -7219
rect 19323 -8059 19333 -7219
rect 19385 -8059 19395 -7219
rect 19471 -8059 19481 -7219
rect 19533 -8059 19543 -7219
rect 19619 -8059 19629 -7219
rect 19681 -8059 19691 -7219
rect 19767 -8059 19777 -7219
rect 19829 -8059 19839 -7219
rect 19915 -8059 19925 -7219
rect 19977 -8059 19987 -7219
rect 20063 -8059 20073 -7219
rect 20125 -8059 20135 -7219
rect 20211 -8059 20221 -7219
rect 20273 -8059 20283 -7219
rect 20359 -8059 20369 -7219
rect 20421 -8059 20431 -7219
rect 20507 -8059 20517 -7219
rect 20569 -8059 20579 -7219
rect 20655 -8059 20665 -7219
rect 20717 -8059 20727 -7219
rect 20803 -8059 20813 -7219
rect 20865 -8059 20875 -7219
rect 20951 -8059 20961 -7219
rect 21013 -8059 21023 -7219
rect 21099 -8059 21109 -7219
rect 21161 -8059 21171 -7219
rect 21247 -8059 21257 -7219
rect 21309 -8059 21319 -7219
rect 21395 -8059 21405 -7219
rect 21457 -8059 21467 -7219
rect 21543 -8059 21553 -7219
rect 21605 -8059 21615 -7219
rect 21691 -8059 21701 -7219
rect 21753 -8059 21763 -7219
rect 21839 -8059 21849 -7219
rect 21901 -8059 21911 -7219
rect 21987 -8059 21997 -7219
rect 22049 -8059 22059 -7219
rect 22135 -8059 22145 -7219
rect 22197 -8059 22207 -7219
rect 22283 -8059 22293 -7219
rect 22345 -8059 22355 -7219
rect 22431 -8059 22441 -7219
rect 22493 -8059 22503 -7219
rect 22579 -8059 22589 -7219
rect 22641 -8059 22651 -7219
rect 22727 -8059 22737 -7219
rect 22789 -8059 22799 -7219
rect 22875 -8059 22885 -7219
rect 22937 -8059 22947 -7219
rect 23023 -8059 23033 -7219
rect 23085 -8059 23095 -7219
rect 23171 -8059 23181 -7219
rect 23233 -8059 23243 -7219
rect 23319 -8059 23329 -7219
rect 23381 -8059 23391 -7219
rect 23467 -8059 23477 -7219
rect 23529 -8059 23539 -7219
rect 23615 -8059 23625 -7219
rect 23677 -8059 23687 -7219
rect 9796 -8111 9834 -8077
rect 9868 -8111 9906 -8077
rect 9940 -8111 9978 -8077
rect 10012 -8111 10050 -8077
rect 10084 -8111 10122 -8077
rect 10156 -8111 10194 -8077
rect 10228 -8111 10266 -8077
rect 10300 -8111 10338 -8077
rect 10372 -8111 10410 -8077
rect 10444 -8111 10482 -8077
rect 12528 -8091 12534 -8059
rect 12568 -8091 12574 -8059
rect 12528 -8103 12574 -8091
rect 12676 -8091 12682 -8059
rect 12716 -8091 12722 -8059
rect 12676 -8103 12722 -8091
rect 12824 -8091 12830 -8059
rect 12864 -8091 12870 -8059
rect 12824 -8103 12870 -8091
rect 12972 -8091 12978 -8059
rect 13012 -8091 13018 -8059
rect 12972 -8103 13018 -8091
rect 13120 -8091 13126 -8059
rect 13160 -8091 13166 -8059
rect 13120 -8103 13166 -8091
rect 13268 -8091 13274 -8059
rect 13308 -8091 13314 -8059
rect 13268 -8103 13314 -8091
rect 13416 -8091 13422 -8059
rect 13456 -8091 13462 -8059
rect 13416 -8103 13462 -8091
rect 13564 -8091 13570 -8059
rect 13604 -8091 13610 -8059
rect 13564 -8103 13610 -8091
rect 13712 -8091 13718 -8059
rect 13752 -8091 13758 -8059
rect 13712 -8103 13758 -8091
rect 13860 -8091 13866 -8059
rect 13900 -8091 13906 -8059
rect 13860 -8103 13906 -8091
rect 14008 -8091 14014 -8059
rect 14048 -8091 14054 -8059
rect 14008 -8103 14054 -8091
rect 14156 -8091 14162 -8059
rect 14196 -8091 14202 -8059
rect 14156 -8103 14202 -8091
rect 14304 -8091 14310 -8059
rect 14344 -8091 14350 -8059
rect 14304 -8103 14350 -8091
rect 14452 -8091 14458 -8059
rect 14492 -8091 14498 -8059
rect 14452 -8103 14498 -8091
rect 14600 -8091 14606 -8059
rect 14640 -8091 14646 -8059
rect 14600 -8103 14646 -8091
rect 14748 -8091 14754 -8059
rect 14788 -8091 14794 -8059
rect 14748 -8103 14794 -8091
rect 14896 -8091 14902 -8059
rect 14936 -8091 14942 -8059
rect 14896 -8103 14942 -8091
rect 15044 -8091 15050 -8059
rect 15084 -8091 15090 -8059
rect 15044 -8103 15090 -8091
rect 15192 -8091 15198 -8059
rect 15232 -8091 15238 -8059
rect 15192 -8103 15238 -8091
rect 15340 -8091 15346 -8059
rect 15380 -8091 15386 -8059
rect 15340 -8103 15386 -8091
rect 15488 -8091 15494 -8059
rect 15528 -8091 15534 -8059
rect 15488 -8103 15534 -8091
rect 15636 -8091 15642 -8059
rect 15676 -8091 15682 -8059
rect 15636 -8103 15682 -8091
rect 15784 -8091 15790 -8059
rect 15824 -8091 15830 -8059
rect 15784 -8103 15830 -8091
rect 15932 -8091 15938 -8059
rect 15972 -8091 15978 -8059
rect 15932 -8103 15978 -8091
rect 16080 -8091 16086 -8059
rect 16120 -8091 16126 -8059
rect 16080 -8103 16126 -8091
rect 16228 -8091 16234 -8059
rect 16268 -8091 16274 -8059
rect 16228 -8103 16274 -8091
rect 16376 -8091 16382 -8059
rect 16416 -8091 16422 -8059
rect 16376 -8103 16422 -8091
rect 16524 -8091 16530 -8059
rect 16564 -8091 16570 -8059
rect 16524 -8103 16570 -8091
rect 16672 -8091 16678 -8059
rect 16712 -8091 16718 -8059
rect 16672 -8103 16718 -8091
rect 16820 -8091 16826 -8059
rect 16860 -8091 16866 -8059
rect 16820 -8103 16866 -8091
rect 16968 -8091 16974 -8059
rect 17008 -8091 17014 -8059
rect 16968 -8103 17014 -8091
rect 17116 -8091 17122 -8059
rect 17156 -8091 17162 -8059
rect 17116 -8103 17162 -8091
rect 17264 -8091 17270 -8059
rect 17304 -8091 17310 -8059
rect 17264 -8103 17310 -8091
rect 17412 -8091 17418 -8059
rect 17452 -8091 17458 -8059
rect 17412 -8103 17458 -8091
rect 17560 -8091 17566 -8059
rect 17600 -8091 17606 -8059
rect 17560 -8103 17606 -8091
rect 17708 -8091 17714 -8059
rect 17748 -8091 17754 -8059
rect 17708 -8103 17754 -8091
rect 17856 -8091 17862 -8059
rect 17896 -8091 17902 -8059
rect 17856 -8103 17902 -8091
rect 18004 -8091 18010 -8059
rect 18044 -8091 18050 -8059
rect 18004 -8103 18050 -8091
rect 18152 -8091 18158 -8059
rect 18192 -8091 18198 -8059
rect 18152 -8103 18198 -8091
rect 18300 -8091 18306 -8059
rect 18340 -8091 18346 -8059
rect 18300 -8103 18346 -8091
rect 18448 -8091 18454 -8059
rect 18488 -8091 18494 -8059
rect 18448 -8103 18494 -8091
rect 18596 -8091 18602 -8059
rect 18636 -8091 18642 -8059
rect 18596 -8103 18642 -8091
rect 18744 -8091 18750 -8059
rect 18784 -8091 18790 -8059
rect 18744 -8103 18790 -8091
rect 18892 -8091 18898 -8059
rect 18932 -8091 18938 -8059
rect 18892 -8103 18938 -8091
rect 19040 -8091 19046 -8059
rect 19080 -8091 19086 -8059
rect 19040 -8103 19086 -8091
rect 19188 -8091 19194 -8059
rect 19228 -8091 19234 -8059
rect 19188 -8103 19234 -8091
rect 19336 -8091 19342 -8059
rect 19376 -8091 19382 -8059
rect 19336 -8103 19382 -8091
rect 19484 -8091 19490 -8059
rect 19524 -8091 19530 -8059
rect 19484 -8103 19530 -8091
rect 19632 -8091 19638 -8059
rect 19672 -8091 19678 -8059
rect 19632 -8103 19678 -8091
rect 19780 -8091 19786 -8059
rect 19820 -8091 19826 -8059
rect 19780 -8103 19826 -8091
rect 19928 -8091 19934 -8059
rect 19968 -8091 19974 -8059
rect 19928 -8103 19974 -8091
rect 20076 -8091 20082 -8059
rect 20116 -8091 20122 -8059
rect 20076 -8103 20122 -8091
rect 20224 -8091 20230 -8059
rect 20264 -8091 20270 -8059
rect 20224 -8103 20270 -8091
rect 20372 -8091 20378 -8059
rect 20412 -8091 20418 -8059
rect 20372 -8103 20418 -8091
rect 20520 -8091 20526 -8059
rect 20560 -8091 20566 -8059
rect 20520 -8103 20566 -8091
rect 20668 -8091 20674 -8059
rect 20708 -8091 20714 -8059
rect 20668 -8103 20714 -8091
rect 20816 -8091 20822 -8059
rect 20856 -8091 20862 -8059
rect 20816 -8103 20862 -8091
rect 20964 -8091 20970 -8059
rect 21004 -8091 21010 -8059
rect 20964 -8103 21010 -8091
rect 21112 -8091 21118 -8059
rect 21152 -8091 21158 -8059
rect 21112 -8103 21158 -8091
rect 21260 -8091 21266 -8059
rect 21300 -8091 21306 -8059
rect 21260 -8103 21306 -8091
rect 21408 -8091 21414 -8059
rect 21448 -8091 21454 -8059
rect 21408 -8103 21454 -8091
rect 21556 -8091 21562 -8059
rect 21596 -8091 21602 -8059
rect 21556 -8103 21602 -8091
rect 21704 -8091 21710 -8059
rect 21744 -8091 21750 -8059
rect 21704 -8103 21750 -8091
rect 21852 -8091 21858 -8059
rect 21892 -8091 21898 -8059
rect 21852 -8103 21898 -8091
rect 22000 -8091 22006 -8059
rect 22040 -8091 22046 -8059
rect 22000 -8103 22046 -8091
rect 22148 -8091 22154 -8059
rect 22188 -8091 22194 -8059
rect 22148 -8103 22194 -8091
rect 22296 -8091 22302 -8059
rect 22336 -8091 22342 -8059
rect 22296 -8103 22342 -8091
rect 22444 -8091 22450 -8059
rect 22484 -8091 22490 -8059
rect 22444 -8103 22490 -8091
rect 22592 -8091 22598 -8059
rect 22632 -8091 22638 -8059
rect 22592 -8103 22638 -8091
rect 22740 -8091 22746 -8059
rect 22780 -8091 22786 -8059
rect 22740 -8103 22786 -8091
rect 22888 -8091 22894 -8059
rect 22928 -8091 22934 -8059
rect 22888 -8103 22934 -8091
rect 23036 -8091 23042 -8059
rect 23076 -8091 23082 -8059
rect 23036 -8103 23082 -8091
rect 23184 -8091 23190 -8059
rect 23224 -8091 23230 -8059
rect 23184 -8103 23230 -8091
rect 23332 -8091 23338 -8059
rect 23372 -8091 23378 -8059
rect 23332 -8103 23378 -8091
rect 23628 -8091 23634 -8059
rect 23668 -8091 23674 -8059
rect 23628 -8103 23674 -8091
rect 9796 -8151 10482 -8111
rect 9796 -8185 9834 -8151
rect 9868 -8185 9906 -8151
rect 9940 -8185 9978 -8151
rect 10012 -8185 10050 -8151
rect 10084 -8185 10122 -8151
rect 10156 -8185 10194 -8151
rect 10228 -8185 10266 -8151
rect 10300 -8185 10338 -8151
rect 10372 -8185 10410 -8151
rect 10444 -8185 10482 -8151
rect 9796 -8225 10482 -8185
rect 9796 -8259 9834 -8225
rect 9868 -8259 9906 -8225
rect 9940 -8259 9978 -8225
rect 10012 -8259 10050 -8225
rect 10084 -8259 10122 -8225
rect 10156 -8259 10194 -8225
rect 10228 -8259 10266 -8225
rect 10300 -8259 10338 -8225
rect 10372 -8259 10410 -8225
rect 10444 -8259 10482 -8225
rect 9796 -8299 10626 -8259
rect 12570 -8289 12580 -8135
rect 12670 -8289 12680 -8135
rect 12718 -8289 12728 -8135
rect 12818 -8289 12828 -8135
rect 12866 -8289 12876 -8135
rect 12966 -8289 12976 -8135
rect 13014 -8289 13024 -8135
rect 13114 -8289 13124 -8135
rect 13162 -8289 13172 -8135
rect 13262 -8289 13272 -8135
rect 13310 -8289 13320 -8135
rect 13410 -8289 13420 -8135
rect 13458 -8289 13468 -8135
rect 13558 -8289 13568 -8135
rect 13606 -8289 13616 -8135
rect 13706 -8289 13716 -8135
rect 13754 -8289 13764 -8135
rect 13854 -8289 13864 -8135
rect 13902 -8289 13912 -8135
rect 14002 -8289 14012 -8135
rect 14050 -8289 14060 -8135
rect 14150 -8289 14160 -8135
rect 14198 -8289 14208 -8135
rect 14298 -8289 14308 -8135
rect 14346 -8289 14356 -8135
rect 14446 -8289 14456 -8135
rect 14494 -8289 14504 -8135
rect 14594 -8289 14604 -8135
rect 14642 -8289 14652 -8135
rect 14742 -8289 14752 -8135
rect 14790 -8289 14800 -8135
rect 14890 -8289 14900 -8135
rect 14938 -8289 14948 -8135
rect 15038 -8289 15048 -8135
rect 15086 -8289 15096 -8135
rect 15186 -8289 15196 -8135
rect 15234 -8289 15244 -8135
rect 15334 -8289 15344 -8135
rect 15382 -8289 15392 -8135
rect 15482 -8289 15492 -8135
rect 15530 -8289 15540 -8135
rect 15630 -8289 15640 -8135
rect 15678 -8289 15688 -8135
rect 15778 -8289 15788 -8135
rect 15826 -8289 15836 -8135
rect 15926 -8289 15936 -8135
rect 15974 -8289 15984 -8135
rect 16074 -8289 16084 -8135
rect 16122 -8289 16132 -8135
rect 16222 -8289 16232 -8135
rect 16270 -8289 16280 -8135
rect 16370 -8289 16380 -8135
rect 16418 -8289 16428 -8135
rect 16518 -8289 16528 -8135
rect 16566 -8289 16576 -8135
rect 16666 -8289 16676 -8135
rect 16714 -8289 16724 -8135
rect 16814 -8289 16824 -8135
rect 16862 -8289 16872 -8135
rect 16962 -8289 16972 -8135
rect 17010 -8289 17020 -8135
rect 17110 -8289 17120 -8135
rect 17158 -8289 17168 -8135
rect 17258 -8289 17268 -8135
rect 17306 -8289 17316 -8135
rect 17406 -8289 17416 -8135
rect 17454 -8289 17464 -8135
rect 17554 -8289 17564 -8135
rect 17602 -8289 17612 -8135
rect 17702 -8289 17712 -8135
rect 17750 -8289 17760 -8135
rect 17850 -8289 17860 -8135
rect 17898 -8289 17908 -8135
rect 17998 -8289 18008 -8135
rect 18046 -8289 18056 -8135
rect 18146 -8289 18156 -8135
rect 18194 -8289 18204 -8135
rect 18294 -8289 18304 -8135
rect 18342 -8289 18352 -8135
rect 18442 -8289 18452 -8135
rect 18490 -8289 18500 -8135
rect 18590 -8289 18600 -8135
rect 18638 -8289 18648 -8135
rect 18738 -8289 18748 -8135
rect 18786 -8289 18796 -8135
rect 18886 -8289 18896 -8135
rect 18934 -8289 18944 -8135
rect 19034 -8289 19044 -8135
rect 19082 -8289 19092 -8135
rect 19182 -8289 19192 -8135
rect 19230 -8289 19240 -8135
rect 19330 -8289 19340 -8135
rect 19378 -8289 19388 -8135
rect 19478 -8289 19488 -8135
rect 19526 -8289 19536 -8135
rect 19626 -8289 19636 -8135
rect 19674 -8289 19684 -8135
rect 19774 -8289 19784 -8135
rect 19822 -8289 19832 -8135
rect 19922 -8289 19932 -8135
rect 19970 -8289 19980 -8135
rect 20070 -8289 20080 -8135
rect 20118 -8289 20128 -8135
rect 20218 -8289 20228 -8135
rect 20266 -8289 20276 -8135
rect 20366 -8289 20376 -8135
rect 20414 -8289 20424 -8135
rect 20514 -8289 20524 -8135
rect 20562 -8289 20572 -8135
rect 20662 -8289 20672 -8135
rect 20710 -8289 20720 -8135
rect 20810 -8289 20820 -8135
rect 20858 -8289 20868 -8135
rect 20958 -8289 20968 -8135
rect 21006 -8289 21016 -8135
rect 21106 -8289 21116 -8135
rect 21154 -8289 21164 -8135
rect 21254 -8289 21264 -8135
rect 21302 -8289 21312 -8135
rect 21402 -8289 21412 -8135
rect 21450 -8289 21460 -8135
rect 21550 -8289 21560 -8135
rect 21598 -8289 21608 -8135
rect 21698 -8289 21708 -8135
rect 21746 -8289 21756 -8135
rect 21846 -8289 21856 -8135
rect 21894 -8289 21904 -8135
rect 21994 -8289 22004 -8135
rect 22042 -8289 22052 -8135
rect 22142 -8289 22152 -8135
rect 22190 -8289 22200 -8135
rect 22290 -8289 22300 -8135
rect 22338 -8289 22348 -8135
rect 22438 -8289 22448 -8135
rect 22486 -8289 22496 -8135
rect 22586 -8289 22596 -8135
rect 22634 -8289 22644 -8135
rect 22734 -8289 22744 -8135
rect 22782 -8289 22792 -8135
rect 22882 -8289 22892 -8135
rect 22930 -8289 22940 -8135
rect 23030 -8289 23040 -8135
rect 23078 -8289 23088 -8135
rect 23178 -8289 23188 -8135
rect 23226 -8289 23236 -8135
rect 23326 -8289 23336 -8135
rect 23374 -8289 23384 -8135
rect 23474 -8289 23484 -8135
rect 23522 -8289 23532 -8135
rect 23622 -8289 23632 -8135
rect 9796 -8333 9834 -8299
rect 9868 -8333 9906 -8299
rect 9940 -8333 9978 -8299
rect 10012 -8333 10050 -8299
rect 10084 -8333 10122 -8299
rect 10156 -8333 10194 -8299
rect 10228 -8333 10266 -8299
rect 10300 -8333 10338 -8299
rect 10372 -8333 10410 -8299
rect 10444 -8333 10482 -8299
rect 10516 -8333 10554 -8299
rect 10588 -8333 10626 -8299
rect 9796 -8373 10626 -8333
rect 12528 -8333 12574 -8321
rect 12528 -8365 12534 -8333
rect 12568 -8365 12574 -8333
rect 12676 -8333 12722 -8321
rect 12676 -8365 12682 -8333
rect 12716 -8365 12722 -8333
rect 12824 -8333 12870 -8321
rect 12824 -8365 12830 -8333
rect 12864 -8365 12870 -8333
rect 12972 -8333 13018 -8321
rect 12972 -8365 12978 -8333
rect 13012 -8365 13018 -8333
rect 13120 -8333 13166 -8321
rect 13120 -8365 13126 -8333
rect 13160 -8365 13166 -8333
rect 13268 -8333 13314 -8321
rect 13268 -8365 13274 -8333
rect 13308 -8365 13314 -8333
rect 13416 -8333 13462 -8321
rect 13416 -8365 13422 -8333
rect 13456 -8365 13462 -8333
rect 13564 -8333 13610 -8321
rect 13564 -8365 13570 -8333
rect 13604 -8365 13610 -8333
rect 13712 -8333 13758 -8321
rect 13712 -8365 13718 -8333
rect 13752 -8365 13758 -8333
rect 13860 -8333 13906 -8321
rect 13860 -8365 13866 -8333
rect 13900 -8365 13906 -8333
rect 14008 -8333 14054 -8321
rect 14008 -8365 14014 -8333
rect 14048 -8365 14054 -8333
rect 14156 -8333 14202 -8321
rect 14156 -8365 14162 -8333
rect 14196 -8365 14202 -8333
rect 14304 -8333 14350 -8321
rect 14304 -8365 14310 -8333
rect 14344 -8365 14350 -8333
rect 14452 -8333 14498 -8321
rect 14452 -8365 14458 -8333
rect 14492 -8365 14498 -8333
rect 14600 -8333 14646 -8321
rect 14600 -8365 14606 -8333
rect 14640 -8365 14646 -8333
rect 14748 -8333 14794 -8321
rect 14748 -8365 14754 -8333
rect 14788 -8365 14794 -8333
rect 14896 -8333 14942 -8321
rect 14896 -8365 14902 -8333
rect 14936 -8365 14942 -8333
rect 15044 -8333 15090 -8321
rect 15044 -8365 15050 -8333
rect 15084 -8365 15090 -8333
rect 15192 -8333 15238 -8321
rect 15192 -8365 15198 -8333
rect 15232 -8365 15238 -8333
rect 15340 -8333 15386 -8321
rect 15340 -8365 15346 -8333
rect 15380 -8365 15386 -8333
rect 15488 -8333 15534 -8321
rect 15488 -8365 15494 -8333
rect 15528 -8365 15534 -8333
rect 15636 -8333 15682 -8321
rect 15636 -8365 15642 -8333
rect 15676 -8365 15682 -8333
rect 15784 -8333 15830 -8321
rect 15784 -8365 15790 -8333
rect 15824 -8365 15830 -8333
rect 15932 -8333 15978 -8321
rect 15932 -8365 15938 -8333
rect 15972 -8365 15978 -8333
rect 16080 -8333 16126 -8321
rect 16080 -8365 16086 -8333
rect 16120 -8365 16126 -8333
rect 16228 -8333 16274 -8321
rect 16228 -8365 16234 -8333
rect 16268 -8365 16274 -8333
rect 16376 -8333 16422 -8321
rect 16376 -8365 16382 -8333
rect 16416 -8365 16422 -8333
rect 16524 -8333 16570 -8321
rect 16524 -8365 16530 -8333
rect 16564 -8365 16570 -8333
rect 16672 -8333 16718 -8321
rect 16672 -8365 16678 -8333
rect 16712 -8365 16718 -8333
rect 16820 -8333 16866 -8321
rect 16820 -8365 16826 -8333
rect 16860 -8365 16866 -8333
rect 16968 -8333 17014 -8321
rect 16968 -8365 16974 -8333
rect 17008 -8365 17014 -8333
rect 17116 -8333 17162 -8321
rect 17116 -8365 17122 -8333
rect 17156 -8365 17162 -8333
rect 17264 -8333 17310 -8321
rect 17264 -8365 17270 -8333
rect 17304 -8365 17310 -8333
rect 17412 -8333 17458 -8321
rect 17412 -8365 17418 -8333
rect 17452 -8365 17458 -8333
rect 17560 -8333 17606 -8321
rect 17560 -8365 17566 -8333
rect 17600 -8365 17606 -8333
rect 17708 -8333 17754 -8321
rect 17708 -8365 17714 -8333
rect 17748 -8365 17754 -8333
rect 17856 -8333 17902 -8321
rect 17856 -8365 17862 -8333
rect 17896 -8365 17902 -8333
rect 18004 -8333 18050 -8321
rect 18004 -8365 18010 -8333
rect 18044 -8365 18050 -8333
rect 18152 -8333 18198 -8321
rect 18152 -8365 18158 -8333
rect 18192 -8365 18198 -8333
rect 18300 -8333 18346 -8321
rect 18300 -8365 18306 -8333
rect 18340 -8365 18346 -8333
rect 18448 -8333 18494 -8321
rect 18448 -8365 18454 -8333
rect 18488 -8365 18494 -8333
rect 18596 -8333 18642 -8321
rect 18596 -8365 18602 -8333
rect 18636 -8365 18642 -8333
rect 18744 -8333 18790 -8321
rect 18744 -8365 18750 -8333
rect 18784 -8365 18790 -8333
rect 18892 -8333 18938 -8321
rect 18892 -8365 18898 -8333
rect 18932 -8365 18938 -8333
rect 19040 -8333 19086 -8321
rect 19040 -8365 19046 -8333
rect 19080 -8365 19086 -8333
rect 19188 -8333 19234 -8321
rect 19188 -8365 19194 -8333
rect 19228 -8365 19234 -8333
rect 19336 -8333 19382 -8321
rect 19336 -8365 19342 -8333
rect 19376 -8365 19382 -8333
rect 19484 -8333 19530 -8321
rect 19484 -8365 19490 -8333
rect 19524 -8365 19530 -8333
rect 19632 -8333 19678 -8321
rect 19632 -8365 19638 -8333
rect 19672 -8365 19678 -8333
rect 19780 -8333 19826 -8321
rect 19780 -8365 19786 -8333
rect 19820 -8365 19826 -8333
rect 19928 -8333 19974 -8321
rect 19928 -8365 19934 -8333
rect 19968 -8365 19974 -8333
rect 20076 -8333 20122 -8321
rect 20076 -8365 20082 -8333
rect 20116 -8365 20122 -8333
rect 20224 -8333 20270 -8321
rect 20224 -8365 20230 -8333
rect 20264 -8365 20270 -8333
rect 20372 -8333 20418 -8321
rect 20372 -8365 20378 -8333
rect 20412 -8365 20418 -8333
rect 20520 -8333 20566 -8321
rect 20520 -8365 20526 -8333
rect 20560 -8365 20566 -8333
rect 20668 -8333 20714 -8321
rect 20668 -8365 20674 -8333
rect 20708 -8365 20714 -8333
rect 20816 -8333 20862 -8321
rect 20816 -8365 20822 -8333
rect 20856 -8365 20862 -8333
rect 20964 -8333 21010 -8321
rect 20964 -8365 20970 -8333
rect 21004 -8365 21010 -8333
rect 21112 -8333 21158 -8321
rect 21112 -8365 21118 -8333
rect 21152 -8365 21158 -8333
rect 21260 -8333 21306 -8321
rect 21260 -8365 21266 -8333
rect 21300 -8365 21306 -8333
rect 21408 -8333 21454 -8321
rect 21408 -8365 21414 -8333
rect 21448 -8365 21454 -8333
rect 21556 -8333 21602 -8321
rect 21556 -8365 21562 -8333
rect 21596 -8365 21602 -8333
rect 21704 -8333 21750 -8321
rect 21704 -8365 21710 -8333
rect 21744 -8365 21750 -8333
rect 21852 -8333 21898 -8321
rect 21852 -8365 21858 -8333
rect 21892 -8365 21898 -8333
rect 22000 -8333 22046 -8321
rect 22000 -8365 22006 -8333
rect 22040 -8365 22046 -8333
rect 22148 -8333 22194 -8321
rect 22148 -8365 22154 -8333
rect 22188 -8365 22194 -8333
rect 22296 -8333 22342 -8321
rect 22296 -8365 22302 -8333
rect 22336 -8365 22342 -8333
rect 22444 -8333 22490 -8321
rect 22444 -8365 22450 -8333
rect 22484 -8365 22490 -8333
rect 22592 -8333 22638 -8321
rect 22592 -8365 22598 -8333
rect 22632 -8365 22638 -8333
rect 22740 -8333 22786 -8321
rect 22740 -8365 22746 -8333
rect 22780 -8365 22786 -8333
rect 22888 -8333 22934 -8321
rect 22888 -8365 22894 -8333
rect 22928 -8365 22934 -8333
rect 23036 -8333 23082 -8321
rect 23036 -8365 23042 -8333
rect 23076 -8365 23082 -8333
rect 23184 -8333 23230 -8321
rect 23184 -8365 23190 -8333
rect 23224 -8365 23230 -8333
rect 23332 -8333 23378 -8321
rect 23332 -8365 23338 -8333
rect 23372 -8365 23378 -8333
rect 9796 -8407 9834 -8373
rect 9868 -8407 9906 -8373
rect 9940 -8407 9978 -8373
rect 10012 -8407 10050 -8373
rect 10084 -8407 10122 -8373
rect 10156 -8407 10194 -8373
rect 10228 -8407 10266 -8373
rect 10300 -8407 10338 -8373
rect 10372 -8407 10410 -8373
rect 10444 -8407 10482 -8373
rect 10516 -8407 10554 -8373
rect 10588 -8407 10626 -8373
rect 9796 -8447 10626 -8407
rect 9796 -8481 9834 -8447
rect 9868 -8481 9906 -8447
rect 9940 -8481 9978 -8447
rect 10012 -8481 10050 -8447
rect 10084 -8481 10122 -8447
rect 10156 -8481 10194 -8447
rect 10228 -8481 10266 -8447
rect 10300 -8481 10338 -8447
rect 10372 -8481 10410 -8447
rect 10444 -8481 10482 -8447
rect 10516 -8481 10554 -8447
rect 10588 -8481 10626 -8447
rect 9796 -8521 10626 -8481
rect 9796 -8555 9834 -8521
rect 9868 -8538 9906 -8521
rect 9940 -8538 9978 -8521
rect 10012 -8538 10050 -8521
rect 10084 -8538 10122 -8521
rect 10156 -8538 10194 -8521
rect 10228 -8538 10266 -8521
rect 10300 -8538 10338 -8521
rect 10372 -8538 10410 -8521
rect 10444 -8538 10482 -8521
rect 10516 -8538 10554 -8521
rect 10588 -8538 10626 -8521
rect 9891 -8555 9906 -8538
rect 9971 -8555 9978 -8538
rect 10156 -8555 10159 -8538
rect 10228 -8555 10239 -8538
rect 10300 -8555 10319 -8538
rect 10372 -8555 10399 -8538
rect 9796 -8590 9839 -8555
rect 9891 -8590 9919 -8555
rect 9971 -8590 9999 -8555
rect 10051 -8590 10079 -8555
rect 10131 -8590 10159 -8555
rect 10211 -8590 10239 -8555
rect 10291 -8590 10319 -8555
rect 10371 -8590 10399 -8555
rect 10451 -8590 10479 -8538
rect 10531 -8555 10554 -8538
rect 10531 -8590 10559 -8555
rect 10611 -8590 10626 -8538
rect 9796 -8595 10626 -8590
rect 5870 -8609 5876 -8601
rect 5910 -8609 5916 -8601
rect 5870 -8621 5916 -8609
rect 5988 -8609 5994 -8601
rect 6028 -8609 6034 -8601
rect 5988 -8621 6034 -8609
rect 6106 -8609 6112 -8601
rect 6146 -8609 6152 -8601
rect 6106 -8621 6152 -8609
rect 6224 -8609 6230 -8601
rect 6264 -8609 6270 -8601
rect 6224 -8621 6270 -8609
rect 6342 -8609 6348 -8601
rect 6382 -8609 6388 -8601
rect 6342 -8621 6388 -8609
rect 6460 -8609 6466 -8601
rect 6500 -8609 6506 -8601
rect 6460 -8621 6506 -8609
rect 6578 -8609 6584 -8601
rect 6618 -8609 6624 -8601
rect 6578 -8621 6624 -8609
rect 6696 -8609 6702 -8601
rect 6736 -8609 6742 -8601
rect 6696 -8621 6742 -8609
rect 6814 -8609 6820 -8601
rect 6854 -8609 6860 -8601
rect 6814 -8621 6860 -8609
rect 6932 -8609 6938 -8601
rect 6972 -8609 6978 -8601
rect 6932 -8621 6978 -8609
rect 7050 -8609 7056 -8601
rect 7090 -8609 7096 -8601
rect 7050 -8621 7096 -8609
rect 7168 -8609 7174 -8601
rect 7208 -8609 7214 -8601
rect 7168 -8621 7214 -8609
rect 7286 -8609 7292 -8601
rect 7326 -8609 7332 -8601
rect 7286 -8621 7332 -8609
rect 7404 -8609 7410 -8601
rect 7444 -8609 7450 -8601
rect 7404 -8621 7450 -8609
rect 7522 -8609 7528 -8601
rect 7562 -8609 7568 -8601
rect 7522 -8621 7568 -8609
rect 7640 -8609 7646 -8601
rect 7680 -8609 7686 -8601
rect 7640 -8621 7686 -8609
rect 7868 -8609 7874 -8601
rect 7908 -8609 7914 -8601
rect 7868 -8621 7914 -8609
rect 7986 -8609 7992 -8601
rect 8026 -8609 8032 -8601
rect 7986 -8621 8032 -8609
rect 8104 -8609 8110 -8601
rect 8144 -8609 8150 -8601
rect 8104 -8621 8150 -8609
rect 8222 -8609 8228 -8601
rect 8262 -8609 8268 -8601
rect 8222 -8621 8268 -8609
rect 8340 -8609 8346 -8601
rect 8380 -8609 8386 -8601
rect 8340 -8621 8386 -8609
rect 8458 -8609 8464 -8601
rect 8498 -8609 8504 -8601
rect 8458 -8621 8504 -8609
rect 8576 -8609 8582 -8601
rect 8616 -8609 8622 -8601
rect 8576 -8621 8622 -8609
rect 8694 -8609 8700 -8601
rect 8734 -8609 8740 -8601
rect 8694 -8621 8740 -8609
rect 8812 -8609 8818 -8601
rect 8852 -8609 8858 -8601
rect 8812 -8621 8858 -8609
rect 8930 -8609 8936 -8601
rect 8970 -8609 8976 -8601
rect 8930 -8621 8976 -8609
rect 9048 -8609 9054 -8601
rect 9088 -8609 9094 -8601
rect 9048 -8621 9094 -8609
rect 9166 -8609 9172 -8601
rect 9206 -8609 9212 -8601
rect 9166 -8621 9212 -8609
rect 9284 -8609 9290 -8601
rect 9324 -8609 9330 -8601
rect 9284 -8621 9330 -8609
rect 9402 -8609 9408 -8601
rect 9442 -8609 9448 -8601
rect 9402 -8621 9448 -8609
rect 9520 -8609 9526 -8601
rect 9560 -8609 9566 -8601
rect 9520 -8621 9566 -8609
rect 9638 -8609 9644 -8601
rect 9678 -8609 9684 -8601
rect 9638 -8621 9684 -8609
rect 9796 -8629 9834 -8595
rect 9868 -8617 9906 -8595
rect 9940 -8617 9978 -8595
rect 10012 -8617 10050 -8595
rect 10084 -8617 10122 -8595
rect 10156 -8617 10194 -8595
rect 10228 -8617 10266 -8595
rect 10300 -8617 10338 -8595
rect 10372 -8617 10410 -8595
rect 10444 -8617 10482 -8595
rect 10516 -8617 10554 -8595
rect 10588 -8617 10626 -8595
rect 9891 -8629 9906 -8617
rect 9971 -8629 9978 -8617
rect 10156 -8629 10159 -8617
rect 10228 -8629 10239 -8617
rect 10300 -8629 10319 -8617
rect 10372 -8629 10399 -8617
rect 9796 -8669 9839 -8629
rect 9891 -8669 9919 -8629
rect 9971 -8669 9999 -8629
rect 10051 -8669 10079 -8629
rect 10131 -8669 10159 -8629
rect 10211 -8669 10239 -8629
rect 10291 -8669 10319 -8629
rect 10371 -8669 10399 -8629
rect 10451 -8669 10479 -8617
rect 10531 -8629 10554 -8617
rect 10531 -8669 10559 -8629
rect 10611 -8669 10626 -8617
rect 9796 -8703 9834 -8669
rect 9868 -8703 9906 -8669
rect 9940 -8703 9978 -8669
rect 10012 -8703 10050 -8669
rect 10084 -8703 10122 -8669
rect 10156 -8703 10194 -8669
rect 10228 -8703 10266 -8669
rect 10300 -8703 10338 -8669
rect 10372 -8703 10410 -8669
rect 10444 -8703 10482 -8669
rect 10516 -8703 10554 -8669
rect 10588 -8703 10626 -8669
rect 9796 -8723 10626 -8703
rect 4056 -8871 5600 -8812
rect 5745 -8829 10875 -8815
rect 4056 -8876 4080 -8871
rect 4056 -8905 4080 -8878
rect 4114 -8876 4152 -8871
rect 4114 -8905 4152 -8878
rect 4186 -8876 4234 -8871
rect 4186 -8905 4234 -8878
rect 4268 -8876 4306 -8871
rect 4268 -8905 4306 -8878
rect 4340 -8876 4388 -8871
rect 4340 -8905 4388 -8878
rect 4422 -8876 4460 -8871
rect 4422 -8905 4460 -8878
rect 4494 -8876 4542 -8871
rect 4494 -8905 4542 -8878
rect 4576 -8876 4614 -8871
rect 4576 -8905 4614 -8878
rect 4648 -8876 4696 -8871
rect 4648 -8905 4696 -8878
rect 4730 -8876 4768 -8871
rect 4730 -8905 4768 -8878
rect 4802 -8876 4850 -8871
rect 4802 -8905 4850 -8878
rect 4884 -8876 4922 -8871
rect 4884 -8905 4922 -8878
rect 4956 -8876 5004 -8871
rect 4956 -8905 5004 -8878
rect 5038 -8876 5076 -8871
rect 5038 -8905 5076 -8878
rect 5110 -8876 5158 -8871
rect 5110 -8905 5158 -8878
rect 5192 -8876 5230 -8871
rect 5192 -8905 5230 -8878
rect 5264 -8876 5312 -8871
rect 5264 -8905 5312 -8878
rect 5346 -8876 5384 -8871
rect 5346 -8905 5384 -8878
rect 5418 -8876 5466 -8871
rect 5418 -8905 5466 -8878
rect 5500 -8876 5538 -8871
rect 5500 -8905 5538 -8878
rect 5572 -8876 5600 -8871
rect 5572 -8905 5620 -8878
rect 5654 -8905 5692 -8878
rect 5745 -8878 5759 -8829
rect 5726 -8881 5759 -8878
rect 5811 -8881 5839 -8829
rect 5891 -8881 5919 -8829
rect 5971 -8881 5999 -8829
rect 6051 -8881 6079 -8829
rect 6131 -8881 6159 -8829
rect 6211 -8881 6239 -8829
rect 6291 -8881 6319 -8829
rect 6371 -8881 6399 -8829
rect 6451 -8881 6479 -8829
rect 6531 -8881 6559 -8829
rect 6611 -8881 6639 -8829
rect 6691 -8881 6719 -8829
rect 6771 -8881 6799 -8829
rect 6851 -8881 6879 -8829
rect 6931 -8881 6959 -8829
rect 7011 -8881 7039 -8829
rect 7091 -8881 7119 -8829
rect 7171 -8881 7199 -8829
rect 7251 -8881 7279 -8829
rect 7331 -8881 7359 -8829
rect 7411 -8881 7439 -8829
rect 7491 -8881 7519 -8829
rect 7571 -8881 7599 -8829
rect 7651 -8881 7679 -8829
rect 7731 -8881 7759 -8829
rect 7811 -8881 7839 -8829
rect 7891 -8881 7919 -8829
rect 7971 -8881 7999 -8829
rect 8051 -8881 8079 -8829
rect 8131 -8881 8159 -8829
rect 8211 -8881 8239 -8829
rect 8291 -8881 8319 -8829
rect 8371 -8881 8399 -8829
rect 8451 -8881 8479 -8829
rect 8531 -8881 8559 -8829
rect 8611 -8881 8639 -8829
rect 8691 -8881 8719 -8829
rect 8771 -8881 8799 -8829
rect 8851 -8881 8879 -8829
rect 8931 -8881 8959 -8829
rect 9011 -8881 9039 -8829
rect 9091 -8881 9119 -8829
rect 9171 -8881 9199 -8829
rect 9251 -8881 9279 -8829
rect 9331 -8881 9359 -8829
rect 9411 -8881 9439 -8829
rect 9491 -8881 9519 -8829
rect 9571 -8881 9599 -8829
rect 9651 -8881 9679 -8829
rect 9731 -8881 9759 -8829
rect 9811 -8881 9839 -8829
rect 9891 -8881 9919 -8829
rect 9971 -8881 9999 -8829
rect 10051 -8881 10079 -8829
rect 10131 -8881 10159 -8829
rect 10211 -8881 10239 -8829
rect 10291 -8881 10319 -8829
rect 10371 -8881 10399 -8829
rect 10451 -8881 10479 -8829
rect 10531 -8881 10559 -8829
rect 10611 -8881 10639 -8829
rect 10691 -8881 10719 -8829
rect 10771 -8881 10799 -8829
rect 10851 -8881 10875 -8829
rect 5726 -8905 10875 -8881
rect 4056 -8909 10875 -8905
rect 4056 -8945 5759 -8909
rect 4056 -8969 4080 -8945
rect 4114 -8969 4152 -8945
rect 4186 -8969 4234 -8945
rect 4268 -8969 4306 -8945
rect 4340 -8969 4388 -8945
rect 4422 -8969 4460 -8945
rect 4494 -8969 4542 -8945
rect 4576 -8969 4614 -8945
rect 4648 -8969 4696 -8945
rect 4730 -8969 4768 -8945
rect 4802 -8969 4850 -8945
rect 4884 -8969 4922 -8945
rect 4956 -8969 5004 -8945
rect 5038 -8969 5076 -8945
rect 5110 -8969 5158 -8945
rect 5192 -8969 5230 -8945
rect 5264 -8969 5312 -8945
rect 5346 -8969 5384 -8945
rect 5418 -8969 5466 -8945
rect 5500 -8969 5538 -8945
rect 5572 -8969 5620 -8945
rect 5654 -8969 5692 -8945
rect 5726 -8961 5759 -8945
rect 5811 -8961 5839 -8909
rect 5891 -8961 5919 -8909
rect 5971 -8961 5999 -8909
rect 6051 -8961 6079 -8909
rect 6131 -8945 6159 -8909
rect 6211 -8945 6239 -8909
rect 6291 -8945 6319 -8909
rect 6371 -8945 6399 -8909
rect 6451 -8945 6479 -8909
rect 6531 -8945 6559 -8909
rect 6611 -8945 6639 -8909
rect 6691 -8945 6719 -8909
rect 6771 -8945 6799 -8909
rect 6851 -8945 6879 -8909
rect 6931 -8945 6959 -8909
rect 7011 -8945 7039 -8909
rect 7091 -8945 7119 -8909
rect 7171 -8945 7199 -8909
rect 7251 -8945 7279 -8909
rect 7331 -8945 7359 -8909
rect 7411 -8945 7439 -8909
rect 7491 -8945 7519 -8909
rect 7571 -8945 7599 -8909
rect 7651 -8945 7679 -8909
rect 6131 -8961 6154 -8945
rect 6211 -8961 6236 -8945
rect 6291 -8961 6308 -8945
rect 6371 -8961 6390 -8945
rect 6451 -8961 6462 -8945
rect 6531 -8961 6544 -8945
rect 6611 -8961 6616 -8945
rect 6691 -8961 6698 -8945
rect 6851 -8961 6852 -8945
rect 6958 -8961 6959 -8945
rect 7112 -8961 7119 -8945
rect 7194 -8961 7199 -8945
rect 7266 -8961 7279 -8945
rect 7348 -8961 7359 -8945
rect 7420 -8961 7439 -8945
rect 7502 -8961 7519 -8945
rect 7574 -8961 7599 -8945
rect 7656 -8961 7679 -8945
rect 7731 -8961 7759 -8909
rect 7811 -8961 7839 -8909
rect 7891 -8961 7919 -8909
rect 7971 -8961 7999 -8909
rect 8051 -8961 8079 -8909
rect 8131 -8945 8159 -8909
rect 8211 -8945 8239 -8909
rect 8291 -8945 8319 -8909
rect 8371 -8945 8399 -8909
rect 8451 -8945 8479 -8909
rect 8531 -8945 8559 -8909
rect 8611 -8945 8639 -8909
rect 8691 -8945 8719 -8909
rect 8771 -8945 8799 -8909
rect 8851 -8945 8879 -8909
rect 8931 -8945 8959 -8909
rect 9011 -8945 9039 -8909
rect 9091 -8945 9119 -8909
rect 9171 -8945 9199 -8909
rect 9251 -8945 9279 -8909
rect 9331 -8945 9359 -8909
rect 9411 -8945 9439 -8909
rect 9491 -8945 9519 -8909
rect 9571 -8945 9599 -8909
rect 9651 -8945 9679 -8909
rect 8131 -8961 8156 -8945
rect 8211 -8961 8238 -8945
rect 8291 -8961 8310 -8945
rect 8371 -8961 8392 -8945
rect 8451 -8961 8464 -8945
rect 8531 -8961 8546 -8945
rect 8611 -8961 8618 -8945
rect 8691 -8961 8700 -8945
rect 8771 -8961 8772 -8945
rect 8851 -8961 8854 -8945
rect 9114 -8961 9119 -8945
rect 9196 -8961 9199 -8945
rect 9268 -8961 9279 -8945
rect 9350 -8961 9359 -8945
rect 9422 -8961 9439 -8945
rect 9504 -8961 9519 -8945
rect 9576 -8961 9599 -8945
rect 9658 -8961 9679 -8945
rect 9731 -8961 9759 -8909
rect 9811 -8945 9839 -8909
rect 9812 -8961 9839 -8945
rect 9891 -8961 9919 -8909
rect 9971 -8961 9999 -8909
rect 10051 -8961 10079 -8909
rect 10131 -8945 10159 -8909
rect 10131 -8961 10158 -8945
rect 10211 -8961 10239 -8909
rect 10291 -8945 10319 -8909
rect 10371 -8945 10399 -8909
rect 10451 -8945 10479 -8909
rect 10531 -8945 10559 -8909
rect 10611 -8945 10639 -8909
rect 10691 -8945 10719 -8909
rect 10771 -8945 10799 -8909
rect 10851 -8945 10875 -8909
rect 10291 -8961 10312 -8945
rect 10371 -8961 10394 -8945
rect 10451 -8961 10466 -8945
rect 10531 -8961 10548 -8945
rect 10611 -8961 10620 -8945
rect 10691 -8961 10702 -8945
rect 10771 -8961 10774 -8945
rect 10851 -8961 10856 -8945
rect 5726 -8969 5774 -8961
rect 5745 -8975 5774 -8969
rect 5808 -8975 5846 -8961
rect 5880 -8975 5928 -8961
rect 5962 -8975 6000 -8961
rect 6034 -8975 6082 -8961
rect 6116 -8975 6154 -8961
rect 6188 -8975 6236 -8961
rect 6270 -8975 6308 -8961
rect 6342 -8975 6390 -8961
rect 6424 -8975 6462 -8961
rect 6496 -8975 6544 -8961
rect 6578 -8975 6616 -8961
rect 6650 -8975 6698 -8961
rect 6732 -8975 6770 -8961
rect 6804 -8975 6852 -8961
rect 6886 -8975 6924 -8961
rect 6958 -8975 7006 -8961
rect 7040 -8975 7078 -8961
rect 7112 -8975 7160 -8961
rect 7194 -8975 7232 -8961
rect 7266 -8975 7314 -8961
rect 7348 -8975 7386 -8961
rect 7420 -8975 7468 -8961
rect 7502 -8975 7540 -8961
rect 7574 -8975 7622 -8961
rect 7656 -8975 7694 -8961
rect 7728 -8975 7776 -8961
rect 7810 -8975 7848 -8961
rect 7882 -8975 7930 -8961
rect 7964 -8975 8002 -8961
rect 8036 -8975 8084 -8961
rect 8118 -8975 8156 -8961
rect 8190 -8975 8238 -8961
rect 8272 -8975 8310 -8961
rect 8344 -8975 8392 -8961
rect 8426 -8975 8464 -8961
rect 8498 -8975 8546 -8961
rect 8580 -8975 8618 -8961
rect 8652 -8975 8700 -8961
rect 8734 -8975 8772 -8961
rect 8806 -8975 8854 -8961
rect 8888 -8975 8926 -8961
rect 8960 -8975 9008 -8961
rect 9042 -8975 9080 -8961
rect 9114 -8975 9162 -8961
rect 9196 -8975 9234 -8961
rect 9268 -8975 9316 -8961
rect 9350 -8975 9388 -8961
rect 9422 -8975 9470 -8961
rect 9504 -8975 9542 -8961
rect 9576 -8975 9624 -8961
rect 9658 -8975 9696 -8961
rect 9730 -8975 9778 -8961
rect 9812 -8975 9850 -8961
rect 9884 -8975 9932 -8961
rect 9966 -8975 10004 -8961
rect 10038 -8975 10086 -8961
rect 10120 -8975 10158 -8961
rect 10192 -8975 10240 -8961
rect 10274 -8975 10312 -8961
rect 10346 -8975 10394 -8961
rect 10428 -8975 10466 -8961
rect 10500 -8975 10548 -8961
rect 10582 -8975 10620 -8961
rect 10654 -8975 10702 -8961
rect 10736 -8975 10774 -8961
rect 10808 -8975 10856 -8961
rect 12515 -9205 12525 -8365
rect 12577 -9205 12587 -8365
rect 12663 -9205 12673 -8365
rect 12725 -9205 12735 -8365
rect 12811 -9205 12821 -8365
rect 12873 -9205 12883 -8365
rect 12959 -9205 12969 -8365
rect 13021 -9205 13031 -8365
rect 13107 -9205 13117 -8365
rect 13169 -9205 13179 -8365
rect 13255 -9205 13265 -8365
rect 13317 -9205 13327 -8365
rect 13403 -9205 13413 -8365
rect 13465 -9205 13475 -8365
rect 13551 -9205 13561 -8365
rect 13613 -9205 13623 -8365
rect 13699 -9205 13709 -8365
rect 13761 -9205 13771 -8365
rect 13847 -9205 13857 -8365
rect 13909 -9205 13919 -8365
rect 13995 -9205 14005 -8365
rect 14057 -9205 14067 -8365
rect 14143 -9205 14153 -8365
rect 14205 -9205 14215 -8365
rect 14291 -9205 14301 -8365
rect 14353 -9205 14363 -8365
rect 14439 -9205 14449 -8365
rect 14501 -9205 14511 -8365
rect 14587 -9205 14597 -8365
rect 14649 -9205 14659 -8365
rect 14735 -9205 14745 -8365
rect 14797 -9205 14807 -8365
rect 14883 -9205 14893 -8365
rect 14945 -9205 14955 -8365
rect 15031 -9205 15041 -8365
rect 15093 -9205 15103 -8365
rect 15179 -9205 15189 -8365
rect 15241 -9205 15251 -8365
rect 15327 -9205 15337 -8365
rect 15389 -9205 15399 -8365
rect 15475 -9205 15485 -8365
rect 15537 -9205 15547 -8365
rect 15623 -9205 15633 -8365
rect 15685 -9205 15695 -8365
rect 15771 -9205 15781 -8365
rect 15833 -9205 15843 -8365
rect 15919 -9205 15929 -8365
rect 15981 -9205 15991 -8365
rect 16067 -9205 16077 -8365
rect 16129 -9205 16139 -8365
rect 16215 -9205 16225 -8365
rect 16277 -9205 16287 -8365
rect 16363 -9205 16373 -8365
rect 16425 -9205 16435 -8365
rect 16511 -9205 16521 -8365
rect 16573 -9205 16583 -8365
rect 16659 -9205 16669 -8365
rect 16721 -9205 16731 -8365
rect 16807 -9205 16817 -8365
rect 16869 -9205 16879 -8365
rect 16955 -9205 16965 -8365
rect 17017 -9205 17027 -8365
rect 17103 -9205 17113 -8365
rect 17165 -9205 17175 -8365
rect 17251 -9205 17261 -8365
rect 17313 -9205 17323 -8365
rect 17399 -9205 17409 -8365
rect 17461 -9205 17471 -8365
rect 17547 -9205 17557 -8365
rect 17609 -9205 17619 -8365
rect 17695 -9205 17705 -8365
rect 17757 -9205 17767 -8365
rect 17843 -9205 17853 -8365
rect 17905 -9205 17915 -8365
rect 17991 -9205 18001 -8365
rect 18053 -9205 18063 -8365
rect 18139 -9205 18149 -8365
rect 18201 -9205 18211 -8365
rect 18287 -9205 18297 -8365
rect 18349 -9205 18359 -8365
rect 18435 -9205 18445 -8365
rect 18497 -9205 18507 -8365
rect 18583 -9205 18593 -8365
rect 18645 -9205 18655 -8365
rect 18731 -9205 18741 -8365
rect 18793 -9205 18803 -8365
rect 18879 -9205 18889 -8365
rect 18941 -9205 18951 -8365
rect 19027 -9205 19037 -8365
rect 19089 -9205 19099 -8365
rect 19175 -9205 19185 -8365
rect 19237 -9205 19247 -8365
rect 19323 -9205 19333 -8365
rect 19385 -9205 19395 -8365
rect 19471 -9205 19481 -8365
rect 19533 -9205 19543 -8365
rect 19619 -9205 19629 -8365
rect 19681 -9205 19691 -8365
rect 19767 -9205 19777 -8365
rect 19829 -9205 19839 -8365
rect 19915 -9205 19925 -8365
rect 19977 -9205 19987 -8365
rect 20063 -9205 20073 -8365
rect 20125 -9205 20135 -8365
rect 20211 -9205 20221 -8365
rect 20273 -9205 20283 -8365
rect 20359 -9205 20369 -8365
rect 20421 -9205 20431 -8365
rect 20507 -9205 20517 -8365
rect 20569 -9205 20579 -8365
rect 20655 -9205 20665 -8365
rect 20717 -9205 20727 -8365
rect 20803 -9205 20813 -8365
rect 20865 -9205 20875 -8365
rect 20951 -9205 20961 -8365
rect 21013 -9205 21023 -8365
rect 21099 -9205 21109 -8365
rect 21161 -9205 21171 -8365
rect 21247 -9205 21257 -8365
rect 21309 -9205 21319 -8365
rect 21395 -9205 21405 -8365
rect 21457 -9205 21467 -8365
rect 21543 -9205 21553 -8365
rect 21605 -9205 21615 -8365
rect 21691 -9205 21701 -8365
rect 21753 -9205 21763 -8365
rect 21839 -9205 21849 -8365
rect 21901 -9205 21911 -8365
rect 21987 -9205 21997 -8365
rect 22049 -9205 22059 -8365
rect 22135 -9205 22145 -8365
rect 22197 -9205 22207 -8365
rect 22283 -9205 22293 -8365
rect 22345 -9205 22355 -8365
rect 22431 -9205 22441 -8365
rect 22493 -9205 22503 -8365
rect 22579 -9205 22589 -8365
rect 22641 -9205 22651 -8365
rect 22727 -9205 22737 -8365
rect 22789 -9205 22799 -8365
rect 22875 -9205 22885 -8365
rect 22937 -9205 22947 -8365
rect 23023 -9205 23033 -8365
rect 23085 -9205 23095 -8365
rect 23171 -9205 23181 -8365
rect 23233 -9205 23243 -8365
rect 23319 -9205 23329 -8365
rect 23381 -9205 23391 -8365
rect 23467 -9205 23477 -8365
rect 23529 -9205 23539 -8365
rect 23615 -9205 23625 -8365
rect 23677 -9205 23687 -8365
rect 12528 -9209 12534 -9205
rect 12568 -9209 12574 -9205
rect 12528 -9221 12574 -9209
rect 12676 -9209 12682 -9205
rect 12716 -9209 12722 -9205
rect 12676 -9221 12722 -9209
rect 12824 -9209 12830 -9205
rect 12864 -9209 12870 -9205
rect 12824 -9221 12870 -9209
rect 12972 -9209 12978 -9205
rect 13012 -9209 13018 -9205
rect 12972 -9221 13018 -9209
rect 13120 -9209 13126 -9205
rect 13160 -9209 13166 -9205
rect 13120 -9221 13166 -9209
rect 13268 -9209 13274 -9205
rect 13308 -9209 13314 -9205
rect 13268 -9221 13314 -9209
rect 13416 -9209 13422 -9205
rect 13456 -9209 13462 -9205
rect 13416 -9221 13462 -9209
rect 13564 -9209 13570 -9205
rect 13604 -9209 13610 -9205
rect 13564 -9221 13610 -9209
rect 13712 -9209 13718 -9205
rect 13752 -9209 13758 -9205
rect 13712 -9221 13758 -9209
rect 13860 -9209 13866 -9205
rect 13900 -9209 13906 -9205
rect 13860 -9221 13906 -9209
rect 14008 -9209 14014 -9205
rect 14048 -9209 14054 -9205
rect 14008 -9221 14054 -9209
rect 14156 -9209 14162 -9205
rect 14196 -9209 14202 -9205
rect 14156 -9221 14202 -9209
rect 14304 -9209 14310 -9205
rect 14344 -9209 14350 -9205
rect 14304 -9221 14350 -9209
rect 14452 -9209 14458 -9205
rect 14492 -9209 14498 -9205
rect 14452 -9221 14498 -9209
rect 14600 -9209 14606 -9205
rect 14640 -9209 14646 -9205
rect 14600 -9221 14646 -9209
rect 14748 -9209 14754 -9205
rect 14788 -9209 14794 -9205
rect 14748 -9221 14794 -9209
rect 14896 -9209 14902 -9205
rect 14936 -9209 14942 -9205
rect 14896 -9221 14942 -9209
rect 15044 -9209 15050 -9205
rect 15084 -9209 15090 -9205
rect 15044 -9221 15090 -9209
rect 15192 -9209 15198 -9205
rect 15232 -9209 15238 -9205
rect 15192 -9221 15238 -9209
rect 15340 -9209 15346 -9205
rect 15380 -9209 15386 -9205
rect 15340 -9221 15386 -9209
rect 15488 -9209 15494 -9205
rect 15528 -9209 15534 -9205
rect 15488 -9221 15534 -9209
rect 15636 -9209 15642 -9205
rect 15676 -9209 15682 -9205
rect 15636 -9221 15682 -9209
rect 15784 -9209 15790 -9205
rect 15824 -9209 15830 -9205
rect 15784 -9221 15830 -9209
rect 15932 -9209 15938 -9205
rect 15972 -9209 15978 -9205
rect 15932 -9221 15978 -9209
rect 16080 -9209 16086 -9205
rect 16120 -9209 16126 -9205
rect 16080 -9221 16126 -9209
rect 16228 -9209 16234 -9205
rect 16268 -9209 16274 -9205
rect 16228 -9221 16274 -9209
rect 16376 -9209 16382 -9205
rect 16416 -9209 16422 -9205
rect 16376 -9221 16422 -9209
rect 16524 -9209 16530 -9205
rect 16564 -9209 16570 -9205
rect 16524 -9221 16570 -9209
rect 16672 -9209 16678 -9205
rect 16712 -9209 16718 -9205
rect 16672 -9221 16718 -9209
rect 16820 -9209 16826 -9205
rect 16860 -9209 16866 -9205
rect 16820 -9221 16866 -9209
rect 16968 -9209 16974 -9205
rect 17008 -9209 17014 -9205
rect 16968 -9221 17014 -9209
rect 17116 -9209 17122 -9205
rect 17156 -9209 17162 -9205
rect 17116 -9221 17162 -9209
rect 17264 -9209 17270 -9205
rect 17304 -9209 17310 -9205
rect 17264 -9221 17310 -9209
rect 17412 -9209 17418 -9205
rect 17452 -9209 17458 -9205
rect 17412 -9221 17458 -9209
rect 17560 -9209 17566 -9205
rect 17600 -9209 17606 -9205
rect 17560 -9221 17606 -9209
rect 17708 -9209 17714 -9205
rect 17748 -9209 17754 -9205
rect 17708 -9221 17754 -9209
rect 17856 -9209 17862 -9205
rect 17896 -9209 17902 -9205
rect 17856 -9221 17902 -9209
rect 18004 -9209 18010 -9205
rect 18044 -9209 18050 -9205
rect 18004 -9221 18050 -9209
rect 18152 -9209 18158 -9205
rect 18192 -9209 18198 -9205
rect 18152 -9221 18198 -9209
rect 18300 -9209 18306 -9205
rect 18340 -9209 18346 -9205
rect 18300 -9221 18346 -9209
rect 18448 -9209 18454 -9205
rect 18488 -9209 18494 -9205
rect 18448 -9221 18494 -9209
rect 18596 -9209 18602 -9205
rect 18636 -9209 18642 -9205
rect 18596 -9221 18642 -9209
rect 18744 -9209 18750 -9205
rect 18784 -9209 18790 -9205
rect 18744 -9221 18790 -9209
rect 18892 -9209 18898 -9205
rect 18932 -9209 18938 -9205
rect 18892 -9221 18938 -9209
rect 19040 -9209 19046 -9205
rect 19080 -9209 19086 -9205
rect 19040 -9221 19086 -9209
rect 19188 -9209 19194 -9205
rect 19228 -9209 19234 -9205
rect 19188 -9221 19234 -9209
rect 19336 -9209 19342 -9205
rect 19376 -9209 19382 -9205
rect 19336 -9221 19382 -9209
rect 19484 -9209 19490 -9205
rect 19524 -9209 19530 -9205
rect 19484 -9221 19530 -9209
rect 19632 -9209 19638 -9205
rect 19672 -9209 19678 -9205
rect 19632 -9221 19678 -9209
rect 19780 -9209 19786 -9205
rect 19820 -9209 19826 -9205
rect 19780 -9221 19826 -9209
rect 19928 -9209 19934 -9205
rect 19968 -9209 19974 -9205
rect 19928 -9221 19974 -9209
rect 20076 -9209 20082 -9205
rect 20116 -9209 20122 -9205
rect 20076 -9221 20122 -9209
rect 20224 -9209 20230 -9205
rect 20264 -9209 20270 -9205
rect 20224 -9221 20270 -9209
rect 20372 -9209 20378 -9205
rect 20412 -9209 20418 -9205
rect 20372 -9221 20418 -9209
rect 20520 -9209 20526 -9205
rect 20560 -9209 20566 -9205
rect 20520 -9221 20566 -9209
rect 20668 -9209 20674 -9205
rect 20708 -9209 20714 -9205
rect 20668 -9221 20714 -9209
rect 20816 -9209 20822 -9205
rect 20856 -9209 20862 -9205
rect 20816 -9221 20862 -9209
rect 20964 -9209 20970 -9205
rect 21004 -9209 21010 -9205
rect 20964 -9221 21010 -9209
rect 21112 -9209 21118 -9205
rect 21152 -9209 21158 -9205
rect 21112 -9221 21158 -9209
rect 21260 -9209 21266 -9205
rect 21300 -9209 21306 -9205
rect 21260 -9221 21306 -9209
rect 21408 -9209 21414 -9205
rect 21448 -9209 21454 -9205
rect 21408 -9221 21454 -9209
rect 21556 -9209 21562 -9205
rect 21596 -9209 21602 -9205
rect 21556 -9221 21602 -9209
rect 21704 -9209 21710 -9205
rect 21744 -9209 21750 -9205
rect 21704 -9221 21750 -9209
rect 21852 -9209 21858 -9205
rect 21892 -9209 21898 -9205
rect 21852 -9221 21898 -9209
rect 22000 -9209 22006 -9205
rect 22040 -9209 22046 -9205
rect 22000 -9221 22046 -9209
rect 22148 -9209 22154 -9205
rect 22188 -9209 22194 -9205
rect 22148 -9221 22194 -9209
rect 22296 -9209 22302 -9205
rect 22336 -9209 22342 -9205
rect 22296 -9221 22342 -9209
rect 22444 -9209 22450 -9205
rect 22484 -9209 22490 -9205
rect 22444 -9221 22490 -9209
rect 22592 -9209 22598 -9205
rect 22632 -9209 22638 -9205
rect 22592 -9221 22638 -9209
rect 22740 -9209 22746 -9205
rect 22780 -9209 22786 -9205
rect 22740 -9221 22786 -9209
rect 22888 -9209 22894 -9205
rect 22928 -9209 22934 -9205
rect 22888 -9221 22934 -9209
rect 23036 -9209 23042 -9205
rect 23076 -9209 23082 -9205
rect 23036 -9221 23082 -9209
rect 23184 -9209 23190 -9205
rect 23224 -9209 23230 -9205
rect 23184 -9221 23230 -9209
rect 23332 -9209 23338 -9205
rect 23372 -9209 23378 -9205
rect 23332 -9221 23378 -9209
rect 4123 -9954 4126 -9658
rect 4197 -9954 4200 -9658
rect 4271 -9954 4274 -9658
rect 4345 -9683 4348 -9658
rect 4419 -9683 4422 -9658
rect 4493 -9683 4496 -9658
rect 4567 -9683 4570 -9658
rect 4641 -9683 4644 -9658
rect 4715 -9683 4718 -9658
rect 4789 -9683 4792 -9658
rect 4345 -9787 4348 -9735
rect 4419 -9787 4422 -9735
rect 4493 -9787 4496 -9735
rect 4567 -9787 4570 -9735
rect 4641 -9787 4644 -9735
rect 4715 -9787 4718 -9735
rect 4789 -9787 4792 -9735
rect 4345 -9891 4348 -9839
rect 4419 -9891 4422 -9839
rect 4493 -9891 4496 -9839
rect 4567 -9891 4570 -9839
rect 4641 -9891 4644 -9839
rect 4715 -9891 4718 -9839
rect 4789 -9891 4792 -9839
rect 4345 -9954 4348 -9943
rect 4419 -9954 4422 -9943
rect 4493 -9954 4496 -9943
rect 4567 -9954 4570 -9943
rect 4641 -9954 4644 -9943
rect 4715 -9954 4718 -9943
rect 4789 -9954 4792 -9943
rect 4863 -9954 4866 -9658
rect 4937 -9954 4940 -9658
rect 5011 -9954 5014 -9658
rect 5085 -9954 5088 -9658
rect 5159 -9683 5162 -9658
rect 5233 -9683 5236 -9658
rect 5307 -9683 5310 -9658
rect 5381 -9683 5384 -9658
rect 5455 -9683 5458 -9658
rect 5529 -9683 5532 -9658
rect 5603 -9683 5606 -9658
rect 5677 -9683 5680 -9658
rect 5161 -9735 5162 -9683
rect 5159 -9787 5162 -9735
rect 5233 -9787 5236 -9735
rect 5307 -9787 5310 -9735
rect 5381 -9787 5384 -9735
rect 5455 -9787 5458 -9735
rect 5529 -9787 5532 -9735
rect 5603 -9787 5606 -9735
rect 5677 -9787 5680 -9735
rect 5161 -9839 5162 -9787
rect 5159 -9891 5162 -9839
rect 5233 -9891 5236 -9839
rect 5307 -9891 5310 -9839
rect 5381 -9891 5384 -9839
rect 5455 -9891 5458 -9839
rect 5529 -9891 5532 -9839
rect 5603 -9891 5606 -9839
rect 5677 -9891 5680 -9839
rect 5161 -9943 5162 -9891
rect 5159 -9954 5162 -9943
rect 5233 -9954 5236 -9943
rect 5307 -9954 5310 -9943
rect 5381 -9954 5384 -9943
rect 5455 -9954 5458 -9943
rect 5529 -9954 5532 -9943
rect 5603 -9954 5606 -9943
rect 5677 -9954 5680 -9943
rect 5751 -9954 5754 -9658
rect 5825 -9954 5828 -9658
rect 5899 -9954 5902 -9658
rect 5973 -9954 5976 -9658
rect 6047 -9683 6050 -9658
rect 6121 -9683 6124 -9658
rect 6195 -9683 6198 -9658
rect 6269 -9683 6272 -9658
rect 6343 -9683 6346 -9658
rect 6417 -9683 6420 -9658
rect 6491 -9683 6494 -9658
rect 6047 -9787 6050 -9735
rect 6121 -9787 6124 -9735
rect 6195 -9787 6198 -9735
rect 6269 -9787 6272 -9735
rect 6343 -9787 6346 -9735
rect 6417 -9787 6420 -9735
rect 6491 -9787 6494 -9735
rect 6047 -9891 6050 -9839
rect 6121 -9891 6124 -9839
rect 6195 -9891 6198 -9839
rect 6269 -9891 6272 -9839
rect 6343 -9891 6346 -9839
rect 6417 -9891 6420 -9839
rect 6491 -9891 6494 -9839
rect 6047 -9954 6050 -9943
rect 6121 -9954 6124 -9943
rect 6195 -9954 6198 -9943
rect 6269 -9954 6272 -9943
rect 6343 -9954 6346 -9943
rect 6417 -9954 6420 -9943
rect 6491 -9954 6494 -9943
rect 6565 -9954 6568 -9658
rect 6639 -9954 6642 -9658
rect 6713 -9954 6716 -9658
rect 6787 -9954 6790 -9658
rect 6861 -9683 6864 -9658
rect 6935 -9683 6938 -9658
rect 7009 -9683 7012 -9658
rect 7083 -9683 7086 -9658
rect 7157 -9683 7160 -9658
rect 7231 -9683 7234 -9658
rect 7305 -9683 7308 -9658
rect 7379 -9683 7382 -9658
rect 7379 -9735 7381 -9683
rect 6861 -9787 6864 -9735
rect 6935 -9787 6938 -9735
rect 7009 -9787 7012 -9735
rect 7083 -9787 7086 -9735
rect 7157 -9787 7160 -9735
rect 7231 -9787 7234 -9735
rect 7305 -9787 7308 -9735
rect 7379 -9787 7382 -9735
rect 7379 -9839 7381 -9787
rect 6861 -9891 6864 -9839
rect 6935 -9891 6938 -9839
rect 7009 -9891 7012 -9839
rect 7083 -9891 7086 -9839
rect 7157 -9891 7160 -9839
rect 7231 -9891 7234 -9839
rect 7305 -9891 7308 -9839
rect 7379 -9891 7382 -9839
rect 7379 -9943 7381 -9891
rect 6861 -9954 6864 -9943
rect 6935 -9954 6938 -9943
rect 7009 -9954 7012 -9943
rect 7083 -9954 7086 -9943
rect 7157 -9954 7160 -9943
rect 7231 -9954 7234 -9943
rect 7305 -9954 7308 -9943
rect 7379 -9954 7382 -9943
rect 7453 -9954 7456 -9658
rect 7527 -9954 7530 -9658
rect 7601 -9954 7604 -9658
rect 7675 -9683 7678 -9658
rect 7749 -9683 7752 -9658
rect 7823 -9683 7826 -9658
rect 7897 -9683 7900 -9658
rect 7971 -9683 7974 -9658
rect 8045 -9683 8048 -9658
rect 8119 -9683 8122 -9658
rect 8193 -9683 8196 -9658
rect 7677 -9735 7678 -9683
rect 7675 -9787 7678 -9735
rect 7749 -9787 7752 -9735
rect 7823 -9787 7826 -9735
rect 7897 -9787 7900 -9735
rect 7971 -9787 7974 -9735
rect 8045 -9787 8048 -9735
rect 8119 -9787 8122 -9735
rect 8193 -9787 8196 -9735
rect 7677 -9839 7678 -9787
rect 7675 -9891 7678 -9839
rect 7749 -9891 7752 -9839
rect 7823 -9891 7826 -9839
rect 7897 -9891 7900 -9839
rect 7971 -9891 7974 -9839
rect 8045 -9891 8048 -9839
rect 8119 -9891 8122 -9839
rect 8193 -9891 8196 -9839
rect 7677 -9943 7678 -9891
rect 7675 -9954 7678 -9943
rect 7749 -9954 7752 -9943
rect 7823 -9954 7826 -9943
rect 7897 -9954 7900 -9943
rect 7971 -9954 7974 -9943
rect 8045 -9954 8048 -9943
rect 8119 -9954 8122 -9943
rect 8193 -9954 8196 -9943
rect 8267 -9954 8270 -9658
rect 8341 -9954 8344 -9658
rect 8415 -9954 8418 -9658
rect 8489 -9954 8492 -9658
rect 8563 -9683 8566 -9658
rect 8637 -9683 8640 -9658
rect 8711 -9683 8714 -9658
rect 8785 -9683 8788 -9658
rect 8859 -9683 8862 -9658
rect 8933 -9683 8936 -9658
rect 9007 -9683 9010 -9658
rect 8563 -9787 8566 -9735
rect 8637 -9787 8640 -9735
rect 8711 -9787 8714 -9735
rect 8785 -9787 8788 -9735
rect 8859 -9787 8862 -9735
rect 8933 -9787 8936 -9735
rect 9007 -9787 9010 -9735
rect 8563 -9891 8566 -9839
rect 8637 -9891 8640 -9839
rect 8711 -9891 8714 -9839
rect 8785 -9891 8788 -9839
rect 8859 -9891 8862 -9839
rect 8933 -9891 8936 -9839
rect 9007 -9891 9010 -9839
rect 8563 -9954 8566 -9943
rect 8637 -9954 8640 -9943
rect 8711 -9954 8714 -9943
rect 8785 -9954 8788 -9943
rect 8859 -9954 8862 -9943
rect 8933 -9954 8936 -9943
rect 9007 -9954 9010 -9943
rect 9081 -9954 9084 -9658
rect 9155 -9954 9158 -9658
rect 9229 -9954 9232 -9658
rect 9303 -9954 9306 -9658
rect 9377 -9683 9380 -9658
rect 9451 -9683 9454 -9658
rect 9525 -9683 9528 -9658
rect 9599 -9683 9602 -9658
rect 9673 -9683 9676 -9658
rect 9747 -9683 9750 -9658
rect 9821 -9683 9824 -9658
rect 9895 -9683 9898 -9658
rect 9895 -9735 9897 -9683
rect 9377 -9787 9380 -9735
rect 9451 -9787 9454 -9735
rect 9525 -9787 9528 -9735
rect 9599 -9787 9602 -9735
rect 9673 -9787 9676 -9735
rect 9747 -9787 9750 -9735
rect 9821 -9787 9824 -9735
rect 9895 -9787 9898 -9735
rect 9895 -9839 9897 -9787
rect 9377 -9891 9380 -9839
rect 9451 -9891 9454 -9839
rect 9525 -9891 9528 -9839
rect 9599 -9891 9602 -9839
rect 9673 -9891 9676 -9839
rect 9747 -9891 9750 -9839
rect 9821 -9891 9824 -9839
rect 9895 -9891 9898 -9839
rect 9895 -9943 9897 -9891
rect 9377 -9954 9380 -9943
rect 9451 -9954 9454 -9943
rect 9525 -9954 9528 -9943
rect 9599 -9954 9602 -9943
rect 9673 -9954 9676 -9943
rect 9747 -9954 9750 -9943
rect 9821 -9954 9824 -9943
rect 9895 -9954 9898 -9943
rect 9969 -9954 9972 -9658
rect 10043 -9954 10046 -9658
rect 10117 -9954 10120 -9658
rect 10191 -9683 10194 -9658
rect 10265 -9683 10268 -9658
rect 10339 -9683 10342 -9658
rect 10413 -9683 10416 -9658
rect 10487 -9683 10490 -9658
rect 10561 -9683 10564 -9658
rect 10635 -9683 10638 -9658
rect 10709 -9683 10712 -9658
rect 10192 -9735 10194 -9683
rect 10191 -9787 10194 -9735
rect 10265 -9787 10268 -9735
rect 10339 -9787 10342 -9735
rect 10413 -9787 10416 -9735
rect 10487 -9787 10490 -9735
rect 10561 -9787 10564 -9735
rect 10635 -9787 10638 -9735
rect 10709 -9787 10712 -9735
rect 10192 -9839 10194 -9787
rect 10191 -9891 10194 -9839
rect 10265 -9891 10268 -9839
rect 10339 -9891 10342 -9839
rect 10413 -9891 10416 -9839
rect 10487 -9891 10490 -9839
rect 10561 -9891 10564 -9839
rect 10635 -9891 10638 -9839
rect 10709 -9891 10712 -9839
rect 10192 -9943 10194 -9891
rect 10191 -9954 10194 -9943
rect 10265 -9954 10268 -9943
rect 10339 -9954 10342 -9943
rect 10413 -9954 10416 -9943
rect 10487 -9954 10490 -9943
rect 10561 -9954 10564 -9943
rect 10635 -9954 10638 -9943
rect 10709 -9954 10712 -9943
rect 10783 -9954 10786 -9658
rect 10857 -9954 10860 -9658
rect 10931 -9954 10934 -9658
rect 11005 -9954 11008 -9658
rect 11079 -9683 11082 -9658
rect 11153 -9683 11156 -9658
rect 11227 -9683 11230 -9658
rect 11301 -9683 11304 -9658
rect 11375 -9683 11378 -9658
rect 11449 -9683 11452 -9658
rect 11523 -9683 11526 -9658
rect 11079 -9787 11082 -9735
rect 11153 -9787 11156 -9735
rect 11227 -9787 11230 -9735
rect 11301 -9787 11304 -9735
rect 11375 -9787 11378 -9735
rect 11449 -9787 11452 -9735
rect 11523 -9787 11526 -9735
rect 11079 -9891 11082 -9839
rect 11153 -9891 11156 -9839
rect 11227 -9891 11230 -9839
rect 11301 -9891 11304 -9839
rect 11375 -9891 11378 -9839
rect 11449 -9891 11452 -9839
rect 11523 -9891 11526 -9839
rect 11079 -9954 11082 -9943
rect 11153 -9954 11156 -9943
rect 11227 -9954 11230 -9943
rect 11301 -9954 11304 -9943
rect 11375 -9954 11378 -9943
rect 11449 -9954 11452 -9943
rect 11523 -9954 11526 -9943
rect 11597 -9954 11600 -9658
rect 11671 -9954 11674 -9658
rect 11745 -9954 11748 -9658
rect 11819 -9954 11822 -9658
rect 11893 -9683 11896 -9658
rect 11967 -9683 11970 -9658
rect 12041 -9683 12044 -9658
rect 12115 -9683 12118 -9658
rect 12189 -9683 12192 -9658
rect 12263 -9683 12266 -9658
rect 12337 -9683 12340 -9658
rect 12411 -9683 12414 -9658
rect 12411 -9735 12412 -9683
rect 11893 -9787 11896 -9735
rect 11967 -9787 11970 -9735
rect 12041 -9787 12044 -9735
rect 12115 -9787 12118 -9735
rect 12189 -9787 12192 -9735
rect 12263 -9787 12266 -9735
rect 12337 -9787 12340 -9735
rect 12411 -9787 12414 -9735
rect 12411 -9839 12412 -9787
rect 11893 -9891 11896 -9839
rect 11967 -9891 11970 -9839
rect 12041 -9891 12044 -9839
rect 12115 -9891 12118 -9839
rect 12189 -9891 12192 -9839
rect 12263 -9891 12266 -9839
rect 12337 -9891 12340 -9839
rect 12411 -9891 12414 -9839
rect 12411 -9943 12412 -9891
rect 11893 -9954 11896 -9943
rect 11967 -9954 11970 -9943
rect 12041 -9954 12044 -9943
rect 12115 -9954 12118 -9943
rect 12189 -9954 12192 -9943
rect 12263 -9954 12266 -9943
rect 12337 -9954 12340 -9943
rect 12411 -9954 12414 -9943
rect 12485 -9954 12488 -9658
rect 12559 -9954 12562 -9658
rect 12633 -9954 12636 -9658
rect 12707 -9683 12710 -9658
rect 12781 -9683 12784 -9658
rect 12855 -9683 12858 -9658
rect 12929 -9683 12932 -9658
rect 13003 -9683 13006 -9658
rect 13077 -9683 13080 -9658
rect 13151 -9683 13154 -9658
rect 13225 -9683 13228 -9658
rect 12708 -9735 12710 -9683
rect 12707 -9787 12710 -9735
rect 12781 -9787 12784 -9735
rect 12855 -9787 12858 -9735
rect 12929 -9787 12932 -9735
rect 13003 -9787 13006 -9735
rect 13077 -9787 13080 -9735
rect 13151 -9787 13154 -9735
rect 13225 -9787 13228 -9735
rect 12708 -9839 12710 -9787
rect 12707 -9891 12710 -9839
rect 12781 -9891 12784 -9839
rect 12855 -9891 12858 -9839
rect 12929 -9891 12932 -9839
rect 13003 -9891 13006 -9839
rect 13077 -9891 13080 -9839
rect 13151 -9891 13154 -9839
rect 13225 -9891 13228 -9839
rect 12708 -9943 12710 -9891
rect 12707 -9954 12710 -9943
rect 12781 -9954 12784 -9943
rect 12855 -9954 12858 -9943
rect 12929 -9954 12932 -9943
rect 13003 -9954 13006 -9943
rect 13077 -9954 13080 -9943
rect 13151 -9954 13154 -9943
rect 13225 -9954 13228 -9943
rect 13299 -9954 13302 -9658
rect 13373 -9954 13376 -9658
rect 13447 -9954 13450 -9658
rect 13521 -9954 13524 -9658
rect 13595 -9683 13598 -9658
rect 13669 -9683 13672 -9658
rect 13743 -9683 13746 -9658
rect 13817 -9683 13820 -9658
rect 13891 -9683 13894 -9658
rect 13965 -9683 13968 -9658
rect 14039 -9683 14042 -9658
rect 13595 -9787 13598 -9735
rect 13669 -9787 13672 -9735
rect 13743 -9787 13746 -9735
rect 13817 -9787 13820 -9735
rect 13891 -9787 13894 -9735
rect 13965 -9787 13968 -9735
rect 14039 -9787 14042 -9735
rect 13595 -9891 13598 -9839
rect 13669 -9891 13672 -9839
rect 13743 -9891 13746 -9839
rect 13817 -9891 13820 -9839
rect 13891 -9891 13894 -9839
rect 13965 -9891 13968 -9839
rect 14039 -9891 14042 -9839
rect 13595 -9954 13598 -9943
rect 13669 -9954 13672 -9943
rect 13743 -9954 13746 -9943
rect 13817 -9954 13820 -9943
rect 13891 -9954 13894 -9943
rect 13965 -9954 13968 -9943
rect 14039 -9954 14042 -9943
rect 14113 -9954 14116 -9658
rect 14187 -9954 14190 -9658
rect 14261 -9954 14264 -9658
rect 14335 -9954 14338 -9658
rect 14409 -9683 14412 -9658
rect 14483 -9683 14486 -9658
rect 14557 -9683 14560 -9658
rect 14631 -9683 14634 -9658
rect 14705 -9683 14708 -9658
rect 14779 -9683 14782 -9658
rect 14853 -9683 14856 -9658
rect 14927 -9683 14930 -9658
rect 14927 -9735 14928 -9683
rect 14409 -9787 14412 -9735
rect 14483 -9787 14486 -9735
rect 14557 -9787 14560 -9735
rect 14631 -9787 14634 -9735
rect 14705 -9787 14708 -9735
rect 14779 -9787 14782 -9735
rect 14853 -9787 14856 -9735
rect 14927 -9787 14930 -9735
rect 14927 -9839 14928 -9787
rect 14409 -9891 14412 -9839
rect 14483 -9891 14486 -9839
rect 14557 -9891 14560 -9839
rect 14631 -9891 14634 -9839
rect 14705 -9891 14708 -9839
rect 14779 -9891 14782 -9839
rect 14853 -9891 14856 -9839
rect 14927 -9891 14930 -9839
rect 14927 -9943 14928 -9891
rect 14409 -9954 14412 -9943
rect 14483 -9954 14486 -9943
rect 14557 -9954 14560 -9943
rect 14631 -9954 14634 -9943
rect 14705 -9954 14708 -9943
rect 14779 -9954 14782 -9943
rect 14853 -9954 14856 -9943
rect 14927 -9954 14930 -9943
rect 15001 -9954 15004 -9658
rect 15075 -9954 15078 -9658
rect 15149 -9954 15152 -9658
rect 15223 -9954 15226 -9658
rect 15297 -9683 15300 -9658
rect 15371 -9683 15374 -9658
rect 15445 -9683 15448 -9658
rect 15519 -9683 15522 -9658
rect 15593 -9683 15596 -9658
rect 15667 -9683 15670 -9658
rect 15741 -9683 15744 -9658
rect 15297 -9787 15300 -9735
rect 15371 -9787 15374 -9735
rect 15445 -9787 15448 -9735
rect 15519 -9787 15522 -9735
rect 15593 -9787 15596 -9735
rect 15667 -9787 15670 -9735
rect 15741 -9787 15744 -9735
rect 15297 -9891 15300 -9839
rect 15371 -9891 15374 -9839
rect 15445 -9891 15448 -9839
rect 15519 -9891 15522 -9839
rect 15593 -9891 15596 -9839
rect 15667 -9891 15670 -9839
rect 15741 -9891 15744 -9839
rect 15297 -9954 15300 -9943
rect 15371 -9954 15374 -9943
rect 15445 -9954 15448 -9943
rect 15519 -9954 15522 -9943
rect 15593 -9954 15596 -9943
rect 15667 -9954 15670 -9943
rect 15741 -9954 15744 -9943
rect 15815 -9954 15818 -9658
rect 15889 -9954 15892 -9658
rect 15963 -9954 15966 -9658
rect 16037 -9954 16040 -9658
rect 16111 -9683 16114 -9658
rect 16185 -9683 16188 -9658
rect 16259 -9683 16262 -9658
rect 16333 -9683 16336 -9658
rect 16407 -9683 16410 -9658
rect 16481 -9683 16484 -9658
rect 16555 -9683 16558 -9658
rect 16111 -9787 16114 -9735
rect 16185 -9787 16188 -9735
rect 16259 -9787 16262 -9735
rect 16333 -9787 16336 -9735
rect 16407 -9787 16410 -9735
rect 16481 -9787 16484 -9735
rect 16555 -9787 16558 -9735
rect 16111 -9891 16114 -9839
rect 16185 -9891 16188 -9839
rect 16259 -9891 16262 -9839
rect 16333 -9891 16336 -9839
rect 16407 -9891 16410 -9839
rect 16481 -9891 16484 -9839
rect 16555 -9891 16558 -9839
rect 16111 -9954 16114 -9943
rect 16185 -9954 16188 -9943
rect 16259 -9954 16262 -9943
rect 16333 -9954 16336 -9943
rect 16407 -9954 16410 -9943
rect 16481 -9954 16484 -9943
rect 16555 -9954 16558 -9943
rect 16629 -9954 16632 -9658
rect 16703 -9954 16706 -9658
rect 16777 -9954 16780 -9658
rect 16851 -9954 16854 -9658
rect 16925 -9683 16928 -9658
rect 16999 -9683 17002 -9658
rect 17073 -9683 17076 -9658
rect 17147 -9683 17150 -9658
rect 17221 -9683 17224 -9658
rect 17295 -9683 17298 -9658
rect 17369 -9683 17372 -9658
rect 17443 -9683 17446 -9658
rect 16927 -9735 16928 -9683
rect 16925 -9787 16928 -9735
rect 16999 -9787 17002 -9735
rect 17073 -9787 17076 -9735
rect 17147 -9787 17150 -9735
rect 17221 -9787 17224 -9735
rect 17295 -9787 17298 -9735
rect 17369 -9787 17372 -9735
rect 17443 -9787 17446 -9735
rect 16927 -9839 16928 -9787
rect 16925 -9891 16928 -9839
rect 16999 -9891 17002 -9839
rect 17073 -9891 17076 -9839
rect 17147 -9891 17150 -9839
rect 17221 -9891 17224 -9839
rect 17295 -9891 17298 -9839
rect 17369 -9891 17372 -9839
rect 17443 -9891 17446 -9839
rect 16927 -9943 16928 -9891
rect 16925 -9954 16928 -9943
rect 16999 -9954 17002 -9943
rect 17073 -9954 17076 -9943
rect 17147 -9954 17150 -9943
rect 17221 -9954 17224 -9943
rect 17295 -9954 17298 -9943
rect 17369 -9954 17372 -9943
rect 17443 -9954 17446 -9943
rect 17517 -9954 17520 -9658
rect 17591 -9954 17594 -9658
rect 17665 -9954 17668 -9658
rect 17739 -9954 17742 -9658
rect 17813 -9683 17816 -9658
rect 17887 -9683 17890 -9658
rect 17961 -9683 17964 -9658
rect 18035 -9683 18038 -9658
rect 18109 -9683 18112 -9658
rect 18183 -9683 18186 -9658
rect 18257 -9683 18260 -9658
rect 17813 -9787 17816 -9735
rect 17887 -9787 17890 -9735
rect 17961 -9787 17964 -9735
rect 18035 -9787 18038 -9735
rect 18109 -9787 18112 -9735
rect 18183 -9787 18186 -9735
rect 18257 -9787 18260 -9735
rect 17813 -9891 17816 -9839
rect 17887 -9891 17890 -9839
rect 17961 -9891 17964 -9839
rect 18035 -9891 18038 -9839
rect 18109 -9891 18112 -9839
rect 18183 -9891 18186 -9839
rect 18257 -9891 18260 -9839
rect 17813 -9954 17816 -9943
rect 17887 -9954 17890 -9943
rect 17961 -9954 17964 -9943
rect 18035 -9954 18038 -9943
rect 18109 -9954 18112 -9943
rect 18183 -9954 18186 -9943
rect 18257 -9954 18260 -9943
rect 18331 -9954 18334 -9658
rect 18405 -9954 18408 -9658
rect 18479 -9954 18482 -9658
rect 18553 -9954 18556 -9658
rect 18627 -9683 18630 -9658
rect 18701 -9683 18704 -9658
rect 18775 -9683 18778 -9658
rect 18849 -9683 18852 -9658
rect 18923 -9683 18926 -9658
rect 18997 -9683 19000 -9658
rect 19071 -9683 19074 -9658
rect 19145 -9683 19148 -9658
rect 19145 -9735 19146 -9683
rect 18627 -9787 18630 -9735
rect 18701 -9787 18704 -9735
rect 18775 -9787 18778 -9735
rect 18849 -9787 18852 -9735
rect 18923 -9787 18926 -9735
rect 18997 -9787 19000 -9735
rect 19071 -9787 19074 -9735
rect 19145 -9787 19148 -9735
rect 19145 -9839 19146 -9787
rect 18627 -9891 18630 -9839
rect 18701 -9891 18704 -9839
rect 18775 -9891 18778 -9839
rect 18849 -9891 18852 -9839
rect 18923 -9891 18926 -9839
rect 18997 -9891 19000 -9839
rect 19071 -9891 19074 -9839
rect 19145 -9891 19148 -9839
rect 19145 -9943 19146 -9891
rect 18627 -9954 18630 -9943
rect 18701 -9954 18704 -9943
rect 18775 -9954 18778 -9943
rect 18849 -9954 18852 -9943
rect 18923 -9954 18926 -9943
rect 18997 -9954 19000 -9943
rect 19071 -9954 19074 -9943
rect 19145 -9954 19148 -9943
rect 19219 -9954 19222 -9658
rect 19293 -9954 19296 -9658
rect 19367 -9954 19370 -9658
rect 19441 -9683 19444 -9658
rect 19515 -9683 19518 -9658
rect 19589 -9683 19592 -9658
rect 19663 -9683 19666 -9658
rect 19737 -9683 19740 -9658
rect 19811 -9683 19814 -9658
rect 19885 -9683 19888 -9658
rect 19959 -9683 19962 -9658
rect 19442 -9735 19444 -9683
rect 19441 -9787 19444 -9735
rect 19515 -9787 19518 -9735
rect 19589 -9787 19592 -9735
rect 19663 -9787 19666 -9735
rect 19737 -9787 19740 -9735
rect 19811 -9787 19814 -9735
rect 19885 -9787 19888 -9735
rect 19959 -9787 19962 -9735
rect 19442 -9839 19444 -9787
rect 19441 -9891 19444 -9839
rect 19515 -9891 19518 -9839
rect 19589 -9891 19592 -9839
rect 19663 -9891 19666 -9839
rect 19737 -9891 19740 -9839
rect 19811 -9891 19814 -9839
rect 19885 -9891 19888 -9839
rect 19959 -9891 19962 -9839
rect 19442 -9943 19444 -9891
rect 19441 -9954 19444 -9943
rect 19515 -9954 19518 -9943
rect 19589 -9954 19592 -9943
rect 19663 -9954 19666 -9943
rect 19737 -9954 19740 -9943
rect 19811 -9954 19814 -9943
rect 19885 -9954 19888 -9943
rect 19959 -9954 19962 -9943
rect 20033 -9954 20036 -9658
rect 20107 -9954 20110 -9658
rect 20181 -9954 20184 -9658
rect 20255 -9954 20258 -9658
rect 20329 -9683 20332 -9658
rect 20403 -9683 20406 -9658
rect 20477 -9683 20480 -9658
rect 20551 -9683 20554 -9658
rect 20625 -9683 20628 -9658
rect 20699 -9683 20702 -9658
rect 20773 -9683 20776 -9658
rect 20329 -9787 20332 -9735
rect 20403 -9787 20406 -9735
rect 20477 -9787 20480 -9735
rect 20551 -9787 20554 -9735
rect 20625 -9787 20628 -9735
rect 20699 -9787 20702 -9735
rect 20773 -9787 20776 -9735
rect 20329 -9891 20332 -9839
rect 20403 -9891 20406 -9839
rect 20477 -9891 20480 -9839
rect 20551 -9891 20554 -9839
rect 20625 -9891 20628 -9839
rect 20699 -9891 20702 -9839
rect 20773 -9891 20776 -9839
rect 20329 -9954 20332 -9943
rect 20403 -9954 20406 -9943
rect 20477 -9954 20480 -9943
rect 20551 -9954 20554 -9943
rect 20625 -9954 20628 -9943
rect 20699 -9954 20702 -9943
rect 20773 -9954 20776 -9943
rect 20847 -9954 20850 -9658
rect 20921 -9954 20924 -9658
rect 20995 -9954 20998 -9658
rect 21069 -9954 21072 -9658
rect 21143 -9683 21146 -9658
rect 21217 -9683 21220 -9658
rect 21291 -9683 21294 -9658
rect 21365 -9683 21368 -9658
rect 21439 -9683 21442 -9658
rect 21513 -9683 21516 -9658
rect 21587 -9683 21590 -9658
rect 21661 -9683 21664 -9658
rect 21661 -9735 21662 -9683
rect 21143 -9787 21146 -9735
rect 21217 -9787 21220 -9735
rect 21291 -9787 21294 -9735
rect 21365 -9787 21368 -9735
rect 21439 -9787 21442 -9735
rect 21513 -9787 21516 -9735
rect 21587 -9787 21590 -9735
rect 21661 -9787 21664 -9735
rect 21661 -9839 21662 -9787
rect 21143 -9891 21146 -9839
rect 21217 -9891 21220 -9839
rect 21291 -9891 21294 -9839
rect 21365 -9891 21368 -9839
rect 21439 -9891 21442 -9839
rect 21513 -9891 21516 -9839
rect 21587 -9891 21590 -9839
rect 21661 -9891 21664 -9839
rect 21661 -9943 21662 -9891
rect 21143 -9954 21146 -9943
rect 21217 -9954 21220 -9943
rect 21291 -9954 21294 -9943
rect 21365 -9954 21368 -9943
rect 21439 -9954 21442 -9943
rect 21513 -9954 21516 -9943
rect 21587 -9954 21590 -9943
rect 21661 -9954 21664 -9943
rect 21735 -9954 21738 -9658
rect 21809 -9954 21812 -9658
rect 21883 -9954 21886 -9658
rect 21957 -9954 21960 -9658
rect 22031 -9683 22034 -9658
rect 22105 -9683 22108 -9658
rect 22179 -9683 22182 -9658
rect 22253 -9683 22256 -9658
rect 22327 -9683 22330 -9658
rect 22401 -9683 22404 -9658
rect 22475 -9683 22478 -9658
rect 22031 -9787 22034 -9735
rect 22105 -9787 22108 -9735
rect 22179 -9787 22182 -9735
rect 22253 -9787 22256 -9735
rect 22327 -9787 22330 -9735
rect 22401 -9787 22404 -9735
rect 22475 -9787 22478 -9735
rect 22031 -9891 22034 -9839
rect 22105 -9891 22108 -9839
rect 22179 -9891 22182 -9839
rect 22253 -9891 22256 -9839
rect 22327 -9891 22330 -9839
rect 22401 -9891 22404 -9839
rect 22475 -9891 22478 -9839
rect 22031 -9954 22034 -9943
rect 22105 -9954 22108 -9943
rect 22179 -9954 22182 -9943
rect 22253 -9954 22256 -9943
rect 22327 -9954 22330 -9943
rect 22401 -9954 22404 -9943
rect 22475 -9954 22478 -9943
rect 22549 -9954 22552 -9658
rect 22623 -9954 22626 -9658
rect 22697 -9954 22700 -9658
rect 22771 -9954 22774 -9658
rect 22845 -9683 22848 -9658
rect 22919 -9683 22922 -9658
rect 22993 -9683 22996 -9658
rect 23067 -9683 23070 -9658
rect 23141 -9683 23144 -9658
rect 23215 -9683 23218 -9658
rect 23289 -9683 23292 -9658
rect 22845 -9787 22848 -9735
rect 22919 -9787 22922 -9735
rect 22993 -9787 22996 -9735
rect 23067 -9787 23070 -9735
rect 23141 -9787 23144 -9735
rect 23215 -9787 23218 -9735
rect 23289 -9787 23292 -9735
rect 22845 -9891 22848 -9839
rect 22919 -9891 22922 -9839
rect 22993 -9891 22996 -9839
rect 23067 -9891 23070 -9839
rect 23141 -9891 23144 -9839
rect 23215 -9891 23218 -9839
rect 23289 -9891 23292 -9839
rect 22845 -9954 22848 -9943
rect 22919 -9954 22922 -9943
rect 22993 -9954 22996 -9943
rect 23067 -9954 23070 -9943
rect 23141 -9954 23144 -9943
rect 23215 -9954 23218 -9943
rect 23289 -9954 23292 -9943
rect 23363 -9954 23366 -9658
rect 23437 -9954 23440 -9658
rect 23511 -9954 23514 -9658
rect 23585 -9954 23588 -9658
rect 23659 -9683 23662 -9658
rect 23733 -9683 23736 -9658
rect 23807 -9683 23810 -9658
rect 23881 -9683 23884 -9658
rect 23955 -9683 23958 -9658
rect 24029 -9683 24032 -9658
rect 24103 -9683 24106 -9658
rect 24177 -9683 24180 -9658
rect 23661 -9735 23662 -9683
rect 23659 -9787 23662 -9735
rect 23733 -9787 23736 -9735
rect 23807 -9787 23810 -9735
rect 23881 -9787 23884 -9735
rect 23955 -9787 23958 -9735
rect 24029 -9787 24032 -9735
rect 24103 -9787 24106 -9735
rect 24177 -9787 24180 -9735
rect 23661 -9839 23662 -9787
rect 23659 -9891 23662 -9839
rect 23733 -9891 23736 -9839
rect 23807 -9891 23810 -9839
rect 23881 -9891 23884 -9839
rect 23955 -9891 23958 -9839
rect 24029 -9891 24032 -9839
rect 24103 -9891 24106 -9839
rect 24177 -9891 24180 -9839
rect 23661 -9943 23662 -9891
rect 23659 -9954 23662 -9943
rect 23733 -9954 23736 -9943
rect 23807 -9954 23810 -9943
rect 23881 -9954 23884 -9943
rect 23955 -9954 23958 -9943
rect 24029 -9954 24032 -9943
rect 24103 -9954 24106 -9943
rect 24177 -9954 24180 -9943
rect 24251 -9954 24254 -9658
rect 24325 -9954 24328 -9658
rect 24399 -9954 24402 -9658
rect 24473 -9954 24476 -9658
rect 24547 -9683 24550 -9658
rect 24621 -9683 24624 -9658
rect 24695 -9683 24698 -9658
rect 24769 -9683 24772 -9658
rect 24843 -9683 24846 -9658
rect 24917 -9683 24920 -9658
rect 24991 -9683 24994 -9658
rect 24547 -9787 24550 -9735
rect 24621 -9787 24624 -9735
rect 24695 -9787 24698 -9735
rect 24769 -9787 24772 -9735
rect 24843 -9787 24846 -9735
rect 24917 -9787 24920 -9735
rect 24991 -9787 24994 -9735
rect 24547 -9891 24550 -9839
rect 24621 -9891 24624 -9839
rect 24695 -9891 24698 -9839
rect 24769 -9891 24772 -9839
rect 24843 -9891 24846 -9839
rect 24917 -9891 24920 -9839
rect 24991 -9891 24994 -9839
rect 24547 -9954 24550 -9943
rect 24621 -9954 24624 -9943
rect 24695 -9954 24698 -9943
rect 24769 -9954 24772 -9943
rect 24843 -9954 24846 -9943
rect 24917 -9954 24920 -9943
rect 24991 -9954 24994 -9943
rect 25065 -9954 25068 -9658
rect 25139 -9954 25142 -9658
rect 25213 -9954 25216 -9658
rect 25287 -9954 25290 -9658
rect 25361 -9683 25364 -9658
rect 25435 -9683 25438 -9658
rect 25509 -9683 25512 -9658
rect 25583 -9683 25586 -9658
rect 25657 -9683 25660 -9658
rect 25731 -9683 25734 -9658
rect 25805 -9683 25808 -9658
rect 25879 -9683 25882 -9658
rect 25879 -9735 25881 -9683
rect 25361 -9787 25364 -9735
rect 25435 -9787 25438 -9735
rect 25509 -9787 25512 -9735
rect 25583 -9787 25586 -9735
rect 25657 -9787 25660 -9735
rect 25731 -9787 25734 -9735
rect 25805 -9787 25808 -9735
rect 25879 -9787 25882 -9735
rect 25879 -9839 25881 -9787
rect 25361 -9891 25364 -9839
rect 25435 -9891 25438 -9839
rect 25509 -9891 25512 -9839
rect 25583 -9891 25586 -9839
rect 25657 -9891 25660 -9839
rect 25731 -9891 25734 -9839
rect 25805 -9891 25808 -9839
rect 25879 -9891 25882 -9839
rect 25879 -9943 25881 -9891
rect 25361 -9954 25364 -9943
rect 25435 -9954 25438 -9943
rect 25509 -9954 25512 -9943
rect 25583 -9954 25586 -9943
rect 25657 -9954 25660 -9943
rect 25731 -9954 25734 -9943
rect 25805 -9954 25808 -9943
rect 25879 -9954 25882 -9943
rect 25953 -9954 25956 -9658
rect 26027 -9954 26030 -9658
rect 26101 -9954 26104 -9658
rect 26175 -9683 26178 -9658
rect 26249 -9683 26258 -9658
rect 26177 -9735 26178 -9683
rect 26175 -9787 26178 -9735
rect 26249 -9787 26258 -9735
rect 26177 -9839 26178 -9787
rect 26175 -9891 26178 -9839
rect 26249 -9891 26258 -9839
rect 26177 -9943 26178 -9891
rect 26175 -9954 26178 -9943
rect 26249 -9952 26258 -9943
rect 26247 -9954 26258 -9952
<< via1 >>
rect 3038 3120 3090 3172
rect 3120 3120 3172 3172
rect 3201 3120 3253 3172
rect 3282 3120 3334 3172
rect 3363 3120 3415 3172
rect 3444 3120 3496 3172
rect 3525 3120 3577 3172
rect 3606 3120 3658 3172
rect 3688 3120 3740 3172
rect 3769 3120 3821 3172
rect 3850 3120 3902 3172
rect 3931 3120 3983 3172
rect 4012 3120 4064 3172
rect 4093 3120 4145 3172
rect 4174 3120 4226 3172
rect 4256 3120 4308 3172
rect 4337 3120 4389 3172
rect 4418 3120 4470 3172
rect 4499 3120 4551 3172
rect 4580 3120 4632 3172
rect 4661 3120 4713 3172
rect 4742 3152 4794 3172
rect 4824 3152 4876 3172
rect 4742 3120 4768 3152
rect 4768 3120 4794 3152
rect 4824 3120 4840 3152
rect 4840 3120 4874 3152
rect 4874 3120 4876 3152
rect 4905 3152 4957 3172
rect 4986 3152 5038 3172
rect 5067 3152 5119 3172
rect 5148 3152 5200 3172
rect 5229 3152 5281 3172
rect 5310 3152 5362 3172
rect 5392 3152 5444 3172
rect 5473 3152 5525 3172
rect 4905 3120 4912 3152
rect 4912 3120 4946 3152
rect 4946 3120 4957 3152
rect 4986 3120 5018 3152
rect 5018 3120 5038 3152
rect 5067 3120 5090 3152
rect 5090 3120 5119 3152
rect 5148 3120 5162 3152
rect 5162 3120 5200 3152
rect 5229 3120 5234 3152
rect 5234 3120 5272 3152
rect 5272 3120 5281 3152
rect 5310 3120 5344 3152
rect 5344 3120 5362 3152
rect 5392 3120 5416 3152
rect 5416 3120 5444 3152
rect 5473 3120 5488 3152
rect 5488 3120 5522 3152
rect 5522 3120 5525 3152
rect 5554 3152 5606 3172
rect 5635 3152 5687 3172
rect 5716 3152 5768 3172
rect 5797 3152 5849 3172
rect 5878 3152 5930 3172
rect 5960 3152 6012 3172
rect 6041 3152 6093 3172
rect 6122 3152 6174 3172
rect 5554 3120 5560 3152
rect 5560 3120 5594 3152
rect 5594 3120 5606 3152
rect 5635 3120 5666 3152
rect 5666 3120 5687 3152
rect 5716 3120 5738 3152
rect 5738 3120 5768 3152
rect 5797 3120 5810 3152
rect 5810 3120 5848 3152
rect 5848 3120 5849 3152
rect 5878 3120 5882 3152
rect 5882 3120 5920 3152
rect 5920 3120 5930 3152
rect 5960 3120 5992 3152
rect 5992 3120 6012 3152
rect 6041 3120 6064 3152
rect 6064 3120 6093 3152
rect 6122 3120 6136 3152
rect 6136 3120 6170 3152
rect 6170 3120 6174 3152
rect 6203 3152 6255 3172
rect 6284 3152 6336 3172
rect 6365 3152 6417 3172
rect 6446 3152 6498 3172
rect 6528 3152 6580 3172
rect 6609 3152 6661 3172
rect 6690 3152 6742 3172
rect 6771 3152 6823 3172
rect 6203 3120 6208 3152
rect 6208 3120 6242 3152
rect 6242 3120 6255 3152
rect 6284 3120 6314 3152
rect 6314 3120 6336 3152
rect 6365 3120 6386 3152
rect 6386 3120 6417 3152
rect 6446 3120 6458 3152
rect 6458 3120 6496 3152
rect 6496 3120 6498 3152
rect 6528 3120 6530 3152
rect 6530 3120 6568 3152
rect 6568 3120 6580 3152
rect 6609 3120 6640 3152
rect 6640 3120 6661 3152
rect 6690 3120 6712 3152
rect 6712 3120 6742 3152
rect 6771 3120 6784 3152
rect 6784 3120 6818 3152
rect 6818 3120 6823 3152
rect 6852 3152 6904 3172
rect 6933 3152 6985 3172
rect 7014 3152 7066 3172
rect 7096 3152 7148 3172
rect 7177 3152 7229 3172
rect 7258 3152 7310 3172
rect 7339 3152 7391 3172
rect 7420 3152 7472 3172
rect 6852 3120 6856 3152
rect 6856 3120 6890 3152
rect 6890 3120 6904 3152
rect 6933 3120 6962 3152
rect 6962 3120 6985 3152
rect 7014 3120 7034 3152
rect 7034 3120 7066 3152
rect 7096 3120 7106 3152
rect 7106 3120 7144 3152
rect 7144 3120 7148 3152
rect 7177 3120 7178 3152
rect 7178 3120 7216 3152
rect 7216 3120 7229 3152
rect 7258 3120 7288 3152
rect 7288 3120 7310 3152
rect 7339 3120 7360 3152
rect 7360 3120 7391 3152
rect 7420 3120 7432 3152
rect 7432 3120 7466 3152
rect 7466 3120 7472 3152
rect 7501 3152 7553 3172
rect 7582 3152 7634 3172
rect 7664 3152 7716 3172
rect 7745 3152 7797 3172
rect 7826 3152 7878 3172
rect 7907 3152 7959 3172
rect 7988 3152 8040 3172
rect 8069 3152 8121 3172
rect 7501 3120 7504 3152
rect 7504 3120 7538 3152
rect 7538 3120 7553 3152
rect 7582 3120 7610 3152
rect 7610 3120 7634 3152
rect 7664 3120 7682 3152
rect 7682 3120 7716 3152
rect 7745 3120 7754 3152
rect 7754 3120 7792 3152
rect 7792 3120 7797 3152
rect 7826 3120 7864 3152
rect 7864 3120 7878 3152
rect 7907 3120 7936 3152
rect 7936 3120 7959 3152
rect 7988 3120 8008 3152
rect 8008 3120 8040 3152
rect 8069 3120 8080 3152
rect 8080 3120 8114 3152
rect 8114 3120 8121 3152
rect 8150 3152 8202 3172
rect 8232 3152 8284 3172
rect 8313 3152 8365 3172
rect 8394 3152 8446 3172
rect 8475 3152 8527 3172
rect 8556 3152 8608 3172
rect 8637 3152 8689 3172
rect 8718 3152 8770 3172
rect 8150 3120 8152 3152
rect 8152 3120 8186 3152
rect 8186 3120 8202 3152
rect 8232 3120 8258 3152
rect 8258 3120 8284 3152
rect 8313 3120 8330 3152
rect 8330 3120 8365 3152
rect 8394 3120 8402 3152
rect 8402 3120 8440 3152
rect 8440 3120 8446 3152
rect 8475 3120 8512 3152
rect 8512 3120 8527 3152
rect 8556 3120 8584 3152
rect 8584 3120 8608 3152
rect 8637 3120 8656 3152
rect 8656 3120 8689 3152
rect 8718 3120 8728 3152
rect 8728 3120 8762 3152
rect 8762 3120 8770 3152
rect 8800 3152 8852 3172
rect 8881 3152 8933 3172
rect 8962 3152 9014 3172
rect 9043 3152 9095 3172
rect 9124 3152 9176 3172
rect 9205 3152 9257 3172
rect 9286 3152 9338 3172
rect 8800 3120 8834 3152
rect 8834 3120 8852 3152
rect 8881 3120 8906 3152
rect 8906 3120 8933 3152
rect 8962 3120 8978 3152
rect 8978 3120 9014 3152
rect 9043 3120 9050 3152
rect 9050 3120 9088 3152
rect 9088 3120 9095 3152
rect 9124 3120 9160 3152
rect 9160 3120 9176 3152
rect 9205 3120 9232 3152
rect 9232 3120 9257 3152
rect 9286 3120 9304 3152
rect 9304 3120 9338 3152
rect 9368 3152 9420 3172
rect 9449 3152 9501 3172
rect 9530 3152 9582 3172
rect 9611 3152 9663 3172
rect 9692 3152 9744 3172
rect 9773 3152 9825 3172
rect 9854 3152 9906 3172
rect 9936 3152 9988 3172
rect 9368 3120 9376 3152
rect 9376 3120 9410 3152
rect 9410 3120 9420 3152
rect 9449 3120 9482 3152
rect 9482 3120 9501 3152
rect 9530 3120 9554 3152
rect 9554 3120 9582 3152
rect 9611 3120 9626 3152
rect 9626 3120 9663 3152
rect 9692 3120 9698 3152
rect 9698 3120 9736 3152
rect 9736 3120 9744 3152
rect 9773 3120 9808 3152
rect 9808 3120 9825 3152
rect 9854 3120 9880 3152
rect 9880 3120 9906 3152
rect 9936 3120 9952 3152
rect 9952 3120 9986 3152
rect 9986 3120 9988 3152
rect 10017 3152 10069 3172
rect 10098 3152 10150 3172
rect 10179 3152 10231 3172
rect 10260 3152 10312 3172
rect 10341 3152 10393 3172
rect 10422 3152 10474 3172
rect 10504 3152 10556 3172
rect 10585 3152 10637 3172
rect 10017 3120 10024 3152
rect 10024 3120 10058 3152
rect 10058 3120 10069 3152
rect 10098 3120 10130 3152
rect 10130 3120 10150 3152
rect 10179 3120 10202 3152
rect 10202 3120 10231 3152
rect 10260 3120 10274 3152
rect 10274 3120 10312 3152
rect 10341 3120 10346 3152
rect 10346 3120 10384 3152
rect 10384 3120 10393 3152
rect 10422 3120 10456 3152
rect 10456 3120 10474 3152
rect 10504 3120 10528 3152
rect 10528 3120 10556 3152
rect 10585 3120 10600 3152
rect 10600 3120 10634 3152
rect 10634 3120 10637 3152
rect 10666 3152 10718 3172
rect 10747 3152 10799 3172
rect 10666 3120 10672 3152
rect 10672 3120 10706 3152
rect 10706 3120 10718 3152
rect 10747 3120 10778 3152
rect 10778 3120 10799 3152
rect 10828 3120 10880 3172
rect 10909 3120 10961 3172
rect 10990 3120 11042 3172
rect 11118 3120 11170 3172
rect 11199 3120 11251 3172
rect 11280 3120 11332 3172
rect 11361 3120 11413 3172
rect 11442 3120 11494 3172
rect 11523 3120 11575 3172
rect 11604 3120 11656 3172
rect 11686 3120 11738 3172
rect 11767 3120 11819 3172
rect 11848 3120 11900 3172
rect 11929 3120 11981 3172
rect 12010 3120 12062 3172
rect 12091 3120 12143 3172
rect 12172 3120 12224 3172
rect 12254 3120 12306 3172
rect 12335 3120 12387 3172
rect 12416 3151 12468 3172
rect 12497 3151 12549 3172
rect 12578 3151 12630 3172
rect 12659 3151 12711 3172
rect 12416 3120 12458 3151
rect 12458 3120 12468 3151
rect 12497 3120 12530 3151
rect 12530 3120 12549 3151
rect 12578 3120 12602 3151
rect 12602 3120 12630 3151
rect 12659 3120 12674 3151
rect 12674 3120 12708 3151
rect 12708 3120 12711 3151
rect 12740 3151 12792 3172
rect 12822 3151 12874 3172
rect 12903 3151 12955 3172
rect 12984 3151 13036 3172
rect 13065 3151 13117 3172
rect 13146 3151 13198 3172
rect 13227 3151 13279 3172
rect 13308 3151 13360 3172
rect 12740 3120 12746 3151
rect 12746 3120 12780 3151
rect 12780 3120 12792 3151
rect 12822 3120 12852 3151
rect 12852 3120 12874 3151
rect 12903 3120 12924 3151
rect 12924 3120 12955 3151
rect 12984 3120 12996 3151
rect 12996 3120 13034 3151
rect 13034 3120 13036 3151
rect 13065 3120 13068 3151
rect 13068 3120 13106 3151
rect 13106 3120 13117 3151
rect 13146 3120 13178 3151
rect 13178 3120 13198 3151
rect 13227 3120 13250 3151
rect 13250 3120 13279 3151
rect 13308 3120 13322 3151
rect 13322 3120 13356 3151
rect 13356 3120 13360 3151
rect 13390 3151 13442 3172
rect 13471 3151 13523 3172
rect 13552 3151 13604 3172
rect 13633 3151 13685 3172
rect 13714 3151 13766 3172
rect 13795 3151 13847 3172
rect 13876 3151 13928 3172
rect 13958 3151 14010 3172
rect 13390 3120 13394 3151
rect 13394 3120 13428 3151
rect 13428 3120 13442 3151
rect 13471 3120 13500 3151
rect 13500 3120 13523 3151
rect 13552 3120 13572 3151
rect 13572 3120 13604 3151
rect 13633 3120 13644 3151
rect 13644 3120 13682 3151
rect 13682 3120 13685 3151
rect 13714 3120 13716 3151
rect 13716 3120 13754 3151
rect 13754 3120 13766 3151
rect 13795 3120 13826 3151
rect 13826 3120 13847 3151
rect 13876 3120 13898 3151
rect 13898 3120 13928 3151
rect 13958 3120 13970 3151
rect 13970 3120 14004 3151
rect 14004 3120 14010 3151
rect 14039 3151 14091 3172
rect 14120 3151 14172 3172
rect 14201 3151 14253 3172
rect 14282 3151 14334 3172
rect 14363 3151 14415 3172
rect 14444 3151 14496 3172
rect 14526 3151 14578 3172
rect 14607 3151 14659 3172
rect 14039 3120 14042 3151
rect 14042 3120 14076 3151
rect 14076 3120 14091 3151
rect 14120 3120 14148 3151
rect 14148 3120 14172 3151
rect 14201 3120 14220 3151
rect 14220 3120 14253 3151
rect 14282 3120 14292 3151
rect 14292 3120 14330 3151
rect 14330 3120 14334 3151
rect 14363 3120 14364 3151
rect 14364 3120 14402 3151
rect 14402 3120 14415 3151
rect 14444 3120 14474 3151
rect 14474 3120 14496 3151
rect 14526 3120 14546 3151
rect 14546 3120 14578 3151
rect 14607 3120 14618 3151
rect 14618 3120 14652 3151
rect 14652 3120 14659 3151
rect 14688 3151 14740 3172
rect 14769 3151 14821 3172
rect 14850 3151 14902 3172
rect 14931 3151 14983 3172
rect 15012 3151 15064 3172
rect 15094 3151 15146 3172
rect 15175 3151 15227 3172
rect 15256 3151 15308 3172
rect 14688 3120 14690 3151
rect 14690 3120 14724 3151
rect 14724 3120 14740 3151
rect 14769 3120 14796 3151
rect 14796 3120 14821 3151
rect 14850 3120 14868 3151
rect 14868 3120 14902 3151
rect 14931 3120 14940 3151
rect 14940 3120 14978 3151
rect 14978 3120 14983 3151
rect 15012 3120 15050 3151
rect 15050 3120 15064 3151
rect 15094 3120 15122 3151
rect 15122 3120 15146 3151
rect 15175 3120 15194 3151
rect 15194 3120 15227 3151
rect 15256 3120 15266 3151
rect 15266 3120 15300 3151
rect 15300 3120 15308 3151
rect 15337 3151 15389 3172
rect 15418 3151 15470 3172
rect 15499 3151 15551 3172
rect 15580 3151 15632 3172
rect 15662 3151 15714 3172
rect 15743 3151 15795 3172
rect 15824 3151 15876 3172
rect 15337 3120 15338 3151
rect 15338 3120 15372 3151
rect 15372 3120 15389 3151
rect 15418 3120 15444 3151
rect 15444 3120 15470 3151
rect 15499 3120 15516 3151
rect 15516 3120 15551 3151
rect 15580 3120 15588 3151
rect 15588 3120 15626 3151
rect 15626 3120 15632 3151
rect 15662 3120 15698 3151
rect 15698 3120 15714 3151
rect 15743 3120 15770 3151
rect 15770 3120 15795 3151
rect 15824 3120 15842 3151
rect 15842 3120 15876 3151
rect 15905 3151 15957 3172
rect 15905 3120 15914 3151
rect 15914 3120 15948 3151
rect 15948 3120 15957 3151
rect 15986 3151 16038 3172
rect 16067 3151 16119 3172
rect 16148 3151 16200 3172
rect 16230 3151 16282 3172
rect 16311 3151 16363 3172
rect 16392 3151 16444 3172
rect 16473 3151 16525 3172
rect 15986 3120 16020 3151
rect 16020 3120 16038 3151
rect 16067 3120 16092 3151
rect 16092 3120 16119 3151
rect 16148 3120 16164 3151
rect 16164 3120 16200 3151
rect 16230 3120 16236 3151
rect 16236 3120 16274 3151
rect 16274 3120 16282 3151
rect 16311 3120 16346 3151
rect 16346 3120 16363 3151
rect 16392 3120 16418 3151
rect 16418 3120 16444 3151
rect 16473 3120 16490 3151
rect 16490 3120 16524 3151
rect 16524 3120 16525 3151
rect 16554 3151 16606 3172
rect 16635 3151 16687 3172
rect 16716 3151 16768 3172
rect 16798 3151 16850 3172
rect 16879 3151 16931 3172
rect 16960 3151 17012 3172
rect 17041 3151 17093 3172
rect 17122 3151 17174 3172
rect 16554 3120 16562 3151
rect 16562 3120 16596 3151
rect 16596 3120 16606 3151
rect 16635 3120 16668 3151
rect 16668 3120 16687 3151
rect 16716 3120 16740 3151
rect 16740 3120 16768 3151
rect 16798 3120 16812 3151
rect 16812 3120 16850 3151
rect 16879 3120 16884 3151
rect 16884 3120 16922 3151
rect 16922 3120 16931 3151
rect 16960 3120 16994 3151
rect 16994 3120 17012 3151
rect 17041 3120 17066 3151
rect 17066 3120 17093 3151
rect 17122 3120 17138 3151
rect 17138 3120 17172 3151
rect 17172 3120 17174 3151
rect 17203 3151 17255 3172
rect 17284 3151 17336 3172
rect 17366 3151 17418 3172
rect 17447 3151 17499 3172
rect 17528 3151 17580 3172
rect 17609 3151 17661 3172
rect 17690 3151 17742 3172
rect 17771 3151 17823 3172
rect 17203 3120 17210 3151
rect 17210 3120 17244 3151
rect 17244 3120 17255 3151
rect 17284 3120 17316 3151
rect 17316 3120 17336 3151
rect 17366 3120 17388 3151
rect 17388 3120 17418 3151
rect 17447 3120 17460 3151
rect 17460 3120 17498 3151
rect 17498 3120 17499 3151
rect 17528 3120 17532 3151
rect 17532 3120 17570 3151
rect 17570 3120 17580 3151
rect 17609 3120 17642 3151
rect 17642 3120 17661 3151
rect 17690 3120 17714 3151
rect 17714 3120 17742 3151
rect 17771 3120 17786 3151
rect 17786 3120 17820 3151
rect 17820 3120 17823 3151
rect 17852 3151 17904 3172
rect 17934 3151 17986 3172
rect 18015 3151 18067 3172
rect 18096 3151 18148 3172
rect 18177 3151 18229 3172
rect 18258 3151 18310 3172
rect 18339 3151 18391 3172
rect 18420 3151 18472 3172
rect 17852 3120 17858 3151
rect 17858 3120 17892 3151
rect 17892 3120 17904 3151
rect 17934 3120 17964 3151
rect 17964 3120 17986 3151
rect 18015 3120 18036 3151
rect 18036 3120 18067 3151
rect 18096 3120 18108 3151
rect 18108 3120 18146 3151
rect 18146 3120 18148 3151
rect 18177 3120 18180 3151
rect 18180 3120 18218 3151
rect 18218 3120 18229 3151
rect 18258 3120 18290 3151
rect 18290 3120 18310 3151
rect 18339 3120 18362 3151
rect 18362 3120 18391 3151
rect 18420 3120 18434 3151
rect 18434 3120 18468 3151
rect 18468 3120 18472 3151
rect 18502 3120 18554 3172
rect 18583 3151 18635 3172
rect 18583 3120 18597 3151
rect 18597 3120 18631 3151
rect 18631 3120 18635 3151
rect 18664 3151 18716 3172
rect 18745 3151 18797 3172
rect 18826 3151 18878 3172
rect 18907 3151 18959 3172
rect 18988 3151 19040 3172
rect 19070 3151 19122 3172
rect 19151 3151 19203 3172
rect 19232 3151 19284 3172
rect 18664 3120 18669 3151
rect 18669 3120 18703 3151
rect 18703 3120 18716 3151
rect 18745 3120 18775 3151
rect 18775 3120 18797 3151
rect 18826 3120 18847 3151
rect 18847 3120 18878 3151
rect 18907 3120 18919 3151
rect 18919 3120 18957 3151
rect 18957 3120 18959 3151
rect 18988 3120 18991 3151
rect 18991 3120 19029 3151
rect 19029 3120 19040 3151
rect 19070 3120 19101 3151
rect 19101 3120 19122 3151
rect 19151 3120 19173 3151
rect 19173 3120 19203 3151
rect 19232 3120 19245 3151
rect 19245 3120 19279 3151
rect 19279 3120 19284 3151
rect 19313 3151 19365 3172
rect 19394 3151 19446 3172
rect 19475 3151 19527 3172
rect 19556 3151 19608 3172
rect 19638 3151 19690 3172
rect 19719 3151 19771 3172
rect 19800 3151 19852 3172
rect 19881 3151 19933 3172
rect 19313 3120 19317 3151
rect 19317 3120 19351 3151
rect 19351 3120 19365 3151
rect 19394 3120 19423 3151
rect 19423 3120 19446 3151
rect 19475 3120 19495 3151
rect 19495 3120 19527 3151
rect 19556 3120 19567 3151
rect 19567 3120 19605 3151
rect 19605 3120 19608 3151
rect 19638 3120 19639 3151
rect 19639 3120 19677 3151
rect 19677 3120 19690 3151
rect 19719 3120 19749 3151
rect 19749 3120 19771 3151
rect 19800 3120 19821 3151
rect 19821 3120 19852 3151
rect 19881 3120 19893 3151
rect 19893 3120 19927 3151
rect 19927 3120 19933 3151
rect 19962 3151 20014 3172
rect 20043 3151 20095 3172
rect 20124 3151 20176 3172
rect 20206 3151 20258 3172
rect 20287 3151 20339 3172
rect 20368 3151 20420 3172
rect 20449 3151 20501 3172
rect 20530 3151 20582 3172
rect 19962 3120 19965 3151
rect 19965 3120 19999 3151
rect 19999 3120 20014 3151
rect 20043 3120 20071 3151
rect 20071 3120 20095 3151
rect 20124 3120 20143 3151
rect 20143 3120 20176 3151
rect 20206 3120 20215 3151
rect 20215 3120 20253 3151
rect 20253 3120 20258 3151
rect 20287 3120 20325 3151
rect 20325 3120 20339 3151
rect 20368 3120 20397 3151
rect 20397 3120 20420 3151
rect 20449 3120 20469 3151
rect 20469 3120 20501 3151
rect 20530 3120 20541 3151
rect 20541 3120 20575 3151
rect 20575 3120 20582 3151
rect 20611 3151 20663 3172
rect 20692 3151 20744 3172
rect 20774 3151 20826 3172
rect 20855 3151 20907 3172
rect 20936 3151 20988 3172
rect 21017 3151 21069 3172
rect 21098 3151 21150 3172
rect 21179 3151 21231 3172
rect 20611 3120 20613 3151
rect 20613 3120 20647 3151
rect 20647 3120 20663 3151
rect 20692 3120 20719 3151
rect 20719 3120 20744 3151
rect 20774 3120 20791 3151
rect 20791 3120 20826 3151
rect 20855 3120 20863 3151
rect 20863 3120 20901 3151
rect 20901 3120 20907 3151
rect 20936 3120 20973 3151
rect 20973 3120 20988 3151
rect 21017 3120 21045 3151
rect 21045 3120 21069 3151
rect 21098 3120 21117 3151
rect 21117 3120 21150 3151
rect 21179 3120 21189 3151
rect 21189 3120 21223 3151
rect 21223 3120 21231 3151
rect 21260 3151 21312 3172
rect 21342 3151 21394 3172
rect 21423 3151 21475 3172
rect 21504 3151 21556 3172
rect 21585 3151 21637 3172
rect 21666 3151 21718 3172
rect 21747 3151 21799 3172
rect 21260 3120 21261 3151
rect 21261 3120 21295 3151
rect 21295 3120 21312 3151
rect 21342 3120 21367 3151
rect 21367 3120 21394 3151
rect 21423 3120 21439 3151
rect 21439 3120 21475 3151
rect 21504 3120 21511 3151
rect 21511 3120 21549 3151
rect 21549 3120 21556 3151
rect 21585 3120 21621 3151
rect 21621 3120 21637 3151
rect 21666 3120 21693 3151
rect 21693 3120 21718 3151
rect 21747 3120 21765 3151
rect 21765 3120 21799 3151
rect 21828 3151 21880 3172
rect 21910 3151 21962 3172
rect 21991 3151 22043 3172
rect 22072 3151 22124 3172
rect 22153 3151 22205 3172
rect 22234 3151 22286 3172
rect 22315 3151 22367 3172
rect 22396 3151 22448 3172
rect 21828 3120 21837 3151
rect 21837 3120 21871 3151
rect 21871 3120 21880 3151
rect 21910 3120 21943 3151
rect 21943 3120 21962 3151
rect 21991 3120 22015 3151
rect 22015 3120 22043 3151
rect 22072 3120 22087 3151
rect 22087 3120 22124 3151
rect 22153 3120 22159 3151
rect 22159 3120 22197 3151
rect 22197 3120 22205 3151
rect 22234 3120 22269 3151
rect 22269 3120 22286 3151
rect 22315 3120 22341 3151
rect 22341 3120 22367 3151
rect 22396 3120 22413 3151
rect 22413 3120 22447 3151
rect 22447 3120 22448 3151
rect 22478 3151 22530 3172
rect 22559 3151 22611 3172
rect 22640 3151 22692 3172
rect 22721 3151 22773 3172
rect 22802 3151 22854 3172
rect 22883 3151 22935 3172
rect 22964 3151 23016 3172
rect 23046 3151 23098 3172
rect 22478 3120 22485 3151
rect 22485 3120 22519 3151
rect 22519 3120 22530 3151
rect 22559 3120 22591 3151
rect 22591 3120 22611 3151
rect 22640 3120 22663 3151
rect 22663 3120 22692 3151
rect 22721 3120 22735 3151
rect 22735 3120 22773 3151
rect 22802 3120 22807 3151
rect 22807 3120 22845 3151
rect 22845 3120 22854 3151
rect 22883 3120 22917 3151
rect 22917 3120 22935 3151
rect 22964 3120 22989 3151
rect 22989 3120 23016 3151
rect 23046 3120 23061 3151
rect 23061 3120 23095 3151
rect 23095 3120 23098 3151
rect 23127 3151 23179 3172
rect 23208 3151 23260 3172
rect 23289 3151 23341 3172
rect 23370 3151 23422 3172
rect 23451 3151 23503 3172
rect 23532 3151 23584 3172
rect 23614 3151 23666 3172
rect 23695 3151 23747 3172
rect 23127 3120 23133 3151
rect 23133 3120 23167 3151
rect 23167 3120 23179 3151
rect 23208 3120 23239 3151
rect 23239 3120 23260 3151
rect 23289 3120 23311 3151
rect 23311 3120 23341 3151
rect 23370 3120 23383 3151
rect 23383 3120 23421 3151
rect 23421 3120 23422 3151
rect 23451 3120 23455 3151
rect 23455 3120 23493 3151
rect 23493 3120 23503 3151
rect 23532 3120 23565 3151
rect 23565 3120 23584 3151
rect 23614 3120 23637 3151
rect 23637 3120 23666 3151
rect 23695 3120 23709 3151
rect 23709 3120 23743 3151
rect 23743 3120 23747 3151
rect 23776 3151 23828 3172
rect 23857 3151 23909 3172
rect 23938 3151 23990 3172
rect 24019 3151 24071 3172
rect 24100 3151 24152 3172
rect 24182 3151 24234 3172
rect 24263 3151 24315 3172
rect 24344 3151 24396 3172
rect 23776 3120 23781 3151
rect 23781 3120 23815 3151
rect 23815 3120 23828 3151
rect 23857 3120 23887 3151
rect 23887 3120 23909 3151
rect 23938 3120 23959 3151
rect 23959 3120 23990 3151
rect 24019 3120 24031 3151
rect 24031 3120 24069 3151
rect 24069 3120 24071 3151
rect 24100 3120 24103 3151
rect 24103 3120 24141 3151
rect 24141 3120 24152 3151
rect 24182 3120 24213 3151
rect 24213 3120 24234 3151
rect 24263 3120 24285 3151
rect 24285 3120 24315 3151
rect 24344 3120 24357 3151
rect 24357 3120 24391 3151
rect 24391 3120 24396 3151
rect 24425 3151 24477 3172
rect 24506 3151 24558 3172
rect 24587 3151 24639 3172
rect 24425 3120 24429 3151
rect 24429 3120 24463 3151
rect 24463 3120 24477 3151
rect 24506 3120 24535 3151
rect 24535 3120 24558 3151
rect 24587 3120 24607 3151
rect 24607 3120 24639 3151
rect 24668 3120 24720 3172
rect 3038 3016 3090 3068
rect 3120 3016 3172 3068
rect 3201 3016 3253 3068
rect 3282 3016 3334 3068
rect 3363 3016 3415 3068
rect 3444 3016 3496 3068
rect 3525 3016 3577 3068
rect 3606 3016 3658 3068
rect 3688 3016 3740 3068
rect 3769 3016 3821 3068
rect 3850 3016 3902 3068
rect 3931 3016 3983 3068
rect 4012 3016 4064 3068
rect 4093 3016 4145 3068
rect 4174 3016 4226 3068
rect 4256 3016 4308 3068
rect 4337 3016 4389 3068
rect 4418 3016 4470 3068
rect 4499 3016 4551 3068
rect 4580 3016 4632 3068
rect 4661 3016 4713 3068
rect 4742 3064 4794 3068
rect 4824 3064 4876 3068
rect 4742 3030 4768 3064
rect 4768 3030 4794 3064
rect 4824 3030 4840 3064
rect 4840 3030 4874 3064
rect 4874 3030 4876 3064
rect 4742 3016 4794 3030
rect 4824 3016 4876 3030
rect 4905 3064 4957 3068
rect 4986 3064 5038 3068
rect 5067 3064 5119 3068
rect 5148 3064 5200 3068
rect 5229 3064 5281 3068
rect 5310 3064 5362 3068
rect 5392 3064 5444 3068
rect 5473 3064 5525 3068
rect 4905 3030 4912 3064
rect 4912 3030 4946 3064
rect 4946 3030 4957 3064
rect 4986 3030 5018 3064
rect 5018 3030 5038 3064
rect 5067 3030 5090 3064
rect 5090 3030 5119 3064
rect 5148 3030 5162 3064
rect 5162 3030 5200 3064
rect 5229 3030 5234 3064
rect 5234 3030 5272 3064
rect 5272 3030 5281 3064
rect 5310 3030 5344 3064
rect 5344 3030 5362 3064
rect 5392 3030 5416 3064
rect 5416 3030 5444 3064
rect 5473 3030 5488 3064
rect 5488 3030 5522 3064
rect 5522 3030 5525 3064
rect 4905 3016 4957 3030
rect 4986 3016 5038 3030
rect 5067 3016 5119 3030
rect 5148 3016 5200 3030
rect 5229 3016 5281 3030
rect 5310 3016 5362 3030
rect 5392 3016 5444 3030
rect 5473 3016 5525 3030
rect 5554 3064 5606 3068
rect 5635 3064 5687 3068
rect 5716 3064 5768 3068
rect 5797 3064 5849 3068
rect 5878 3064 5930 3068
rect 5960 3064 6012 3068
rect 6041 3064 6093 3068
rect 6122 3064 6174 3068
rect 5554 3030 5560 3064
rect 5560 3030 5594 3064
rect 5594 3030 5606 3064
rect 5635 3030 5666 3064
rect 5666 3030 5687 3064
rect 5716 3030 5738 3064
rect 5738 3030 5768 3064
rect 5797 3030 5810 3064
rect 5810 3030 5848 3064
rect 5848 3030 5849 3064
rect 5878 3030 5882 3064
rect 5882 3030 5920 3064
rect 5920 3030 5930 3064
rect 5960 3030 5992 3064
rect 5992 3030 6012 3064
rect 6041 3030 6064 3064
rect 6064 3030 6093 3064
rect 6122 3030 6136 3064
rect 6136 3030 6170 3064
rect 6170 3030 6174 3064
rect 5554 3016 5606 3030
rect 5635 3016 5687 3030
rect 5716 3016 5768 3030
rect 5797 3016 5849 3030
rect 5878 3016 5930 3030
rect 5960 3016 6012 3030
rect 6041 3016 6093 3030
rect 6122 3016 6174 3030
rect 6203 3064 6255 3068
rect 6284 3064 6336 3068
rect 6365 3064 6417 3068
rect 6446 3064 6498 3068
rect 6528 3064 6580 3068
rect 6609 3064 6661 3068
rect 6690 3064 6742 3068
rect 6771 3064 6823 3068
rect 6203 3030 6208 3064
rect 6208 3030 6242 3064
rect 6242 3030 6255 3064
rect 6284 3030 6314 3064
rect 6314 3030 6336 3064
rect 6365 3030 6386 3064
rect 6386 3030 6417 3064
rect 6446 3030 6458 3064
rect 6458 3030 6496 3064
rect 6496 3030 6498 3064
rect 6528 3030 6530 3064
rect 6530 3030 6568 3064
rect 6568 3030 6580 3064
rect 6609 3030 6640 3064
rect 6640 3030 6661 3064
rect 6690 3030 6712 3064
rect 6712 3030 6742 3064
rect 6771 3030 6784 3064
rect 6784 3030 6818 3064
rect 6818 3030 6823 3064
rect 6203 3016 6255 3030
rect 6284 3016 6336 3030
rect 6365 3016 6417 3030
rect 6446 3016 6498 3030
rect 6528 3016 6580 3030
rect 6609 3016 6661 3030
rect 6690 3016 6742 3030
rect 6771 3016 6823 3030
rect 6852 3064 6904 3068
rect 6933 3064 6985 3068
rect 7014 3064 7066 3068
rect 7096 3064 7148 3068
rect 7177 3064 7229 3068
rect 7258 3064 7310 3068
rect 7339 3064 7391 3068
rect 7420 3064 7472 3068
rect 6852 3030 6856 3064
rect 6856 3030 6890 3064
rect 6890 3030 6904 3064
rect 6933 3030 6962 3064
rect 6962 3030 6985 3064
rect 7014 3030 7034 3064
rect 7034 3030 7066 3064
rect 7096 3030 7106 3064
rect 7106 3030 7144 3064
rect 7144 3030 7148 3064
rect 7177 3030 7178 3064
rect 7178 3030 7216 3064
rect 7216 3030 7229 3064
rect 7258 3030 7288 3064
rect 7288 3030 7310 3064
rect 7339 3030 7360 3064
rect 7360 3030 7391 3064
rect 7420 3030 7432 3064
rect 7432 3030 7466 3064
rect 7466 3030 7472 3064
rect 6852 3016 6904 3030
rect 6933 3016 6985 3030
rect 7014 3016 7066 3030
rect 7096 3016 7148 3030
rect 7177 3016 7229 3030
rect 7258 3016 7310 3030
rect 7339 3016 7391 3030
rect 7420 3016 7472 3030
rect 7501 3064 7553 3068
rect 7582 3064 7634 3068
rect 7664 3064 7716 3068
rect 7745 3064 7797 3068
rect 7826 3064 7878 3068
rect 7907 3064 7959 3068
rect 7988 3064 8040 3068
rect 8069 3064 8121 3068
rect 7501 3030 7504 3064
rect 7504 3030 7538 3064
rect 7538 3030 7553 3064
rect 7582 3030 7610 3064
rect 7610 3030 7634 3064
rect 7664 3030 7682 3064
rect 7682 3030 7716 3064
rect 7745 3030 7754 3064
rect 7754 3030 7792 3064
rect 7792 3030 7797 3064
rect 7826 3030 7864 3064
rect 7864 3030 7878 3064
rect 7907 3030 7936 3064
rect 7936 3030 7959 3064
rect 7988 3030 8008 3064
rect 8008 3030 8040 3064
rect 8069 3030 8080 3064
rect 8080 3030 8114 3064
rect 8114 3030 8121 3064
rect 7501 3016 7553 3030
rect 7582 3016 7634 3030
rect 7664 3016 7716 3030
rect 7745 3016 7797 3030
rect 7826 3016 7878 3030
rect 7907 3016 7959 3030
rect 7988 3016 8040 3030
rect 8069 3016 8121 3030
rect 8150 3064 8202 3068
rect 8232 3064 8284 3068
rect 8313 3064 8365 3068
rect 8394 3064 8446 3068
rect 8475 3064 8527 3068
rect 8556 3064 8608 3068
rect 8637 3064 8689 3068
rect 8718 3064 8770 3068
rect 8150 3030 8152 3064
rect 8152 3030 8186 3064
rect 8186 3030 8202 3064
rect 8232 3030 8258 3064
rect 8258 3030 8284 3064
rect 8313 3030 8330 3064
rect 8330 3030 8365 3064
rect 8394 3030 8402 3064
rect 8402 3030 8440 3064
rect 8440 3030 8446 3064
rect 8475 3030 8512 3064
rect 8512 3030 8527 3064
rect 8556 3030 8584 3064
rect 8584 3030 8608 3064
rect 8637 3030 8656 3064
rect 8656 3030 8689 3064
rect 8718 3030 8728 3064
rect 8728 3030 8762 3064
rect 8762 3030 8770 3064
rect 8150 3016 8202 3030
rect 8232 3016 8284 3030
rect 8313 3016 8365 3030
rect 8394 3016 8446 3030
rect 8475 3016 8527 3030
rect 8556 3016 8608 3030
rect 8637 3016 8689 3030
rect 8718 3016 8770 3030
rect 8800 3064 8852 3068
rect 8881 3064 8933 3068
rect 8962 3064 9014 3068
rect 9043 3064 9095 3068
rect 9124 3064 9176 3068
rect 9205 3064 9257 3068
rect 9286 3064 9338 3068
rect 8800 3030 8834 3064
rect 8834 3030 8852 3064
rect 8881 3030 8906 3064
rect 8906 3030 8933 3064
rect 8962 3030 8978 3064
rect 8978 3030 9014 3064
rect 9043 3030 9050 3064
rect 9050 3030 9088 3064
rect 9088 3030 9095 3064
rect 9124 3030 9160 3064
rect 9160 3030 9176 3064
rect 9205 3030 9232 3064
rect 9232 3030 9257 3064
rect 9286 3030 9304 3064
rect 9304 3030 9338 3064
rect 8800 3016 8852 3030
rect 8881 3016 8933 3030
rect 8962 3016 9014 3030
rect 9043 3016 9095 3030
rect 9124 3016 9176 3030
rect 9205 3016 9257 3030
rect 9286 3016 9338 3030
rect 9368 3064 9420 3068
rect 9449 3064 9501 3068
rect 9530 3064 9582 3068
rect 9611 3064 9663 3068
rect 9692 3064 9744 3068
rect 9773 3064 9825 3068
rect 9854 3064 9906 3068
rect 9936 3064 9988 3068
rect 9368 3030 9376 3064
rect 9376 3030 9410 3064
rect 9410 3030 9420 3064
rect 9449 3030 9482 3064
rect 9482 3030 9501 3064
rect 9530 3030 9554 3064
rect 9554 3030 9582 3064
rect 9611 3030 9626 3064
rect 9626 3030 9663 3064
rect 9692 3030 9698 3064
rect 9698 3030 9736 3064
rect 9736 3030 9744 3064
rect 9773 3030 9808 3064
rect 9808 3030 9825 3064
rect 9854 3030 9880 3064
rect 9880 3030 9906 3064
rect 9936 3030 9952 3064
rect 9952 3030 9986 3064
rect 9986 3030 9988 3064
rect 9368 3016 9420 3030
rect 9449 3016 9501 3030
rect 9530 3016 9582 3030
rect 9611 3016 9663 3030
rect 9692 3016 9744 3030
rect 9773 3016 9825 3030
rect 9854 3016 9906 3030
rect 9936 3016 9988 3030
rect 10017 3064 10069 3068
rect 10098 3064 10150 3068
rect 10179 3064 10231 3068
rect 10260 3064 10312 3068
rect 10341 3064 10393 3068
rect 10422 3064 10474 3068
rect 10504 3064 10556 3068
rect 10585 3064 10637 3068
rect 10017 3030 10024 3064
rect 10024 3030 10058 3064
rect 10058 3030 10069 3064
rect 10098 3030 10130 3064
rect 10130 3030 10150 3064
rect 10179 3030 10202 3064
rect 10202 3030 10231 3064
rect 10260 3030 10274 3064
rect 10274 3030 10312 3064
rect 10341 3030 10346 3064
rect 10346 3030 10384 3064
rect 10384 3030 10393 3064
rect 10422 3030 10456 3064
rect 10456 3030 10474 3064
rect 10504 3030 10528 3064
rect 10528 3030 10556 3064
rect 10585 3030 10600 3064
rect 10600 3030 10634 3064
rect 10634 3030 10637 3064
rect 10017 3016 10069 3030
rect 10098 3016 10150 3030
rect 10179 3016 10231 3030
rect 10260 3016 10312 3030
rect 10341 3016 10393 3030
rect 10422 3016 10474 3030
rect 10504 3016 10556 3030
rect 10585 3016 10637 3030
rect 10666 3064 10718 3068
rect 10747 3064 10799 3068
rect 10666 3030 10672 3064
rect 10672 3030 10706 3064
rect 10706 3030 10718 3064
rect 10747 3030 10778 3064
rect 10778 3030 10799 3064
rect 10666 3016 10718 3030
rect 10747 3016 10799 3030
rect 10828 3016 10880 3068
rect 10909 3016 10961 3068
rect 10990 3016 11042 3068
rect 11118 3016 11170 3068
rect 11199 3016 11251 3068
rect 11280 3016 11332 3068
rect 11361 3016 11413 3068
rect 11442 3016 11494 3068
rect 11523 3016 11575 3068
rect 11604 3016 11656 3068
rect 11686 3016 11738 3068
rect 11767 3016 11819 3068
rect 11848 3016 11900 3068
rect 11929 3016 11981 3068
rect 12010 3016 12062 3068
rect 12091 3016 12143 3068
rect 12172 3016 12224 3068
rect 12254 3016 12306 3068
rect 12335 3016 12387 3068
rect 12416 3063 12468 3068
rect 12497 3063 12549 3068
rect 12578 3063 12630 3068
rect 12659 3063 12711 3068
rect 12416 3029 12458 3063
rect 12458 3029 12468 3063
rect 12497 3029 12530 3063
rect 12530 3029 12549 3063
rect 12578 3029 12602 3063
rect 12602 3029 12630 3063
rect 12659 3029 12674 3063
rect 12674 3029 12708 3063
rect 12708 3029 12711 3063
rect 12416 3016 12468 3029
rect 12497 3016 12549 3029
rect 12578 3016 12630 3029
rect 12659 3016 12711 3029
rect 12740 3063 12792 3068
rect 12822 3063 12874 3068
rect 12903 3063 12955 3068
rect 12984 3063 13036 3068
rect 13065 3063 13117 3068
rect 13146 3063 13198 3068
rect 13227 3063 13279 3068
rect 13308 3063 13360 3068
rect 12740 3029 12746 3063
rect 12746 3029 12780 3063
rect 12780 3029 12792 3063
rect 12822 3029 12852 3063
rect 12852 3029 12874 3063
rect 12903 3029 12924 3063
rect 12924 3029 12955 3063
rect 12984 3029 12996 3063
rect 12996 3029 13034 3063
rect 13034 3029 13036 3063
rect 13065 3029 13068 3063
rect 13068 3029 13106 3063
rect 13106 3029 13117 3063
rect 13146 3029 13178 3063
rect 13178 3029 13198 3063
rect 13227 3029 13250 3063
rect 13250 3029 13279 3063
rect 13308 3029 13322 3063
rect 13322 3029 13356 3063
rect 13356 3029 13360 3063
rect 12740 3016 12792 3029
rect 12822 3016 12874 3029
rect 12903 3016 12955 3029
rect 12984 3016 13036 3029
rect 13065 3016 13117 3029
rect 13146 3016 13198 3029
rect 13227 3016 13279 3029
rect 13308 3016 13360 3029
rect 13390 3063 13442 3068
rect 13471 3063 13523 3068
rect 13552 3063 13604 3068
rect 13633 3063 13685 3068
rect 13714 3063 13766 3068
rect 13795 3063 13847 3068
rect 13876 3063 13928 3068
rect 13958 3063 14010 3068
rect 13390 3029 13394 3063
rect 13394 3029 13428 3063
rect 13428 3029 13442 3063
rect 13471 3029 13500 3063
rect 13500 3029 13523 3063
rect 13552 3029 13572 3063
rect 13572 3029 13604 3063
rect 13633 3029 13644 3063
rect 13644 3029 13682 3063
rect 13682 3029 13685 3063
rect 13714 3029 13716 3063
rect 13716 3029 13754 3063
rect 13754 3029 13766 3063
rect 13795 3029 13826 3063
rect 13826 3029 13847 3063
rect 13876 3029 13898 3063
rect 13898 3029 13928 3063
rect 13958 3029 13970 3063
rect 13970 3029 14004 3063
rect 14004 3029 14010 3063
rect 13390 3016 13442 3029
rect 13471 3016 13523 3029
rect 13552 3016 13604 3029
rect 13633 3016 13685 3029
rect 13714 3016 13766 3029
rect 13795 3016 13847 3029
rect 13876 3016 13928 3029
rect 13958 3016 14010 3029
rect 14039 3063 14091 3068
rect 14120 3063 14172 3068
rect 14201 3063 14253 3068
rect 14282 3063 14334 3068
rect 14363 3063 14415 3068
rect 14444 3063 14496 3068
rect 14526 3063 14578 3068
rect 14607 3063 14659 3068
rect 14039 3029 14042 3063
rect 14042 3029 14076 3063
rect 14076 3029 14091 3063
rect 14120 3029 14148 3063
rect 14148 3029 14172 3063
rect 14201 3029 14220 3063
rect 14220 3029 14253 3063
rect 14282 3029 14292 3063
rect 14292 3029 14330 3063
rect 14330 3029 14334 3063
rect 14363 3029 14364 3063
rect 14364 3029 14402 3063
rect 14402 3029 14415 3063
rect 14444 3029 14474 3063
rect 14474 3029 14496 3063
rect 14526 3029 14546 3063
rect 14546 3029 14578 3063
rect 14607 3029 14618 3063
rect 14618 3029 14652 3063
rect 14652 3029 14659 3063
rect 14039 3016 14091 3029
rect 14120 3016 14172 3029
rect 14201 3016 14253 3029
rect 14282 3016 14334 3029
rect 14363 3016 14415 3029
rect 14444 3016 14496 3029
rect 14526 3016 14578 3029
rect 14607 3016 14659 3029
rect 14688 3063 14740 3068
rect 14769 3063 14821 3068
rect 14850 3063 14902 3068
rect 14931 3063 14983 3068
rect 15012 3063 15064 3068
rect 15094 3063 15146 3068
rect 15175 3063 15227 3068
rect 15256 3063 15308 3068
rect 14688 3029 14690 3063
rect 14690 3029 14724 3063
rect 14724 3029 14740 3063
rect 14769 3029 14796 3063
rect 14796 3029 14821 3063
rect 14850 3029 14868 3063
rect 14868 3029 14902 3063
rect 14931 3029 14940 3063
rect 14940 3029 14978 3063
rect 14978 3029 14983 3063
rect 15012 3029 15050 3063
rect 15050 3029 15064 3063
rect 15094 3029 15122 3063
rect 15122 3029 15146 3063
rect 15175 3029 15194 3063
rect 15194 3029 15227 3063
rect 15256 3029 15266 3063
rect 15266 3029 15300 3063
rect 15300 3029 15308 3063
rect 14688 3016 14740 3029
rect 14769 3016 14821 3029
rect 14850 3016 14902 3029
rect 14931 3016 14983 3029
rect 15012 3016 15064 3029
rect 15094 3016 15146 3029
rect 15175 3016 15227 3029
rect 15256 3016 15308 3029
rect 15337 3063 15389 3068
rect 15418 3063 15470 3068
rect 15499 3063 15551 3068
rect 15580 3063 15632 3068
rect 15662 3063 15714 3068
rect 15743 3063 15795 3068
rect 15824 3063 15876 3068
rect 15337 3029 15338 3063
rect 15338 3029 15372 3063
rect 15372 3029 15389 3063
rect 15418 3029 15444 3063
rect 15444 3029 15470 3063
rect 15499 3029 15516 3063
rect 15516 3029 15551 3063
rect 15580 3029 15588 3063
rect 15588 3029 15626 3063
rect 15626 3029 15632 3063
rect 15662 3029 15698 3063
rect 15698 3029 15714 3063
rect 15743 3029 15770 3063
rect 15770 3029 15795 3063
rect 15824 3029 15842 3063
rect 15842 3029 15876 3063
rect 15337 3016 15389 3029
rect 15418 3016 15470 3029
rect 15499 3016 15551 3029
rect 15580 3016 15632 3029
rect 15662 3016 15714 3029
rect 15743 3016 15795 3029
rect 15824 3016 15876 3029
rect 15905 3063 15957 3068
rect 15905 3029 15914 3063
rect 15914 3029 15948 3063
rect 15948 3029 15957 3063
rect 15905 3016 15957 3029
rect 15986 3063 16038 3068
rect 16067 3063 16119 3068
rect 16148 3063 16200 3068
rect 16230 3063 16282 3068
rect 16311 3063 16363 3068
rect 16392 3063 16444 3068
rect 16473 3063 16525 3068
rect 15986 3029 16020 3063
rect 16020 3029 16038 3063
rect 16067 3029 16092 3063
rect 16092 3029 16119 3063
rect 16148 3029 16164 3063
rect 16164 3029 16200 3063
rect 16230 3029 16236 3063
rect 16236 3029 16274 3063
rect 16274 3029 16282 3063
rect 16311 3029 16346 3063
rect 16346 3029 16363 3063
rect 16392 3029 16418 3063
rect 16418 3029 16444 3063
rect 16473 3029 16490 3063
rect 16490 3029 16524 3063
rect 16524 3029 16525 3063
rect 15986 3016 16038 3029
rect 16067 3016 16119 3029
rect 16148 3016 16200 3029
rect 16230 3016 16282 3029
rect 16311 3016 16363 3029
rect 16392 3016 16444 3029
rect 16473 3016 16525 3029
rect 16554 3063 16606 3068
rect 16635 3063 16687 3068
rect 16716 3063 16768 3068
rect 16798 3063 16850 3068
rect 16879 3063 16931 3068
rect 16960 3063 17012 3068
rect 17041 3063 17093 3068
rect 17122 3063 17174 3068
rect 16554 3029 16562 3063
rect 16562 3029 16596 3063
rect 16596 3029 16606 3063
rect 16635 3029 16668 3063
rect 16668 3029 16687 3063
rect 16716 3029 16740 3063
rect 16740 3029 16768 3063
rect 16798 3029 16812 3063
rect 16812 3029 16850 3063
rect 16879 3029 16884 3063
rect 16884 3029 16922 3063
rect 16922 3029 16931 3063
rect 16960 3029 16994 3063
rect 16994 3029 17012 3063
rect 17041 3029 17066 3063
rect 17066 3029 17093 3063
rect 17122 3029 17138 3063
rect 17138 3029 17172 3063
rect 17172 3029 17174 3063
rect 16554 3016 16606 3029
rect 16635 3016 16687 3029
rect 16716 3016 16768 3029
rect 16798 3016 16850 3029
rect 16879 3016 16931 3029
rect 16960 3016 17012 3029
rect 17041 3016 17093 3029
rect 17122 3016 17174 3029
rect 17203 3063 17255 3068
rect 17284 3063 17336 3068
rect 17366 3063 17418 3068
rect 17447 3063 17499 3068
rect 17528 3063 17580 3068
rect 17609 3063 17661 3068
rect 17690 3063 17742 3068
rect 17771 3063 17823 3068
rect 17203 3029 17210 3063
rect 17210 3029 17244 3063
rect 17244 3029 17255 3063
rect 17284 3029 17316 3063
rect 17316 3029 17336 3063
rect 17366 3029 17388 3063
rect 17388 3029 17418 3063
rect 17447 3029 17460 3063
rect 17460 3029 17498 3063
rect 17498 3029 17499 3063
rect 17528 3029 17532 3063
rect 17532 3029 17570 3063
rect 17570 3029 17580 3063
rect 17609 3029 17642 3063
rect 17642 3029 17661 3063
rect 17690 3029 17714 3063
rect 17714 3029 17742 3063
rect 17771 3029 17786 3063
rect 17786 3029 17820 3063
rect 17820 3029 17823 3063
rect 17203 3016 17255 3029
rect 17284 3016 17336 3029
rect 17366 3016 17418 3029
rect 17447 3016 17499 3029
rect 17528 3016 17580 3029
rect 17609 3016 17661 3029
rect 17690 3016 17742 3029
rect 17771 3016 17823 3029
rect 17852 3063 17904 3068
rect 17934 3063 17986 3068
rect 18015 3063 18067 3068
rect 18096 3063 18148 3068
rect 18177 3063 18229 3068
rect 18258 3063 18310 3068
rect 18339 3063 18391 3068
rect 18420 3063 18472 3068
rect 17852 3029 17858 3063
rect 17858 3029 17892 3063
rect 17892 3029 17904 3063
rect 17934 3029 17964 3063
rect 17964 3029 17986 3063
rect 18015 3029 18036 3063
rect 18036 3029 18067 3063
rect 18096 3029 18108 3063
rect 18108 3029 18146 3063
rect 18146 3029 18148 3063
rect 18177 3029 18180 3063
rect 18180 3029 18218 3063
rect 18218 3029 18229 3063
rect 18258 3029 18290 3063
rect 18290 3029 18310 3063
rect 18339 3029 18362 3063
rect 18362 3029 18391 3063
rect 18420 3029 18434 3063
rect 18434 3029 18468 3063
rect 18468 3029 18472 3063
rect 17852 3016 17904 3029
rect 17934 3016 17986 3029
rect 18015 3016 18067 3029
rect 18096 3016 18148 3029
rect 18177 3016 18229 3029
rect 18258 3016 18310 3029
rect 18339 3016 18391 3029
rect 18420 3016 18472 3029
rect 18502 3016 18554 3068
rect 18583 3063 18635 3068
rect 18583 3029 18597 3063
rect 18597 3029 18631 3063
rect 18631 3029 18635 3063
rect 18583 3016 18635 3029
rect 18664 3063 18716 3068
rect 18745 3063 18797 3068
rect 18826 3063 18878 3068
rect 18907 3063 18959 3068
rect 18988 3063 19040 3068
rect 19070 3063 19122 3068
rect 19151 3063 19203 3068
rect 19232 3063 19284 3068
rect 18664 3029 18669 3063
rect 18669 3029 18703 3063
rect 18703 3029 18716 3063
rect 18745 3029 18775 3063
rect 18775 3029 18797 3063
rect 18826 3029 18847 3063
rect 18847 3029 18878 3063
rect 18907 3029 18919 3063
rect 18919 3029 18957 3063
rect 18957 3029 18959 3063
rect 18988 3029 18991 3063
rect 18991 3029 19029 3063
rect 19029 3029 19040 3063
rect 19070 3029 19101 3063
rect 19101 3029 19122 3063
rect 19151 3029 19173 3063
rect 19173 3029 19203 3063
rect 19232 3029 19245 3063
rect 19245 3029 19279 3063
rect 19279 3029 19284 3063
rect 18664 3016 18716 3029
rect 18745 3016 18797 3029
rect 18826 3016 18878 3029
rect 18907 3016 18959 3029
rect 18988 3016 19040 3029
rect 19070 3016 19122 3029
rect 19151 3016 19203 3029
rect 19232 3016 19284 3029
rect 19313 3063 19365 3068
rect 19394 3063 19446 3068
rect 19475 3063 19527 3068
rect 19556 3063 19608 3068
rect 19638 3063 19690 3068
rect 19719 3063 19771 3068
rect 19800 3063 19852 3068
rect 19881 3063 19933 3068
rect 19313 3029 19317 3063
rect 19317 3029 19351 3063
rect 19351 3029 19365 3063
rect 19394 3029 19423 3063
rect 19423 3029 19446 3063
rect 19475 3029 19495 3063
rect 19495 3029 19527 3063
rect 19556 3029 19567 3063
rect 19567 3029 19605 3063
rect 19605 3029 19608 3063
rect 19638 3029 19639 3063
rect 19639 3029 19677 3063
rect 19677 3029 19690 3063
rect 19719 3029 19749 3063
rect 19749 3029 19771 3063
rect 19800 3029 19821 3063
rect 19821 3029 19852 3063
rect 19881 3029 19893 3063
rect 19893 3029 19927 3063
rect 19927 3029 19933 3063
rect 19313 3016 19365 3029
rect 19394 3016 19446 3029
rect 19475 3016 19527 3029
rect 19556 3016 19608 3029
rect 19638 3016 19690 3029
rect 19719 3016 19771 3029
rect 19800 3016 19852 3029
rect 19881 3016 19933 3029
rect 19962 3063 20014 3068
rect 20043 3063 20095 3068
rect 20124 3063 20176 3068
rect 20206 3063 20258 3068
rect 20287 3063 20339 3068
rect 20368 3063 20420 3068
rect 20449 3063 20501 3068
rect 20530 3063 20582 3068
rect 19962 3029 19965 3063
rect 19965 3029 19999 3063
rect 19999 3029 20014 3063
rect 20043 3029 20071 3063
rect 20071 3029 20095 3063
rect 20124 3029 20143 3063
rect 20143 3029 20176 3063
rect 20206 3029 20215 3063
rect 20215 3029 20253 3063
rect 20253 3029 20258 3063
rect 20287 3029 20325 3063
rect 20325 3029 20339 3063
rect 20368 3029 20397 3063
rect 20397 3029 20420 3063
rect 20449 3029 20469 3063
rect 20469 3029 20501 3063
rect 20530 3029 20541 3063
rect 20541 3029 20575 3063
rect 20575 3029 20582 3063
rect 19962 3016 20014 3029
rect 20043 3016 20095 3029
rect 20124 3016 20176 3029
rect 20206 3016 20258 3029
rect 20287 3016 20339 3029
rect 20368 3016 20420 3029
rect 20449 3016 20501 3029
rect 20530 3016 20582 3029
rect 20611 3063 20663 3068
rect 20692 3063 20744 3068
rect 20774 3063 20826 3068
rect 20855 3063 20907 3068
rect 20936 3063 20988 3068
rect 21017 3063 21069 3068
rect 21098 3063 21150 3068
rect 21179 3063 21231 3068
rect 20611 3029 20613 3063
rect 20613 3029 20647 3063
rect 20647 3029 20663 3063
rect 20692 3029 20719 3063
rect 20719 3029 20744 3063
rect 20774 3029 20791 3063
rect 20791 3029 20826 3063
rect 20855 3029 20863 3063
rect 20863 3029 20901 3063
rect 20901 3029 20907 3063
rect 20936 3029 20973 3063
rect 20973 3029 20988 3063
rect 21017 3029 21045 3063
rect 21045 3029 21069 3063
rect 21098 3029 21117 3063
rect 21117 3029 21150 3063
rect 21179 3029 21189 3063
rect 21189 3029 21223 3063
rect 21223 3029 21231 3063
rect 20611 3016 20663 3029
rect 20692 3016 20744 3029
rect 20774 3016 20826 3029
rect 20855 3016 20907 3029
rect 20936 3016 20988 3029
rect 21017 3016 21069 3029
rect 21098 3016 21150 3029
rect 21179 3016 21231 3029
rect 21260 3063 21312 3068
rect 21342 3063 21394 3068
rect 21423 3063 21475 3068
rect 21504 3063 21556 3068
rect 21585 3063 21637 3068
rect 21666 3063 21718 3068
rect 21747 3063 21799 3068
rect 21260 3029 21261 3063
rect 21261 3029 21295 3063
rect 21295 3029 21312 3063
rect 21342 3029 21367 3063
rect 21367 3029 21394 3063
rect 21423 3029 21439 3063
rect 21439 3029 21475 3063
rect 21504 3029 21511 3063
rect 21511 3029 21549 3063
rect 21549 3029 21556 3063
rect 21585 3029 21621 3063
rect 21621 3029 21637 3063
rect 21666 3029 21693 3063
rect 21693 3029 21718 3063
rect 21747 3029 21765 3063
rect 21765 3029 21799 3063
rect 21260 3016 21312 3029
rect 21342 3016 21394 3029
rect 21423 3016 21475 3029
rect 21504 3016 21556 3029
rect 21585 3016 21637 3029
rect 21666 3016 21718 3029
rect 21747 3016 21799 3029
rect 21828 3063 21880 3068
rect 21910 3063 21962 3068
rect 21991 3063 22043 3068
rect 22072 3063 22124 3068
rect 22153 3063 22205 3068
rect 22234 3063 22286 3068
rect 22315 3063 22367 3068
rect 22396 3063 22448 3068
rect 21828 3029 21837 3063
rect 21837 3029 21871 3063
rect 21871 3029 21880 3063
rect 21910 3029 21943 3063
rect 21943 3029 21962 3063
rect 21991 3029 22015 3063
rect 22015 3029 22043 3063
rect 22072 3029 22087 3063
rect 22087 3029 22124 3063
rect 22153 3029 22159 3063
rect 22159 3029 22197 3063
rect 22197 3029 22205 3063
rect 22234 3029 22269 3063
rect 22269 3029 22286 3063
rect 22315 3029 22341 3063
rect 22341 3029 22367 3063
rect 22396 3029 22413 3063
rect 22413 3029 22447 3063
rect 22447 3029 22448 3063
rect 21828 3016 21880 3029
rect 21910 3016 21962 3029
rect 21991 3016 22043 3029
rect 22072 3016 22124 3029
rect 22153 3016 22205 3029
rect 22234 3016 22286 3029
rect 22315 3016 22367 3029
rect 22396 3016 22448 3029
rect 22478 3063 22530 3068
rect 22559 3063 22611 3068
rect 22640 3063 22692 3068
rect 22721 3063 22773 3068
rect 22802 3063 22854 3068
rect 22883 3063 22935 3068
rect 22964 3063 23016 3068
rect 23046 3063 23098 3068
rect 22478 3029 22485 3063
rect 22485 3029 22519 3063
rect 22519 3029 22530 3063
rect 22559 3029 22591 3063
rect 22591 3029 22611 3063
rect 22640 3029 22663 3063
rect 22663 3029 22692 3063
rect 22721 3029 22735 3063
rect 22735 3029 22773 3063
rect 22802 3029 22807 3063
rect 22807 3029 22845 3063
rect 22845 3029 22854 3063
rect 22883 3029 22917 3063
rect 22917 3029 22935 3063
rect 22964 3029 22989 3063
rect 22989 3029 23016 3063
rect 23046 3029 23061 3063
rect 23061 3029 23095 3063
rect 23095 3029 23098 3063
rect 22478 3016 22530 3029
rect 22559 3016 22611 3029
rect 22640 3016 22692 3029
rect 22721 3016 22773 3029
rect 22802 3016 22854 3029
rect 22883 3016 22935 3029
rect 22964 3016 23016 3029
rect 23046 3016 23098 3029
rect 23127 3063 23179 3068
rect 23208 3063 23260 3068
rect 23289 3063 23341 3068
rect 23370 3063 23422 3068
rect 23451 3063 23503 3068
rect 23532 3063 23584 3068
rect 23614 3063 23666 3068
rect 23695 3063 23747 3068
rect 23127 3029 23133 3063
rect 23133 3029 23167 3063
rect 23167 3029 23179 3063
rect 23208 3029 23239 3063
rect 23239 3029 23260 3063
rect 23289 3029 23311 3063
rect 23311 3029 23341 3063
rect 23370 3029 23383 3063
rect 23383 3029 23421 3063
rect 23421 3029 23422 3063
rect 23451 3029 23455 3063
rect 23455 3029 23493 3063
rect 23493 3029 23503 3063
rect 23532 3029 23565 3063
rect 23565 3029 23584 3063
rect 23614 3029 23637 3063
rect 23637 3029 23666 3063
rect 23695 3029 23709 3063
rect 23709 3029 23743 3063
rect 23743 3029 23747 3063
rect 23127 3016 23179 3029
rect 23208 3016 23260 3029
rect 23289 3016 23341 3029
rect 23370 3016 23422 3029
rect 23451 3016 23503 3029
rect 23532 3016 23584 3029
rect 23614 3016 23666 3029
rect 23695 3016 23747 3029
rect 23776 3063 23828 3068
rect 23857 3063 23909 3068
rect 23938 3063 23990 3068
rect 24019 3063 24071 3068
rect 24100 3063 24152 3068
rect 24182 3063 24234 3068
rect 24263 3063 24315 3068
rect 24344 3063 24396 3068
rect 23776 3029 23781 3063
rect 23781 3029 23815 3063
rect 23815 3029 23828 3063
rect 23857 3029 23887 3063
rect 23887 3029 23909 3063
rect 23938 3029 23959 3063
rect 23959 3029 23990 3063
rect 24019 3029 24031 3063
rect 24031 3029 24069 3063
rect 24069 3029 24071 3063
rect 24100 3029 24103 3063
rect 24103 3029 24141 3063
rect 24141 3029 24152 3063
rect 24182 3029 24213 3063
rect 24213 3029 24234 3063
rect 24263 3029 24285 3063
rect 24285 3029 24315 3063
rect 24344 3029 24357 3063
rect 24357 3029 24391 3063
rect 24391 3029 24396 3063
rect 23776 3016 23828 3029
rect 23857 3016 23909 3029
rect 23938 3016 23990 3029
rect 24019 3016 24071 3029
rect 24100 3016 24152 3029
rect 24182 3016 24234 3029
rect 24263 3016 24315 3029
rect 24344 3016 24396 3029
rect 24425 3063 24477 3068
rect 24506 3063 24558 3068
rect 24587 3063 24639 3068
rect 24425 3029 24429 3063
rect 24429 3029 24463 3063
rect 24463 3029 24477 3063
rect 24506 3029 24535 3063
rect 24535 3029 24558 3063
rect 24587 3029 24607 3063
rect 24607 3029 24639 3063
rect 24425 3016 24477 3029
rect 24506 3016 24558 3029
rect 24587 3016 24639 3029
rect 24668 3016 24720 3068
rect 3038 2912 3090 2964
rect 3120 2912 3172 2964
rect 3201 2912 3253 2964
rect 3282 2912 3334 2964
rect 3363 2912 3415 2964
rect 3444 2912 3496 2964
rect 3525 2912 3577 2964
rect 3606 2912 3658 2964
rect 3688 2912 3740 2964
rect 3769 2912 3821 2964
rect 3850 2912 3902 2964
rect 3931 2912 3983 2964
rect 4012 2912 4064 2964
rect 4093 2912 4145 2964
rect 4174 2912 4226 2964
rect 4256 2912 4308 2964
rect 4337 2912 4389 2964
rect 4418 2912 4470 2964
rect 4499 2912 4551 2964
rect 4580 2912 4632 2964
rect 4661 2912 4713 2964
rect 4742 2942 4768 2964
rect 4768 2942 4794 2964
rect 4824 2942 4840 2964
rect 4840 2942 4874 2964
rect 4874 2942 4876 2964
rect 4742 2912 4794 2942
rect 4824 2912 4876 2942
rect 4905 2942 4912 2964
rect 4912 2942 4946 2964
rect 4946 2942 4957 2964
rect 4986 2942 5018 2964
rect 5018 2942 5038 2964
rect 5067 2942 5090 2964
rect 5090 2942 5119 2964
rect 5148 2942 5162 2964
rect 5162 2942 5200 2964
rect 5229 2942 5234 2964
rect 5234 2942 5272 2964
rect 5272 2942 5281 2964
rect 5310 2942 5344 2964
rect 5344 2942 5362 2964
rect 5392 2942 5416 2964
rect 5416 2942 5444 2964
rect 5473 2942 5488 2964
rect 5488 2942 5522 2964
rect 5522 2942 5525 2964
rect 4905 2912 4957 2942
rect 4986 2912 5038 2942
rect 5067 2912 5119 2942
rect 5148 2912 5200 2942
rect 5229 2912 5281 2942
rect 5310 2912 5362 2942
rect 5392 2912 5444 2942
rect 5473 2912 5525 2942
rect 5554 2942 5560 2964
rect 5560 2942 5594 2964
rect 5594 2942 5606 2964
rect 5635 2942 5666 2964
rect 5666 2942 5687 2964
rect 5716 2942 5738 2964
rect 5738 2942 5768 2964
rect 5797 2942 5810 2964
rect 5810 2942 5848 2964
rect 5848 2942 5849 2964
rect 5878 2942 5882 2964
rect 5882 2942 5920 2964
rect 5920 2942 5930 2964
rect 5960 2942 5992 2964
rect 5992 2942 6012 2964
rect 6041 2942 6064 2964
rect 6064 2942 6093 2964
rect 6122 2942 6136 2964
rect 6136 2942 6170 2964
rect 6170 2942 6174 2964
rect 5554 2912 5606 2942
rect 5635 2912 5687 2942
rect 5716 2912 5768 2942
rect 5797 2912 5849 2942
rect 5878 2912 5930 2942
rect 5960 2912 6012 2942
rect 6041 2912 6093 2942
rect 6122 2912 6174 2942
rect 6203 2942 6208 2964
rect 6208 2942 6242 2964
rect 6242 2942 6255 2964
rect 6284 2942 6314 2964
rect 6314 2942 6336 2964
rect 6365 2942 6386 2964
rect 6386 2942 6417 2964
rect 6446 2942 6458 2964
rect 6458 2942 6496 2964
rect 6496 2942 6498 2964
rect 6528 2942 6530 2964
rect 6530 2942 6568 2964
rect 6568 2942 6580 2964
rect 6609 2942 6640 2964
rect 6640 2942 6661 2964
rect 6690 2942 6712 2964
rect 6712 2942 6742 2964
rect 6771 2942 6784 2964
rect 6784 2942 6818 2964
rect 6818 2942 6823 2964
rect 6203 2912 6255 2942
rect 6284 2912 6336 2942
rect 6365 2912 6417 2942
rect 6446 2912 6498 2942
rect 6528 2912 6580 2942
rect 6609 2912 6661 2942
rect 6690 2912 6742 2942
rect 6771 2912 6823 2942
rect 6852 2942 6856 2964
rect 6856 2942 6890 2964
rect 6890 2942 6904 2964
rect 6933 2942 6962 2964
rect 6962 2942 6985 2964
rect 7014 2942 7034 2964
rect 7034 2942 7066 2964
rect 7096 2942 7106 2964
rect 7106 2942 7144 2964
rect 7144 2942 7148 2964
rect 7177 2942 7178 2964
rect 7178 2942 7216 2964
rect 7216 2942 7229 2964
rect 7258 2942 7288 2964
rect 7288 2942 7310 2964
rect 7339 2942 7360 2964
rect 7360 2942 7391 2964
rect 7420 2942 7432 2964
rect 7432 2942 7466 2964
rect 7466 2942 7472 2964
rect 6852 2912 6904 2942
rect 6933 2912 6985 2942
rect 7014 2912 7066 2942
rect 7096 2912 7148 2942
rect 7177 2912 7229 2942
rect 7258 2912 7310 2942
rect 7339 2912 7391 2942
rect 7420 2912 7472 2942
rect 7501 2942 7504 2964
rect 7504 2942 7538 2964
rect 7538 2942 7553 2964
rect 7582 2942 7610 2964
rect 7610 2942 7634 2964
rect 7664 2942 7682 2964
rect 7682 2942 7716 2964
rect 7745 2942 7754 2964
rect 7754 2942 7792 2964
rect 7792 2942 7797 2964
rect 7826 2942 7864 2964
rect 7864 2942 7878 2964
rect 7907 2942 7936 2964
rect 7936 2942 7959 2964
rect 7988 2942 8008 2964
rect 8008 2942 8040 2964
rect 8069 2942 8080 2964
rect 8080 2942 8114 2964
rect 8114 2942 8121 2964
rect 7501 2912 7553 2942
rect 7582 2912 7634 2942
rect 7664 2912 7716 2942
rect 7745 2912 7797 2942
rect 7826 2912 7878 2942
rect 7907 2912 7959 2942
rect 7988 2912 8040 2942
rect 8069 2912 8121 2942
rect 8150 2942 8152 2964
rect 8152 2942 8186 2964
rect 8186 2942 8202 2964
rect 8232 2942 8258 2964
rect 8258 2942 8284 2964
rect 8313 2942 8330 2964
rect 8330 2942 8365 2964
rect 8394 2942 8402 2964
rect 8402 2942 8440 2964
rect 8440 2942 8446 2964
rect 8475 2942 8512 2964
rect 8512 2942 8527 2964
rect 8556 2942 8584 2964
rect 8584 2942 8608 2964
rect 8637 2942 8656 2964
rect 8656 2942 8689 2964
rect 8718 2942 8728 2964
rect 8728 2942 8762 2964
rect 8762 2942 8770 2964
rect 8150 2912 8202 2942
rect 8232 2912 8284 2942
rect 8313 2912 8365 2942
rect 8394 2912 8446 2942
rect 8475 2912 8527 2942
rect 8556 2912 8608 2942
rect 8637 2912 8689 2942
rect 8718 2912 8770 2942
rect 8800 2942 8834 2964
rect 8834 2942 8852 2964
rect 8881 2942 8906 2964
rect 8906 2942 8933 2964
rect 8962 2942 8978 2964
rect 8978 2942 9014 2964
rect 9043 2942 9050 2964
rect 9050 2942 9088 2964
rect 9088 2942 9095 2964
rect 9124 2942 9160 2964
rect 9160 2942 9176 2964
rect 9205 2942 9232 2964
rect 9232 2942 9257 2964
rect 9286 2942 9304 2964
rect 9304 2942 9338 2964
rect 8800 2912 8852 2942
rect 8881 2912 8933 2942
rect 8962 2912 9014 2942
rect 9043 2912 9095 2942
rect 9124 2912 9176 2942
rect 9205 2912 9257 2942
rect 9286 2912 9338 2942
rect 9368 2942 9376 2964
rect 9376 2942 9410 2964
rect 9410 2942 9420 2964
rect 9449 2942 9482 2964
rect 9482 2942 9501 2964
rect 9530 2942 9554 2964
rect 9554 2942 9582 2964
rect 9611 2942 9626 2964
rect 9626 2942 9663 2964
rect 9692 2942 9698 2964
rect 9698 2942 9736 2964
rect 9736 2942 9744 2964
rect 9773 2942 9808 2964
rect 9808 2942 9825 2964
rect 9854 2942 9880 2964
rect 9880 2942 9906 2964
rect 9936 2942 9952 2964
rect 9952 2942 9986 2964
rect 9986 2942 9988 2964
rect 9368 2912 9420 2942
rect 9449 2912 9501 2942
rect 9530 2912 9582 2942
rect 9611 2912 9663 2942
rect 9692 2912 9744 2942
rect 9773 2912 9825 2942
rect 9854 2912 9906 2942
rect 9936 2912 9988 2942
rect 10017 2942 10024 2964
rect 10024 2942 10058 2964
rect 10058 2942 10069 2964
rect 10098 2942 10130 2964
rect 10130 2942 10150 2964
rect 10179 2942 10202 2964
rect 10202 2942 10231 2964
rect 10260 2942 10274 2964
rect 10274 2942 10312 2964
rect 10341 2942 10346 2964
rect 10346 2942 10384 2964
rect 10384 2942 10393 2964
rect 10422 2942 10456 2964
rect 10456 2942 10474 2964
rect 10504 2942 10528 2964
rect 10528 2942 10556 2964
rect 10585 2942 10600 2964
rect 10600 2942 10634 2964
rect 10634 2942 10637 2964
rect 10017 2912 10069 2942
rect 10098 2912 10150 2942
rect 10179 2912 10231 2942
rect 10260 2912 10312 2942
rect 10341 2912 10393 2942
rect 10422 2912 10474 2942
rect 10504 2912 10556 2942
rect 10585 2912 10637 2942
rect 10666 2942 10672 2964
rect 10672 2942 10706 2964
rect 10706 2942 10718 2964
rect 10747 2942 10778 2964
rect 10778 2942 10799 2964
rect 10666 2912 10718 2942
rect 10747 2912 10799 2942
rect 10828 2912 10880 2964
rect 10909 2912 10961 2964
rect 10990 2912 11042 2964
rect 11118 2912 11170 2964
rect 11199 2912 11251 2964
rect 11280 2912 11332 2964
rect 11361 2912 11413 2964
rect 11442 2912 11494 2964
rect 11523 2912 11575 2964
rect 11604 2912 11656 2964
rect 11686 2912 11738 2964
rect 11767 2912 11819 2964
rect 11848 2912 11900 2964
rect 11929 2912 11981 2964
rect 12010 2912 12062 2964
rect 12091 2912 12143 2964
rect 12172 2912 12224 2964
rect 12254 2912 12306 2964
rect 12335 2912 12387 2964
rect 12416 2941 12458 2964
rect 12458 2941 12468 2964
rect 12497 2941 12530 2964
rect 12530 2941 12549 2964
rect 12578 2941 12602 2964
rect 12602 2941 12630 2964
rect 12659 2941 12674 2964
rect 12674 2941 12708 2964
rect 12708 2941 12711 2964
rect 12416 2912 12468 2941
rect 12497 2912 12549 2941
rect 12578 2912 12630 2941
rect 12659 2912 12711 2941
rect 12740 2941 12746 2964
rect 12746 2941 12780 2964
rect 12780 2941 12792 2964
rect 12822 2941 12852 2964
rect 12852 2941 12874 2964
rect 12903 2941 12924 2964
rect 12924 2941 12955 2964
rect 12984 2941 12996 2964
rect 12996 2941 13034 2964
rect 13034 2941 13036 2964
rect 13065 2941 13068 2964
rect 13068 2941 13106 2964
rect 13106 2941 13117 2964
rect 13146 2941 13178 2964
rect 13178 2941 13198 2964
rect 13227 2941 13250 2964
rect 13250 2941 13279 2964
rect 13308 2941 13322 2964
rect 13322 2941 13356 2964
rect 13356 2941 13360 2964
rect 12740 2912 12792 2941
rect 12822 2912 12874 2941
rect 12903 2912 12955 2941
rect 12984 2912 13036 2941
rect 13065 2912 13117 2941
rect 13146 2912 13198 2941
rect 13227 2912 13279 2941
rect 13308 2912 13360 2941
rect 13390 2941 13394 2964
rect 13394 2941 13428 2964
rect 13428 2941 13442 2964
rect 13471 2941 13500 2964
rect 13500 2941 13523 2964
rect 13552 2941 13572 2964
rect 13572 2941 13604 2964
rect 13633 2941 13644 2964
rect 13644 2941 13682 2964
rect 13682 2941 13685 2964
rect 13714 2941 13716 2964
rect 13716 2941 13754 2964
rect 13754 2941 13766 2964
rect 13795 2941 13826 2964
rect 13826 2941 13847 2964
rect 13876 2941 13898 2964
rect 13898 2941 13928 2964
rect 13958 2941 13970 2964
rect 13970 2941 14004 2964
rect 14004 2941 14010 2964
rect 13390 2912 13442 2941
rect 13471 2912 13523 2941
rect 13552 2912 13604 2941
rect 13633 2912 13685 2941
rect 13714 2912 13766 2941
rect 13795 2912 13847 2941
rect 13876 2912 13928 2941
rect 13958 2912 14010 2941
rect 14039 2941 14042 2964
rect 14042 2941 14076 2964
rect 14076 2941 14091 2964
rect 14120 2941 14148 2964
rect 14148 2941 14172 2964
rect 14201 2941 14220 2964
rect 14220 2941 14253 2964
rect 14282 2941 14292 2964
rect 14292 2941 14330 2964
rect 14330 2941 14334 2964
rect 14363 2941 14364 2964
rect 14364 2941 14402 2964
rect 14402 2941 14415 2964
rect 14444 2941 14474 2964
rect 14474 2941 14496 2964
rect 14526 2941 14546 2964
rect 14546 2941 14578 2964
rect 14607 2941 14618 2964
rect 14618 2941 14652 2964
rect 14652 2941 14659 2964
rect 14039 2912 14091 2941
rect 14120 2912 14172 2941
rect 14201 2912 14253 2941
rect 14282 2912 14334 2941
rect 14363 2912 14415 2941
rect 14444 2912 14496 2941
rect 14526 2912 14578 2941
rect 14607 2912 14659 2941
rect 14688 2941 14690 2964
rect 14690 2941 14724 2964
rect 14724 2941 14740 2964
rect 14769 2941 14796 2964
rect 14796 2941 14821 2964
rect 14850 2941 14868 2964
rect 14868 2941 14902 2964
rect 14931 2941 14940 2964
rect 14940 2941 14978 2964
rect 14978 2941 14983 2964
rect 15012 2941 15050 2964
rect 15050 2941 15064 2964
rect 15094 2941 15122 2964
rect 15122 2941 15146 2964
rect 15175 2941 15194 2964
rect 15194 2941 15227 2964
rect 15256 2941 15266 2964
rect 15266 2941 15300 2964
rect 15300 2941 15308 2964
rect 14688 2912 14740 2941
rect 14769 2912 14821 2941
rect 14850 2912 14902 2941
rect 14931 2912 14983 2941
rect 15012 2912 15064 2941
rect 15094 2912 15146 2941
rect 15175 2912 15227 2941
rect 15256 2912 15308 2941
rect 15337 2941 15338 2964
rect 15338 2941 15372 2964
rect 15372 2941 15389 2964
rect 15418 2941 15444 2964
rect 15444 2941 15470 2964
rect 15499 2941 15516 2964
rect 15516 2941 15551 2964
rect 15580 2941 15588 2964
rect 15588 2941 15626 2964
rect 15626 2941 15632 2964
rect 15662 2941 15698 2964
rect 15698 2941 15714 2964
rect 15743 2941 15770 2964
rect 15770 2941 15795 2964
rect 15824 2941 15842 2964
rect 15842 2941 15876 2964
rect 15337 2912 15389 2941
rect 15418 2912 15470 2941
rect 15499 2912 15551 2941
rect 15580 2912 15632 2941
rect 15662 2912 15714 2941
rect 15743 2912 15795 2941
rect 15824 2912 15876 2941
rect 15905 2941 15914 2964
rect 15914 2941 15948 2964
rect 15948 2941 15957 2964
rect 15905 2912 15957 2941
rect 15986 2941 16020 2964
rect 16020 2941 16038 2964
rect 16067 2941 16092 2964
rect 16092 2941 16119 2964
rect 16148 2941 16164 2964
rect 16164 2941 16200 2964
rect 16230 2941 16236 2964
rect 16236 2941 16274 2964
rect 16274 2941 16282 2964
rect 16311 2941 16346 2964
rect 16346 2941 16363 2964
rect 16392 2941 16418 2964
rect 16418 2941 16444 2964
rect 16473 2941 16490 2964
rect 16490 2941 16524 2964
rect 16524 2941 16525 2964
rect 15986 2912 16038 2941
rect 16067 2912 16119 2941
rect 16148 2912 16200 2941
rect 16230 2912 16282 2941
rect 16311 2912 16363 2941
rect 16392 2912 16444 2941
rect 16473 2912 16525 2941
rect 16554 2941 16562 2964
rect 16562 2941 16596 2964
rect 16596 2941 16606 2964
rect 16635 2941 16668 2964
rect 16668 2941 16687 2964
rect 16716 2941 16740 2964
rect 16740 2941 16768 2964
rect 16798 2941 16812 2964
rect 16812 2941 16850 2964
rect 16879 2941 16884 2964
rect 16884 2941 16922 2964
rect 16922 2941 16931 2964
rect 16960 2941 16994 2964
rect 16994 2941 17012 2964
rect 17041 2941 17066 2964
rect 17066 2941 17093 2964
rect 17122 2941 17138 2964
rect 17138 2941 17172 2964
rect 17172 2941 17174 2964
rect 16554 2912 16606 2941
rect 16635 2912 16687 2941
rect 16716 2912 16768 2941
rect 16798 2912 16850 2941
rect 16879 2912 16931 2941
rect 16960 2912 17012 2941
rect 17041 2912 17093 2941
rect 17122 2912 17174 2941
rect 17203 2941 17210 2964
rect 17210 2941 17244 2964
rect 17244 2941 17255 2964
rect 17284 2941 17316 2964
rect 17316 2941 17336 2964
rect 17366 2941 17388 2964
rect 17388 2941 17418 2964
rect 17447 2941 17460 2964
rect 17460 2941 17498 2964
rect 17498 2941 17499 2964
rect 17528 2941 17532 2964
rect 17532 2941 17570 2964
rect 17570 2941 17580 2964
rect 17609 2941 17642 2964
rect 17642 2941 17661 2964
rect 17690 2941 17714 2964
rect 17714 2941 17742 2964
rect 17771 2941 17786 2964
rect 17786 2941 17820 2964
rect 17820 2941 17823 2964
rect 17203 2912 17255 2941
rect 17284 2912 17336 2941
rect 17366 2912 17418 2941
rect 17447 2912 17499 2941
rect 17528 2912 17580 2941
rect 17609 2912 17661 2941
rect 17690 2912 17742 2941
rect 17771 2912 17823 2941
rect 17852 2941 17858 2964
rect 17858 2941 17892 2964
rect 17892 2941 17904 2964
rect 17934 2941 17964 2964
rect 17964 2941 17986 2964
rect 18015 2941 18036 2964
rect 18036 2941 18067 2964
rect 18096 2941 18108 2964
rect 18108 2941 18146 2964
rect 18146 2941 18148 2964
rect 18177 2941 18180 2964
rect 18180 2941 18218 2964
rect 18218 2941 18229 2964
rect 18258 2941 18290 2964
rect 18290 2941 18310 2964
rect 18339 2941 18362 2964
rect 18362 2941 18391 2964
rect 18420 2941 18434 2964
rect 18434 2941 18468 2964
rect 18468 2941 18472 2964
rect 17852 2912 17904 2941
rect 17934 2912 17986 2941
rect 18015 2912 18067 2941
rect 18096 2912 18148 2941
rect 18177 2912 18229 2941
rect 18258 2912 18310 2941
rect 18339 2912 18391 2941
rect 18420 2912 18472 2941
rect 18502 2912 18554 2964
rect 18583 2941 18597 2964
rect 18597 2941 18631 2964
rect 18631 2941 18635 2964
rect 18583 2912 18635 2941
rect 18664 2941 18669 2964
rect 18669 2941 18703 2964
rect 18703 2941 18716 2964
rect 18745 2941 18775 2964
rect 18775 2941 18797 2964
rect 18826 2941 18847 2964
rect 18847 2941 18878 2964
rect 18907 2941 18919 2964
rect 18919 2941 18957 2964
rect 18957 2941 18959 2964
rect 18988 2941 18991 2964
rect 18991 2941 19029 2964
rect 19029 2941 19040 2964
rect 19070 2941 19101 2964
rect 19101 2941 19122 2964
rect 19151 2941 19173 2964
rect 19173 2941 19203 2964
rect 19232 2941 19245 2964
rect 19245 2941 19279 2964
rect 19279 2941 19284 2964
rect 18664 2912 18716 2941
rect 18745 2912 18797 2941
rect 18826 2912 18878 2941
rect 18907 2912 18959 2941
rect 18988 2912 19040 2941
rect 19070 2912 19122 2941
rect 19151 2912 19203 2941
rect 19232 2912 19284 2941
rect 19313 2941 19317 2964
rect 19317 2941 19351 2964
rect 19351 2941 19365 2964
rect 19394 2941 19423 2964
rect 19423 2941 19446 2964
rect 19475 2941 19495 2964
rect 19495 2941 19527 2964
rect 19556 2941 19567 2964
rect 19567 2941 19605 2964
rect 19605 2941 19608 2964
rect 19638 2941 19639 2964
rect 19639 2941 19677 2964
rect 19677 2941 19690 2964
rect 19719 2941 19749 2964
rect 19749 2941 19771 2964
rect 19800 2941 19821 2964
rect 19821 2941 19852 2964
rect 19881 2941 19893 2964
rect 19893 2941 19927 2964
rect 19927 2941 19933 2964
rect 19313 2912 19365 2941
rect 19394 2912 19446 2941
rect 19475 2912 19527 2941
rect 19556 2912 19608 2941
rect 19638 2912 19690 2941
rect 19719 2912 19771 2941
rect 19800 2912 19852 2941
rect 19881 2912 19933 2941
rect 19962 2941 19965 2964
rect 19965 2941 19999 2964
rect 19999 2941 20014 2964
rect 20043 2941 20071 2964
rect 20071 2941 20095 2964
rect 20124 2941 20143 2964
rect 20143 2941 20176 2964
rect 20206 2941 20215 2964
rect 20215 2941 20253 2964
rect 20253 2941 20258 2964
rect 20287 2941 20325 2964
rect 20325 2941 20339 2964
rect 20368 2941 20397 2964
rect 20397 2941 20420 2964
rect 20449 2941 20469 2964
rect 20469 2941 20501 2964
rect 20530 2941 20541 2964
rect 20541 2941 20575 2964
rect 20575 2941 20582 2964
rect 19962 2912 20014 2941
rect 20043 2912 20095 2941
rect 20124 2912 20176 2941
rect 20206 2912 20258 2941
rect 20287 2912 20339 2941
rect 20368 2912 20420 2941
rect 20449 2912 20501 2941
rect 20530 2912 20582 2941
rect 20611 2941 20613 2964
rect 20613 2941 20647 2964
rect 20647 2941 20663 2964
rect 20692 2941 20719 2964
rect 20719 2941 20744 2964
rect 20774 2941 20791 2964
rect 20791 2941 20826 2964
rect 20855 2941 20863 2964
rect 20863 2941 20901 2964
rect 20901 2941 20907 2964
rect 20936 2941 20973 2964
rect 20973 2941 20988 2964
rect 21017 2941 21045 2964
rect 21045 2941 21069 2964
rect 21098 2941 21117 2964
rect 21117 2941 21150 2964
rect 21179 2941 21189 2964
rect 21189 2941 21223 2964
rect 21223 2941 21231 2964
rect 20611 2912 20663 2941
rect 20692 2912 20744 2941
rect 20774 2912 20826 2941
rect 20855 2912 20907 2941
rect 20936 2912 20988 2941
rect 21017 2912 21069 2941
rect 21098 2912 21150 2941
rect 21179 2912 21231 2941
rect 21260 2941 21261 2964
rect 21261 2941 21295 2964
rect 21295 2941 21312 2964
rect 21342 2941 21367 2964
rect 21367 2941 21394 2964
rect 21423 2941 21439 2964
rect 21439 2941 21475 2964
rect 21504 2941 21511 2964
rect 21511 2941 21549 2964
rect 21549 2941 21556 2964
rect 21585 2941 21621 2964
rect 21621 2941 21637 2964
rect 21666 2941 21693 2964
rect 21693 2941 21718 2964
rect 21747 2941 21765 2964
rect 21765 2941 21799 2964
rect 21260 2912 21312 2941
rect 21342 2912 21394 2941
rect 21423 2912 21475 2941
rect 21504 2912 21556 2941
rect 21585 2912 21637 2941
rect 21666 2912 21718 2941
rect 21747 2912 21799 2941
rect 21828 2941 21837 2964
rect 21837 2941 21871 2964
rect 21871 2941 21880 2964
rect 21910 2941 21943 2964
rect 21943 2941 21962 2964
rect 21991 2941 22015 2964
rect 22015 2941 22043 2964
rect 22072 2941 22087 2964
rect 22087 2941 22124 2964
rect 22153 2941 22159 2964
rect 22159 2941 22197 2964
rect 22197 2941 22205 2964
rect 22234 2941 22269 2964
rect 22269 2941 22286 2964
rect 22315 2941 22341 2964
rect 22341 2941 22367 2964
rect 22396 2941 22413 2964
rect 22413 2941 22447 2964
rect 22447 2941 22448 2964
rect 21828 2912 21880 2941
rect 21910 2912 21962 2941
rect 21991 2912 22043 2941
rect 22072 2912 22124 2941
rect 22153 2912 22205 2941
rect 22234 2912 22286 2941
rect 22315 2912 22367 2941
rect 22396 2912 22448 2941
rect 22478 2941 22485 2964
rect 22485 2941 22519 2964
rect 22519 2941 22530 2964
rect 22559 2941 22591 2964
rect 22591 2941 22611 2964
rect 22640 2941 22663 2964
rect 22663 2941 22692 2964
rect 22721 2941 22735 2964
rect 22735 2941 22773 2964
rect 22802 2941 22807 2964
rect 22807 2941 22845 2964
rect 22845 2941 22854 2964
rect 22883 2941 22917 2964
rect 22917 2941 22935 2964
rect 22964 2941 22989 2964
rect 22989 2941 23016 2964
rect 23046 2941 23061 2964
rect 23061 2941 23095 2964
rect 23095 2941 23098 2964
rect 22478 2912 22530 2941
rect 22559 2912 22611 2941
rect 22640 2912 22692 2941
rect 22721 2912 22773 2941
rect 22802 2912 22854 2941
rect 22883 2912 22935 2941
rect 22964 2912 23016 2941
rect 23046 2912 23098 2941
rect 23127 2941 23133 2964
rect 23133 2941 23167 2964
rect 23167 2941 23179 2964
rect 23208 2941 23239 2964
rect 23239 2941 23260 2964
rect 23289 2941 23311 2964
rect 23311 2941 23341 2964
rect 23370 2941 23383 2964
rect 23383 2941 23421 2964
rect 23421 2941 23422 2964
rect 23451 2941 23455 2964
rect 23455 2941 23493 2964
rect 23493 2941 23503 2964
rect 23532 2941 23565 2964
rect 23565 2941 23584 2964
rect 23614 2941 23637 2964
rect 23637 2941 23666 2964
rect 23695 2941 23709 2964
rect 23709 2941 23743 2964
rect 23743 2941 23747 2964
rect 23127 2912 23179 2941
rect 23208 2912 23260 2941
rect 23289 2912 23341 2941
rect 23370 2912 23422 2941
rect 23451 2912 23503 2941
rect 23532 2912 23584 2941
rect 23614 2912 23666 2941
rect 23695 2912 23747 2941
rect 23776 2941 23781 2964
rect 23781 2941 23815 2964
rect 23815 2941 23828 2964
rect 23857 2941 23887 2964
rect 23887 2941 23909 2964
rect 23938 2941 23959 2964
rect 23959 2941 23990 2964
rect 24019 2941 24031 2964
rect 24031 2941 24069 2964
rect 24069 2941 24071 2964
rect 24100 2941 24103 2964
rect 24103 2941 24141 2964
rect 24141 2941 24152 2964
rect 24182 2941 24213 2964
rect 24213 2941 24234 2964
rect 24263 2941 24285 2964
rect 24285 2941 24315 2964
rect 24344 2941 24357 2964
rect 24357 2941 24391 2964
rect 24391 2941 24396 2964
rect 23776 2912 23828 2941
rect 23857 2912 23909 2941
rect 23938 2912 23990 2941
rect 24019 2912 24071 2941
rect 24100 2912 24152 2941
rect 24182 2912 24234 2941
rect 24263 2912 24315 2941
rect 24344 2912 24396 2941
rect 24425 2941 24429 2964
rect 24429 2941 24463 2964
rect 24463 2941 24477 2964
rect 24506 2941 24535 2964
rect 24535 2941 24558 2964
rect 24587 2941 24607 2964
rect 24607 2941 24639 2964
rect 24425 2912 24477 2941
rect 24506 2912 24558 2941
rect 24587 2912 24639 2941
rect 24668 2912 24720 2964
rect 4919 2107 4971 2667
rect 5155 2107 5207 2667
rect 5391 2107 5443 2667
rect 5627 2107 5679 2667
rect 5863 2107 5915 2667
rect 6099 2107 6151 2667
rect 6335 2107 6387 2667
rect 6571 2107 6623 2667
rect 6917 2107 6969 2667
rect 7153 2107 7205 2667
rect 7389 2107 7398 2667
rect 7398 2107 7432 2667
rect 7432 2107 7441 2667
rect 7625 2107 7677 2667
rect 7861 2107 7913 2667
rect 8097 2107 8149 2667
rect 8333 2107 8385 2667
rect 8569 2107 8621 2667
rect 8915 2107 8967 2667
rect 9151 2107 9203 2667
rect 9387 2107 9439 2667
rect 9623 2107 9675 2667
rect 9859 2107 9911 2667
rect 10095 2107 10147 2667
rect 10331 2107 10383 2667
rect 10567 2107 10619 2667
rect 12491 2106 12543 2666
rect 12609 2106 12661 2666
rect 12727 2106 12736 2666
rect 12736 2106 12770 2666
rect 12770 2106 12779 2666
rect 12845 2106 12854 2666
rect 12854 2106 12888 2666
rect 12888 2106 12897 2666
rect 12963 2106 12972 2666
rect 12972 2106 13006 2666
rect 13006 2106 13015 2666
rect 13081 2106 13090 2666
rect 13090 2106 13124 2666
rect 13124 2106 13133 2666
rect 13199 2106 13208 2666
rect 13208 2106 13242 2666
rect 13242 2106 13251 2666
rect 13317 2106 13326 2666
rect 13326 2106 13360 2666
rect 13360 2106 13369 2666
rect 13435 2106 13444 2666
rect 13444 2106 13478 2666
rect 13478 2106 13487 2666
rect 13553 2106 13562 2666
rect 13562 2106 13596 2666
rect 13596 2106 13605 2666
rect 13671 2106 13680 2666
rect 13680 2106 13714 2666
rect 13714 2106 13723 2666
rect 13789 2106 13798 2666
rect 13798 2106 13832 2666
rect 13832 2106 13841 2666
rect 13907 2106 13916 2666
rect 13916 2106 13950 2666
rect 13950 2106 13959 2666
rect 14025 2106 14034 2666
rect 14034 2106 14068 2666
rect 14068 2106 14077 2666
rect 14143 2106 14152 2666
rect 14152 2106 14186 2666
rect 14186 2106 14195 2666
rect 14261 2106 14270 2666
rect 14270 2106 14304 2666
rect 14304 2106 14313 2666
rect 14379 2106 14388 2666
rect 14388 2106 14422 2666
rect 14422 2106 14431 2666
rect 14497 2106 14506 2666
rect 14506 2106 14540 2666
rect 14540 2106 14549 2666
rect 14615 2106 14624 2666
rect 14624 2106 14658 2666
rect 14658 2106 14667 2666
rect 14733 2106 14742 2666
rect 14742 2106 14776 2666
rect 14776 2106 14785 2666
rect 14851 2106 14860 2666
rect 14860 2106 14894 2666
rect 14894 2106 14903 2666
rect 14969 2106 14978 2666
rect 14978 2106 15012 2666
rect 15012 2106 15021 2666
rect 15087 2106 15096 2666
rect 15096 2106 15130 2666
rect 15130 2106 15139 2666
rect 15205 2106 15214 2666
rect 15214 2106 15248 2666
rect 15248 2106 15257 2666
rect 15323 2106 15332 2666
rect 15332 2106 15366 2666
rect 15366 2106 15375 2666
rect 15441 2106 15450 2666
rect 15450 2106 15484 2666
rect 15484 2106 15493 2666
rect 16614 2106 16666 2666
rect 16732 2106 16784 2666
rect 16850 2106 16859 2666
rect 16859 2106 16893 2666
rect 16893 2106 16902 2666
rect 16968 2106 16977 2666
rect 16977 2106 17011 2666
rect 17011 2106 17020 2666
rect 17086 2106 17095 2666
rect 17095 2106 17129 2666
rect 17129 2106 17138 2666
rect 17204 2106 17213 2666
rect 17213 2106 17247 2666
rect 17247 2106 17256 2666
rect 17322 2106 17331 2666
rect 17331 2106 17365 2666
rect 17365 2106 17374 2666
rect 17440 2106 17449 2666
rect 17449 2106 17483 2666
rect 17483 2106 17492 2666
rect 17558 2106 17567 2666
rect 17567 2106 17601 2666
rect 17601 2106 17610 2666
rect 17676 2106 17685 2666
rect 17685 2106 17719 2666
rect 17719 2106 17728 2666
rect 17794 2106 17803 2666
rect 17803 2106 17837 2666
rect 17837 2106 17846 2666
rect 17912 2106 17921 2666
rect 17921 2106 17955 2666
rect 17955 2106 17964 2666
rect 18030 2106 18039 2666
rect 18039 2106 18073 2666
rect 18073 2106 18082 2666
rect 18148 2106 18157 2666
rect 18157 2106 18191 2666
rect 18191 2106 18200 2666
rect 18266 2106 18275 2666
rect 18275 2106 18309 2666
rect 18309 2106 18318 2666
rect 18384 2106 18393 2666
rect 18393 2106 18427 2666
rect 18427 2106 18436 2666
rect 18502 2106 18511 2666
rect 18511 2106 18545 2666
rect 18545 2106 18554 2666
rect 18620 2106 18629 2666
rect 18629 2106 18663 2666
rect 18663 2106 18672 2666
rect 18738 2106 18747 2666
rect 18747 2106 18781 2666
rect 18781 2106 18790 2666
rect 18856 2106 18865 2666
rect 18865 2106 18899 2666
rect 18899 2106 18908 2666
rect 18974 2106 18983 2666
rect 18983 2106 19017 2666
rect 19017 2106 19026 2666
rect 19092 2106 19101 2666
rect 19101 2106 19135 2666
rect 19135 2106 19144 2666
rect 19210 2106 19219 2666
rect 19219 2106 19253 2666
rect 19253 2106 19262 2666
rect 19328 2106 19337 2666
rect 19337 2106 19371 2666
rect 19371 2106 19380 2666
rect 19446 2106 19455 2666
rect 19455 2106 19489 2666
rect 19489 2106 19498 2666
rect 19564 2106 19573 2666
rect 19573 2106 19607 2666
rect 19607 2106 19616 2666
rect 20737 2106 20789 2666
rect 20855 2106 20907 2666
rect 20973 2106 20982 2666
rect 20982 2106 21016 2666
rect 21016 2106 21025 2666
rect 21091 2106 21100 2666
rect 21100 2106 21134 2666
rect 21134 2106 21143 2666
rect 21209 2106 21218 2666
rect 21218 2106 21252 2666
rect 21252 2106 21261 2666
rect 21327 2106 21336 2666
rect 21336 2106 21370 2666
rect 21370 2106 21379 2666
rect 21445 2106 21454 2666
rect 21454 2106 21488 2666
rect 21488 2106 21497 2666
rect 21563 2106 21572 2666
rect 21572 2106 21606 2666
rect 21606 2106 21615 2666
rect 21681 2106 21690 2666
rect 21690 2106 21724 2666
rect 21724 2106 21733 2666
rect 21799 2106 21808 2666
rect 21808 2106 21842 2666
rect 21842 2106 21851 2666
rect 21917 2106 21926 2666
rect 21926 2106 21960 2666
rect 21960 2106 21969 2666
rect 22035 2106 22044 2666
rect 22044 2106 22078 2666
rect 22078 2106 22087 2666
rect 22153 2106 22162 2666
rect 22162 2106 22196 2666
rect 22196 2106 22205 2666
rect 22271 2106 22280 2666
rect 22280 2106 22314 2666
rect 22314 2106 22323 2666
rect 22389 2106 22398 2666
rect 22398 2106 22432 2666
rect 22432 2106 22441 2666
rect 22507 2106 22516 2666
rect 22516 2106 22550 2666
rect 22550 2106 22559 2666
rect 22625 2106 22634 2666
rect 22634 2106 22668 2666
rect 22668 2106 22677 2666
rect 22743 2106 22752 2666
rect 22752 2106 22786 2666
rect 22786 2106 22795 2666
rect 22861 2106 22870 2666
rect 22870 2106 22904 2666
rect 22904 2106 22913 2666
rect 22979 2106 22988 2666
rect 22988 2106 23022 2666
rect 23022 2106 23031 2666
rect 23097 2106 23106 2666
rect 23106 2106 23140 2666
rect 23140 2106 23149 2666
rect 23215 2106 23224 2666
rect 23224 2106 23258 2666
rect 23258 2106 23267 2666
rect 23333 2106 23342 2666
rect 23342 2106 23376 2666
rect 23376 2106 23385 2666
rect 23451 2106 23460 2666
rect 23460 2106 23494 2666
rect 23494 2106 23503 2666
rect 23569 2106 23578 2666
rect 23578 2106 23612 2666
rect 23612 2106 23621 2666
rect 23687 2106 23696 2666
rect 23696 2106 23730 2666
rect 23730 2106 23739 2666
rect 23895 2613 23947 2653
rect 23895 2601 23905 2613
rect 23905 2601 23939 2613
rect 23939 2601 23947 2613
rect 23975 2613 24027 2653
rect 24055 2613 24107 2653
rect 24135 2613 24187 2653
rect 24215 2613 24267 2653
rect 24295 2613 24347 2653
rect 24375 2613 24427 2653
rect 24455 2613 24507 2653
rect 24535 2613 24587 2653
rect 23975 2601 23977 2613
rect 23977 2601 24011 2613
rect 24011 2601 24027 2613
rect 24055 2601 24083 2613
rect 24083 2601 24107 2613
rect 24135 2601 24155 2613
rect 24155 2601 24187 2613
rect 24215 2601 24227 2613
rect 24227 2601 24265 2613
rect 24265 2601 24267 2613
rect 24295 2601 24299 2613
rect 24299 2601 24337 2613
rect 24337 2601 24347 2613
rect 24375 2601 24409 2613
rect 24409 2601 24427 2613
rect 24455 2601 24481 2613
rect 24481 2601 24507 2613
rect 24535 2601 24553 2613
rect 24553 2601 24587 2613
rect 24615 2613 24667 2653
rect 24615 2601 24625 2613
rect 24625 2601 24659 2613
rect 24659 2601 24667 2613
rect 24695 2601 24747 2653
rect 24775 2601 24827 2653
rect 24855 2601 24907 2653
rect 24935 2601 24987 2653
rect 25015 2601 25067 2653
rect 23895 2539 23947 2573
rect 23895 2521 23905 2539
rect 23905 2521 23939 2539
rect 23939 2521 23947 2539
rect 23975 2539 24027 2573
rect 24055 2539 24107 2573
rect 24135 2539 24187 2573
rect 24215 2539 24267 2573
rect 24295 2539 24347 2573
rect 24375 2539 24427 2573
rect 24455 2539 24507 2573
rect 24535 2539 24587 2573
rect 23975 2521 23977 2539
rect 23977 2521 24011 2539
rect 24011 2521 24027 2539
rect 24055 2521 24083 2539
rect 24083 2521 24107 2539
rect 24135 2521 24155 2539
rect 24155 2521 24187 2539
rect 24215 2521 24227 2539
rect 24227 2521 24265 2539
rect 24265 2521 24267 2539
rect 24295 2521 24299 2539
rect 24299 2521 24337 2539
rect 24337 2521 24347 2539
rect 24375 2521 24409 2539
rect 24409 2521 24427 2539
rect 24455 2521 24481 2539
rect 24481 2521 24507 2539
rect 24535 2521 24553 2539
rect 24553 2521 24587 2539
rect 24615 2539 24667 2573
rect 24615 2521 24625 2539
rect 24625 2521 24659 2539
rect 24659 2521 24667 2539
rect 24695 2521 24747 2573
rect 24775 2521 24827 2573
rect 24855 2521 24907 2573
rect 24935 2521 24987 2573
rect 25015 2521 25067 2573
rect 23895 2465 23947 2493
rect 23895 2441 23905 2465
rect 23905 2441 23939 2465
rect 23939 2441 23947 2465
rect 23975 2465 24027 2493
rect 24055 2465 24107 2493
rect 24135 2465 24187 2493
rect 24215 2465 24267 2493
rect 24295 2465 24347 2493
rect 24375 2465 24427 2493
rect 24455 2465 24507 2493
rect 24535 2465 24587 2493
rect 23975 2441 23977 2465
rect 23977 2441 24011 2465
rect 24011 2441 24027 2465
rect 24055 2441 24083 2465
rect 24083 2441 24107 2465
rect 24135 2441 24155 2465
rect 24155 2441 24187 2465
rect 24215 2441 24227 2465
rect 24227 2441 24265 2465
rect 24265 2441 24267 2465
rect 24295 2441 24299 2465
rect 24299 2441 24337 2465
rect 24337 2441 24347 2465
rect 24375 2441 24409 2465
rect 24409 2441 24427 2465
rect 24455 2441 24481 2465
rect 24481 2441 24507 2465
rect 24535 2441 24553 2465
rect 24553 2441 24587 2465
rect 24615 2465 24667 2493
rect 24615 2441 24625 2465
rect 24625 2441 24659 2465
rect 24659 2441 24667 2465
rect 24695 2441 24747 2493
rect 24775 2441 24827 2493
rect 24855 2441 24907 2493
rect 24935 2441 24987 2493
rect 25015 2441 25067 2493
rect 23895 2391 23947 2413
rect 23895 2361 23905 2391
rect 23905 2361 23939 2391
rect 23939 2361 23947 2391
rect 23975 2391 24027 2413
rect 24055 2391 24107 2413
rect 24135 2391 24187 2413
rect 24215 2391 24267 2413
rect 24295 2391 24347 2413
rect 24375 2391 24427 2413
rect 24455 2391 24507 2413
rect 24535 2391 24587 2413
rect 23975 2361 23977 2391
rect 23977 2361 24011 2391
rect 24011 2361 24027 2391
rect 24055 2361 24083 2391
rect 24083 2361 24107 2391
rect 24135 2361 24155 2391
rect 24155 2361 24187 2391
rect 24215 2361 24227 2391
rect 24227 2361 24265 2391
rect 24265 2361 24267 2391
rect 24295 2361 24299 2391
rect 24299 2361 24337 2391
rect 24337 2361 24347 2391
rect 24375 2361 24409 2391
rect 24409 2361 24427 2391
rect 24455 2361 24481 2391
rect 24481 2361 24507 2391
rect 24535 2361 24553 2391
rect 24553 2361 24587 2391
rect 24615 2391 24667 2413
rect 24615 2361 24625 2391
rect 24625 2361 24659 2391
rect 24659 2361 24667 2391
rect 24695 2361 24747 2413
rect 24775 2361 24827 2413
rect 24855 2361 24907 2413
rect 24935 2361 24987 2413
rect 25015 2361 25067 2413
rect 23895 2317 23947 2333
rect 23895 2283 23905 2317
rect 23905 2283 23939 2317
rect 23939 2283 23947 2317
rect 23895 2281 23947 2283
rect 23975 2317 24027 2333
rect 24055 2317 24107 2333
rect 24135 2317 24187 2333
rect 24215 2317 24267 2333
rect 24295 2317 24347 2333
rect 24375 2317 24427 2333
rect 24455 2317 24507 2333
rect 24535 2317 24587 2333
rect 23975 2283 23977 2317
rect 23977 2283 24011 2317
rect 24011 2283 24027 2317
rect 24055 2283 24083 2317
rect 24083 2283 24107 2317
rect 24135 2283 24155 2317
rect 24155 2283 24187 2317
rect 24215 2283 24227 2317
rect 24227 2283 24265 2317
rect 24265 2283 24267 2317
rect 24295 2283 24299 2317
rect 24299 2283 24337 2317
rect 24337 2283 24347 2317
rect 24375 2283 24409 2317
rect 24409 2283 24427 2317
rect 24455 2283 24481 2317
rect 24481 2283 24507 2317
rect 24535 2283 24553 2317
rect 24553 2283 24587 2317
rect 23975 2281 24027 2283
rect 24055 2281 24107 2283
rect 24135 2281 24187 2283
rect 24215 2281 24267 2283
rect 24295 2281 24347 2283
rect 24375 2281 24427 2283
rect 24455 2281 24507 2283
rect 24535 2281 24587 2283
rect 24615 2317 24667 2333
rect 24615 2283 24625 2317
rect 24625 2283 24659 2317
rect 24659 2283 24667 2317
rect 24615 2281 24667 2283
rect 24695 2281 24747 2333
rect 24775 2281 24827 2333
rect 24855 2281 24907 2333
rect 24935 2281 24987 2333
rect 25015 2281 25067 2333
rect 23895 2243 23947 2253
rect 23895 2209 23905 2243
rect 23905 2209 23939 2243
rect 23939 2209 23947 2243
rect 23895 2201 23947 2209
rect 23975 2243 24027 2253
rect 24055 2243 24107 2253
rect 24135 2243 24187 2253
rect 24215 2243 24267 2253
rect 24295 2243 24347 2253
rect 24375 2243 24427 2253
rect 24455 2243 24507 2253
rect 24535 2243 24587 2253
rect 23975 2209 23977 2243
rect 23977 2209 24011 2243
rect 24011 2209 24027 2243
rect 24055 2209 24083 2243
rect 24083 2209 24107 2243
rect 24135 2209 24155 2243
rect 24155 2209 24187 2243
rect 24215 2209 24227 2243
rect 24227 2209 24265 2243
rect 24265 2209 24267 2243
rect 24295 2209 24299 2243
rect 24299 2209 24337 2243
rect 24337 2209 24347 2243
rect 24375 2209 24409 2243
rect 24409 2209 24427 2243
rect 24455 2209 24481 2243
rect 24481 2209 24507 2243
rect 24535 2209 24553 2243
rect 24553 2209 24587 2243
rect 23975 2201 24027 2209
rect 24055 2201 24107 2209
rect 24135 2201 24187 2209
rect 24215 2201 24267 2209
rect 24295 2201 24347 2209
rect 24375 2201 24427 2209
rect 24455 2201 24507 2209
rect 24535 2201 24587 2209
rect 24615 2243 24667 2253
rect 24615 2209 24625 2243
rect 24625 2209 24659 2243
rect 24659 2209 24667 2243
rect 24615 2201 24667 2209
rect 24695 2201 24747 2253
rect 24775 2201 24827 2253
rect 24855 2201 24907 2253
rect 24935 2201 24987 2253
rect 25015 2201 25067 2253
rect 23895 2169 23947 2173
rect 23895 2135 23905 2169
rect 23905 2135 23939 2169
rect 23939 2135 23947 2169
rect 23895 2121 23947 2135
rect 23975 2169 24027 2173
rect 24055 2169 24107 2173
rect 24135 2169 24187 2173
rect 24215 2169 24267 2173
rect 24295 2169 24347 2173
rect 24375 2169 24427 2173
rect 24455 2169 24507 2173
rect 24535 2169 24587 2173
rect 23975 2135 23977 2169
rect 23977 2135 24011 2169
rect 24011 2135 24027 2169
rect 24055 2135 24083 2169
rect 24083 2135 24107 2169
rect 24135 2135 24155 2169
rect 24155 2135 24187 2169
rect 24215 2135 24227 2169
rect 24227 2135 24265 2169
rect 24265 2135 24267 2169
rect 24295 2135 24299 2169
rect 24299 2135 24337 2169
rect 24337 2135 24347 2169
rect 24375 2135 24409 2169
rect 24409 2135 24427 2169
rect 24455 2135 24481 2169
rect 24481 2135 24507 2169
rect 24535 2135 24553 2169
rect 24553 2135 24587 2169
rect 23975 2121 24027 2135
rect 24055 2121 24107 2135
rect 24135 2121 24187 2135
rect 24215 2121 24267 2135
rect 24295 2121 24347 2135
rect 24375 2121 24427 2135
rect 24455 2121 24507 2135
rect 24535 2121 24587 2135
rect 24615 2169 24667 2173
rect 24615 2135 24625 2169
rect 24625 2135 24659 2169
rect 24659 2135 24667 2169
rect 24615 2121 24667 2135
rect 24695 2121 24747 2173
rect 24775 2121 24827 2173
rect 24855 2121 24907 2173
rect 24935 2121 24987 2173
rect 25015 2121 25067 2173
rect 4857 2040 4915 2044
rect 4857 2006 4869 2040
rect 4869 2006 4903 2040
rect 4903 2006 4915 2040
rect 4857 1952 4915 2006
rect 4975 2040 5033 2044
rect 4975 2006 4987 2040
rect 4987 2006 5021 2040
rect 5021 2006 5033 2040
rect 4975 1952 5033 2006
rect 5093 2040 5151 2044
rect 5093 2006 5105 2040
rect 5105 2006 5139 2040
rect 5139 2006 5151 2040
rect 5093 1952 5151 2006
rect 5211 2040 5269 2044
rect 5211 2006 5223 2040
rect 5223 2006 5257 2040
rect 5257 2006 5269 2040
rect 5211 1952 5269 2006
rect 5329 2040 5387 2044
rect 5329 2006 5341 2040
rect 5341 2006 5375 2040
rect 5375 2006 5387 2040
rect 5329 1952 5387 2006
rect 5447 2040 5505 2044
rect 5447 2006 5459 2040
rect 5459 2006 5493 2040
rect 5493 2006 5505 2040
rect 5447 1952 5505 2006
rect 5565 2040 5623 2044
rect 5565 2006 5577 2040
rect 5577 2006 5611 2040
rect 5611 2006 5623 2040
rect 5565 1952 5623 2006
rect 5683 2040 5741 2044
rect 5683 2006 5695 2040
rect 5695 2006 5729 2040
rect 5729 2006 5741 2040
rect 5683 1952 5741 2006
rect 5801 2040 5859 2044
rect 5801 2006 5813 2040
rect 5813 2006 5847 2040
rect 5847 2006 5859 2040
rect 5801 1952 5859 2006
rect 5919 2040 5977 2044
rect 5919 2006 5931 2040
rect 5931 2006 5965 2040
rect 5965 2006 5977 2040
rect 5919 1952 5977 2006
rect 6037 2040 6095 2044
rect 6037 2006 6049 2040
rect 6049 2006 6083 2040
rect 6083 2006 6095 2040
rect 6037 1952 6095 2006
rect 6155 2040 6213 2044
rect 6155 2006 6167 2040
rect 6167 2006 6201 2040
rect 6201 2006 6213 2040
rect 6155 1952 6213 2006
rect 6273 2040 6331 2044
rect 6273 2006 6285 2040
rect 6285 2006 6319 2040
rect 6319 2006 6331 2040
rect 6273 1952 6331 2006
rect 6391 2040 6449 2044
rect 6391 2006 6403 2040
rect 6403 2006 6437 2040
rect 6437 2006 6449 2040
rect 6391 1952 6449 2006
rect 6509 2040 6567 2044
rect 6509 2006 6521 2040
rect 6521 2006 6555 2040
rect 6555 2006 6567 2040
rect 6509 1952 6567 2006
rect 6855 1952 6913 2044
rect 6973 1952 7031 2044
rect 7091 2040 7149 2044
rect 7091 2006 7103 2040
rect 7103 2006 7137 2040
rect 7137 2006 7149 2040
rect 7091 1952 7149 2006
rect 7209 2040 7267 2044
rect 7209 2006 7221 2040
rect 7221 2006 7255 2040
rect 7255 2006 7267 2040
rect 7209 1952 7267 2006
rect 7327 2040 7385 2044
rect 7327 2006 7339 2040
rect 7339 2006 7373 2040
rect 7373 2006 7385 2040
rect 7327 1952 7385 2006
rect 7445 2040 7503 2044
rect 7445 2006 7457 2040
rect 7457 2006 7491 2040
rect 7491 2006 7503 2040
rect 7445 1952 7503 2006
rect 7563 2040 7621 2044
rect 7563 2006 7575 2040
rect 7575 2006 7609 2040
rect 7609 2006 7621 2040
rect 7563 1952 7621 2006
rect 7681 2040 7739 2044
rect 7681 2006 7693 2040
rect 7693 2006 7727 2040
rect 7727 2006 7739 2040
rect 7681 1952 7739 2006
rect 7799 2040 7857 2044
rect 7799 2006 7811 2040
rect 7811 2006 7845 2040
rect 7845 2006 7857 2040
rect 7799 1952 7857 2006
rect 7917 2040 7975 2044
rect 7917 2006 7929 2040
rect 7929 2006 7963 2040
rect 7963 2006 7975 2040
rect 7917 1952 7975 2006
rect 8035 2040 8093 2044
rect 8035 2006 8047 2040
rect 8047 2006 8081 2040
rect 8081 2006 8093 2040
rect 8035 1952 8093 2006
rect 8153 2040 8211 2044
rect 8153 2006 8165 2040
rect 8165 2006 8199 2040
rect 8199 2006 8211 2040
rect 8153 1952 8211 2006
rect 8271 2040 8329 2044
rect 8271 2006 8283 2040
rect 8283 2006 8317 2040
rect 8317 2006 8329 2040
rect 8271 1952 8329 2006
rect 8389 2040 8447 2044
rect 8389 2006 8401 2040
rect 8401 2006 8435 2040
rect 8435 2006 8447 2040
rect 8389 1952 8447 2006
rect 8507 2040 8565 2044
rect 8507 2006 8519 2040
rect 8519 2006 8553 2040
rect 8553 2006 8565 2040
rect 8507 1952 8565 2006
rect 8853 2040 8911 2044
rect 8853 2006 8865 2040
rect 8865 2006 8899 2040
rect 8899 2006 8911 2040
rect 8853 1952 8911 2006
rect 8971 2040 9029 2044
rect 8971 2006 8983 2040
rect 8983 2006 9017 2040
rect 9017 2006 9029 2040
rect 8971 1952 9029 2006
rect 9089 2040 9147 2044
rect 9089 2006 9101 2040
rect 9101 2006 9135 2040
rect 9135 2006 9147 2040
rect 9089 1952 9147 2006
rect 9207 2040 9265 2044
rect 9207 2006 9219 2040
rect 9219 2006 9253 2040
rect 9253 2006 9265 2040
rect 9207 1952 9265 2006
rect 9325 2040 9383 2044
rect 9325 2006 9337 2040
rect 9337 2006 9371 2040
rect 9371 2006 9383 2040
rect 9325 1952 9383 2006
rect 9443 2040 9501 2044
rect 9443 2006 9455 2040
rect 9455 2006 9489 2040
rect 9489 2006 9501 2040
rect 9443 1952 9501 2006
rect 9561 2040 9619 2044
rect 9561 2006 9573 2040
rect 9573 2006 9607 2040
rect 9607 2006 9619 2040
rect 9561 1952 9619 2006
rect 9679 2040 9737 2044
rect 9679 2006 9691 2040
rect 9691 2006 9725 2040
rect 9725 2006 9737 2040
rect 9679 1952 9737 2006
rect 9797 2040 9855 2044
rect 9797 2006 9809 2040
rect 9809 2006 9843 2040
rect 9843 2006 9855 2040
rect 9797 1952 9855 2006
rect 9915 2040 9973 2044
rect 9915 2006 9927 2040
rect 9927 2006 9961 2040
rect 9961 2006 9973 2040
rect 9915 1952 9973 2006
rect 10033 2040 10091 2044
rect 10033 2006 10045 2040
rect 10045 2006 10079 2040
rect 10079 2006 10091 2040
rect 10033 1952 10091 2006
rect 10151 2040 10209 2044
rect 10151 2006 10163 2040
rect 10163 2006 10197 2040
rect 10197 2006 10209 2040
rect 10151 1952 10209 2006
rect 10269 2040 10327 2044
rect 10269 2006 10281 2040
rect 10281 2006 10315 2040
rect 10315 2006 10327 2040
rect 10269 1952 10327 2006
rect 10387 2040 10445 2044
rect 10387 2006 10399 2040
rect 10399 2006 10433 2040
rect 10433 2006 10445 2040
rect 10387 1952 10445 2006
rect 10505 2040 10563 2044
rect 10505 2006 10517 2040
rect 10517 2006 10551 2040
rect 10551 2006 10563 2040
rect 10505 1952 10563 2006
rect 12547 1891 12605 2045
rect 12665 2039 12723 2045
rect 12665 2005 12677 2039
rect 12677 2005 12711 2039
rect 12711 2005 12723 2039
rect 12665 1931 12723 2005
rect 12665 1897 12677 1931
rect 12677 1897 12711 1931
rect 12711 1897 12723 1931
rect 12665 1891 12723 1897
rect 12783 2039 12841 2045
rect 12783 2005 12795 2039
rect 12795 2005 12829 2039
rect 12829 2005 12841 2039
rect 12783 1931 12841 2005
rect 12783 1897 12795 1931
rect 12795 1897 12829 1931
rect 12829 1897 12841 1931
rect 12783 1891 12841 1897
rect 12901 2039 12959 2045
rect 12901 2005 12913 2039
rect 12913 2005 12947 2039
rect 12947 2005 12959 2039
rect 12901 1931 12959 2005
rect 12901 1897 12913 1931
rect 12913 1897 12947 1931
rect 12947 1897 12959 1931
rect 12901 1891 12959 1897
rect 13019 2039 13077 2045
rect 13019 2005 13031 2039
rect 13031 2005 13065 2039
rect 13065 2005 13077 2039
rect 13019 1931 13077 2005
rect 13019 1897 13031 1931
rect 13031 1897 13065 1931
rect 13065 1897 13077 1931
rect 13019 1891 13077 1897
rect 13137 2039 13195 2045
rect 13137 2005 13149 2039
rect 13149 2005 13183 2039
rect 13183 2005 13195 2039
rect 13137 1931 13195 2005
rect 13137 1897 13149 1931
rect 13149 1897 13183 1931
rect 13183 1897 13195 1931
rect 13137 1891 13195 1897
rect 13255 2039 13313 2045
rect 13255 2005 13267 2039
rect 13267 2005 13301 2039
rect 13301 2005 13313 2039
rect 13255 1931 13313 2005
rect 13255 1897 13267 1931
rect 13267 1897 13301 1931
rect 13301 1897 13313 1931
rect 13255 1891 13313 1897
rect 13373 2039 13431 2045
rect 13373 2005 13385 2039
rect 13385 2005 13419 2039
rect 13419 2005 13431 2039
rect 13373 1931 13431 2005
rect 13373 1897 13385 1931
rect 13385 1897 13419 1931
rect 13419 1897 13431 1931
rect 13373 1891 13431 1897
rect 13491 2039 13549 2045
rect 13491 2005 13503 2039
rect 13503 2005 13537 2039
rect 13537 2005 13549 2039
rect 13491 1931 13549 2005
rect 13491 1897 13503 1931
rect 13503 1897 13537 1931
rect 13537 1897 13549 1931
rect 13491 1891 13549 1897
rect 13609 2039 13667 2045
rect 13609 2005 13621 2039
rect 13621 2005 13655 2039
rect 13655 2005 13667 2039
rect 13609 1931 13667 2005
rect 13609 1897 13621 1931
rect 13621 1897 13655 1931
rect 13655 1897 13667 1931
rect 13609 1891 13667 1897
rect 13727 2039 13785 2045
rect 13727 2005 13739 2039
rect 13739 2005 13773 2039
rect 13773 2005 13785 2039
rect 13727 1931 13785 2005
rect 13727 1897 13739 1931
rect 13739 1897 13773 1931
rect 13773 1897 13785 1931
rect 13727 1891 13785 1897
rect 13845 2039 13903 2045
rect 13845 2005 13857 2039
rect 13857 2005 13891 2039
rect 13891 2005 13903 2039
rect 13845 1931 13903 2005
rect 13845 1897 13857 1931
rect 13857 1897 13891 1931
rect 13891 1897 13903 1931
rect 13845 1891 13903 1897
rect 13963 2039 14021 2045
rect 13963 2005 13975 2039
rect 13975 2005 14009 2039
rect 14009 2005 14021 2039
rect 13963 1931 14021 2005
rect 13963 1897 13975 1931
rect 13975 1897 14009 1931
rect 14009 1897 14021 1931
rect 13963 1891 14021 1897
rect 14081 2039 14139 2045
rect 14081 2005 14093 2039
rect 14093 2005 14127 2039
rect 14127 2005 14139 2039
rect 14081 1931 14139 2005
rect 14081 1897 14093 1931
rect 14093 1897 14127 1931
rect 14127 1897 14139 1931
rect 14081 1891 14139 1897
rect 14199 2039 14257 2045
rect 14199 2005 14211 2039
rect 14211 2005 14245 2039
rect 14245 2005 14257 2039
rect 14199 1931 14257 2005
rect 14199 1897 14211 1931
rect 14211 1897 14245 1931
rect 14245 1897 14257 1931
rect 14199 1891 14257 1897
rect 14317 2039 14375 2045
rect 14317 2005 14329 2039
rect 14329 2005 14363 2039
rect 14363 2005 14375 2039
rect 14317 1931 14375 2005
rect 14317 1897 14329 1931
rect 14329 1897 14363 1931
rect 14363 1897 14375 1931
rect 14317 1891 14375 1897
rect 14435 2039 14493 2045
rect 14435 2005 14447 2039
rect 14447 2005 14481 2039
rect 14481 2005 14493 2039
rect 14435 1931 14493 2005
rect 14435 1897 14447 1931
rect 14447 1897 14481 1931
rect 14481 1897 14493 1931
rect 14435 1891 14493 1897
rect 14553 2039 14611 2045
rect 14553 2005 14565 2039
rect 14565 2005 14599 2039
rect 14599 2005 14611 2039
rect 14553 1931 14611 2005
rect 14553 1897 14565 1931
rect 14565 1897 14599 1931
rect 14599 1897 14611 1931
rect 14553 1891 14611 1897
rect 14671 2039 14729 2045
rect 14671 2005 14683 2039
rect 14683 2005 14717 2039
rect 14717 2005 14729 2039
rect 14671 1931 14729 2005
rect 14671 1897 14683 1931
rect 14683 1897 14717 1931
rect 14717 1897 14729 1931
rect 14671 1891 14729 1897
rect 14789 2039 14847 2045
rect 14789 2005 14801 2039
rect 14801 2005 14835 2039
rect 14835 2005 14847 2039
rect 14789 1931 14847 2005
rect 14789 1897 14801 1931
rect 14801 1897 14835 1931
rect 14835 1897 14847 1931
rect 14789 1891 14847 1897
rect 14907 2039 14965 2045
rect 14907 2005 14919 2039
rect 14919 2005 14953 2039
rect 14953 2005 14965 2039
rect 14907 1931 14965 2005
rect 14907 1897 14919 1931
rect 14919 1897 14953 1931
rect 14953 1897 14965 1931
rect 14907 1891 14965 1897
rect 15025 2039 15083 2045
rect 15025 2005 15037 2039
rect 15037 2005 15071 2039
rect 15071 2005 15083 2039
rect 15025 1931 15083 2005
rect 15025 1897 15037 1931
rect 15037 1897 15071 1931
rect 15071 1897 15083 1931
rect 15025 1891 15083 1897
rect 15143 2039 15201 2045
rect 15143 2005 15155 2039
rect 15155 2005 15189 2039
rect 15189 2005 15201 2039
rect 15143 1931 15201 2005
rect 15143 1897 15155 1931
rect 15155 1897 15189 1931
rect 15189 1897 15201 1931
rect 15143 1891 15201 1897
rect 15261 2039 15319 2045
rect 15261 2005 15273 2039
rect 15273 2005 15307 2039
rect 15307 2005 15319 2039
rect 15261 1931 15319 2005
rect 15261 1897 15273 1931
rect 15273 1897 15307 1931
rect 15307 1897 15319 1931
rect 15261 1891 15319 1897
rect 15379 2039 15437 2045
rect 15379 2005 15391 2039
rect 15391 2005 15425 2039
rect 15425 2005 15437 2039
rect 15379 1931 15437 2005
rect 15379 1897 15391 1931
rect 15391 1897 15425 1931
rect 15425 1897 15437 1931
rect 15379 1891 15437 1897
rect 16670 1891 16728 2045
rect 16788 2039 16846 2045
rect 16788 2005 16800 2039
rect 16800 2005 16834 2039
rect 16834 2005 16846 2039
rect 16788 1931 16846 2005
rect 16788 1897 16800 1931
rect 16800 1897 16834 1931
rect 16834 1897 16846 1931
rect 16788 1891 16846 1897
rect 16906 2039 16964 2045
rect 16906 2005 16918 2039
rect 16918 2005 16952 2039
rect 16952 2005 16964 2039
rect 16906 1931 16964 2005
rect 16906 1897 16918 1931
rect 16918 1897 16952 1931
rect 16952 1897 16964 1931
rect 16906 1891 16964 1897
rect 17024 2039 17082 2045
rect 17024 2005 17036 2039
rect 17036 2005 17070 2039
rect 17070 2005 17082 2039
rect 17024 1931 17082 2005
rect 17024 1897 17036 1931
rect 17036 1897 17070 1931
rect 17070 1897 17082 1931
rect 17024 1891 17082 1897
rect 17142 2039 17200 2045
rect 17142 2005 17154 2039
rect 17154 2005 17188 2039
rect 17188 2005 17200 2039
rect 17142 1931 17200 2005
rect 17142 1897 17154 1931
rect 17154 1897 17188 1931
rect 17188 1897 17200 1931
rect 17142 1891 17200 1897
rect 17260 2039 17318 2045
rect 17260 2005 17272 2039
rect 17272 2005 17306 2039
rect 17306 2005 17318 2039
rect 17260 1931 17318 2005
rect 17260 1897 17272 1931
rect 17272 1897 17306 1931
rect 17306 1897 17318 1931
rect 17260 1891 17318 1897
rect 17378 2039 17436 2045
rect 17378 2005 17390 2039
rect 17390 2005 17424 2039
rect 17424 2005 17436 2039
rect 17378 1931 17436 2005
rect 17378 1897 17390 1931
rect 17390 1897 17424 1931
rect 17424 1897 17436 1931
rect 17378 1891 17436 1897
rect 17496 2039 17554 2045
rect 17496 2005 17508 2039
rect 17508 2005 17542 2039
rect 17542 2005 17554 2039
rect 17496 1931 17554 2005
rect 17496 1897 17508 1931
rect 17508 1897 17542 1931
rect 17542 1897 17554 1931
rect 17496 1891 17554 1897
rect 17614 2039 17672 2045
rect 17614 2005 17626 2039
rect 17626 2005 17660 2039
rect 17660 2005 17672 2039
rect 17614 1931 17672 2005
rect 17614 1897 17626 1931
rect 17626 1897 17660 1931
rect 17660 1897 17672 1931
rect 17614 1891 17672 1897
rect 17732 2039 17790 2045
rect 17732 2005 17744 2039
rect 17744 2005 17778 2039
rect 17778 2005 17790 2039
rect 17732 1931 17790 2005
rect 17732 1897 17744 1931
rect 17744 1897 17778 1931
rect 17778 1897 17790 1931
rect 17732 1891 17790 1897
rect 17850 2039 17908 2045
rect 17850 2005 17862 2039
rect 17862 2005 17896 2039
rect 17896 2005 17908 2039
rect 17850 1931 17908 2005
rect 17850 1897 17862 1931
rect 17862 1897 17896 1931
rect 17896 1897 17908 1931
rect 17850 1891 17908 1897
rect 17968 2039 18026 2045
rect 17968 2005 17980 2039
rect 17980 2005 18014 2039
rect 18014 2005 18026 2039
rect 17968 1931 18026 2005
rect 17968 1897 17980 1931
rect 17980 1897 18014 1931
rect 18014 1897 18026 1931
rect 17968 1891 18026 1897
rect 18086 2039 18144 2045
rect 18086 2005 18098 2039
rect 18098 2005 18132 2039
rect 18132 2005 18144 2039
rect 18086 1931 18144 2005
rect 18086 1897 18098 1931
rect 18098 1897 18132 1931
rect 18132 1897 18144 1931
rect 18086 1891 18144 1897
rect 18204 2039 18262 2045
rect 18204 2005 18216 2039
rect 18216 2005 18250 2039
rect 18250 2005 18262 2039
rect 18204 1931 18262 2005
rect 18204 1897 18216 1931
rect 18216 1897 18250 1931
rect 18250 1897 18262 1931
rect 18204 1891 18262 1897
rect 18322 2039 18380 2045
rect 18322 2005 18334 2039
rect 18334 2005 18368 2039
rect 18368 2005 18380 2039
rect 18322 1931 18380 2005
rect 18322 1897 18334 1931
rect 18334 1897 18368 1931
rect 18368 1897 18380 1931
rect 18322 1891 18380 1897
rect 18440 2039 18498 2045
rect 18440 2005 18452 2039
rect 18452 2005 18486 2039
rect 18486 2005 18498 2039
rect 18440 1931 18498 2005
rect 18440 1897 18452 1931
rect 18452 1897 18486 1931
rect 18486 1897 18498 1931
rect 18440 1891 18498 1897
rect 18558 2039 18616 2045
rect 18558 2005 18570 2039
rect 18570 2005 18604 2039
rect 18604 2005 18616 2039
rect 18558 1931 18616 2005
rect 18558 1897 18570 1931
rect 18570 1897 18604 1931
rect 18604 1897 18616 1931
rect 18558 1891 18616 1897
rect 18676 2039 18734 2045
rect 18676 2005 18688 2039
rect 18688 2005 18722 2039
rect 18722 2005 18734 2039
rect 18676 1931 18734 2005
rect 18676 1897 18688 1931
rect 18688 1897 18722 1931
rect 18722 1897 18734 1931
rect 18676 1891 18734 1897
rect 18794 2039 18852 2045
rect 18794 2005 18806 2039
rect 18806 2005 18840 2039
rect 18840 2005 18852 2039
rect 18794 1931 18852 2005
rect 18794 1897 18806 1931
rect 18806 1897 18840 1931
rect 18840 1897 18852 1931
rect 18794 1891 18852 1897
rect 18912 2039 18970 2045
rect 18912 2005 18924 2039
rect 18924 2005 18958 2039
rect 18958 2005 18970 2039
rect 18912 1931 18970 2005
rect 18912 1897 18924 1931
rect 18924 1897 18958 1931
rect 18958 1897 18970 1931
rect 18912 1891 18970 1897
rect 19030 2039 19088 2045
rect 19030 2005 19042 2039
rect 19042 2005 19076 2039
rect 19076 2005 19088 2039
rect 19030 1931 19088 2005
rect 19030 1897 19042 1931
rect 19042 1897 19076 1931
rect 19076 1897 19088 1931
rect 19030 1891 19088 1897
rect 19148 2039 19206 2045
rect 19148 2005 19160 2039
rect 19160 2005 19194 2039
rect 19194 2005 19206 2039
rect 19148 1931 19206 2005
rect 19148 1897 19160 1931
rect 19160 1897 19194 1931
rect 19194 1897 19206 1931
rect 19148 1891 19206 1897
rect 19266 2039 19324 2045
rect 19266 2005 19278 2039
rect 19278 2005 19312 2039
rect 19312 2005 19324 2039
rect 19266 1931 19324 2005
rect 19266 1897 19278 1931
rect 19278 1897 19312 1931
rect 19312 1897 19324 1931
rect 19266 1891 19324 1897
rect 19384 2039 19442 2045
rect 19384 2005 19396 2039
rect 19396 2005 19430 2039
rect 19430 2005 19442 2039
rect 19384 1931 19442 2005
rect 19384 1897 19396 1931
rect 19396 1897 19430 1931
rect 19430 1897 19442 1931
rect 19384 1891 19442 1897
rect 19502 2039 19560 2045
rect 19502 2005 19514 2039
rect 19514 2005 19548 2039
rect 19548 2005 19560 2039
rect 19502 1931 19560 2005
rect 19502 1897 19514 1931
rect 19514 1897 19548 1931
rect 19548 1897 19560 1931
rect 19502 1891 19560 1897
rect 20793 1891 20851 2045
rect 20911 2039 20969 2045
rect 20911 2005 20923 2039
rect 20923 2005 20957 2039
rect 20957 2005 20969 2039
rect 20911 1931 20969 2005
rect 20911 1897 20923 1931
rect 20923 1897 20957 1931
rect 20957 1897 20969 1931
rect 20911 1891 20969 1897
rect 21029 2039 21087 2045
rect 21029 2005 21041 2039
rect 21041 2005 21075 2039
rect 21075 2005 21087 2039
rect 21029 1931 21087 2005
rect 21029 1897 21041 1931
rect 21041 1897 21075 1931
rect 21075 1897 21087 1931
rect 21029 1891 21087 1897
rect 21147 2039 21205 2045
rect 21147 2005 21159 2039
rect 21159 2005 21193 2039
rect 21193 2005 21205 2039
rect 21147 1931 21205 2005
rect 21147 1897 21159 1931
rect 21159 1897 21193 1931
rect 21193 1897 21205 1931
rect 21147 1891 21205 1897
rect 21265 2039 21323 2045
rect 21265 2005 21277 2039
rect 21277 2005 21311 2039
rect 21311 2005 21323 2039
rect 21265 1931 21323 2005
rect 21265 1897 21277 1931
rect 21277 1897 21311 1931
rect 21311 1897 21323 1931
rect 21265 1891 21323 1897
rect 21383 2039 21441 2045
rect 21383 2005 21395 2039
rect 21395 2005 21429 2039
rect 21429 2005 21441 2039
rect 21383 1931 21441 2005
rect 21383 1897 21395 1931
rect 21395 1897 21429 1931
rect 21429 1897 21441 1931
rect 21383 1891 21441 1897
rect 21501 2039 21559 2045
rect 21501 2005 21513 2039
rect 21513 2005 21547 2039
rect 21547 2005 21559 2039
rect 21501 1931 21559 2005
rect 21501 1897 21513 1931
rect 21513 1897 21547 1931
rect 21547 1897 21559 1931
rect 21501 1891 21559 1897
rect 21619 2039 21677 2045
rect 21619 2005 21631 2039
rect 21631 2005 21665 2039
rect 21665 2005 21677 2039
rect 21619 1931 21677 2005
rect 21619 1897 21631 1931
rect 21631 1897 21665 1931
rect 21665 1897 21677 1931
rect 21619 1891 21677 1897
rect 21737 2039 21795 2045
rect 21737 2005 21749 2039
rect 21749 2005 21783 2039
rect 21783 2005 21795 2039
rect 21737 1931 21795 2005
rect 21737 1897 21749 1931
rect 21749 1897 21783 1931
rect 21783 1897 21795 1931
rect 21737 1891 21795 1897
rect 21855 2039 21913 2045
rect 21855 2005 21867 2039
rect 21867 2005 21901 2039
rect 21901 2005 21913 2039
rect 21855 1931 21913 2005
rect 21855 1897 21867 1931
rect 21867 1897 21901 1931
rect 21901 1897 21913 1931
rect 21855 1891 21913 1897
rect 21973 2039 22031 2045
rect 21973 2005 21985 2039
rect 21985 2005 22019 2039
rect 22019 2005 22031 2039
rect 21973 1931 22031 2005
rect 21973 1897 21985 1931
rect 21985 1897 22019 1931
rect 22019 1897 22031 1931
rect 21973 1891 22031 1897
rect 22091 2039 22149 2045
rect 22091 2005 22103 2039
rect 22103 2005 22137 2039
rect 22137 2005 22149 2039
rect 22091 1931 22149 2005
rect 22091 1897 22103 1931
rect 22103 1897 22137 1931
rect 22137 1897 22149 1931
rect 22091 1891 22149 1897
rect 22209 2039 22267 2045
rect 22209 2005 22221 2039
rect 22221 2005 22255 2039
rect 22255 2005 22267 2039
rect 22209 1931 22267 2005
rect 22209 1897 22221 1931
rect 22221 1897 22255 1931
rect 22255 1897 22267 1931
rect 22209 1891 22267 1897
rect 22327 2039 22385 2045
rect 22327 2005 22339 2039
rect 22339 2005 22373 2039
rect 22373 2005 22385 2039
rect 22327 1931 22385 2005
rect 22327 1897 22339 1931
rect 22339 1897 22373 1931
rect 22373 1897 22385 1931
rect 22327 1891 22385 1897
rect 22445 2039 22503 2045
rect 22445 2005 22457 2039
rect 22457 2005 22491 2039
rect 22491 2005 22503 2039
rect 22445 1931 22503 2005
rect 22445 1897 22457 1931
rect 22457 1897 22491 1931
rect 22491 1897 22503 1931
rect 22445 1891 22503 1897
rect 22563 2039 22621 2045
rect 22563 2005 22575 2039
rect 22575 2005 22609 2039
rect 22609 2005 22621 2039
rect 22563 1931 22621 2005
rect 22563 1897 22575 1931
rect 22575 1897 22609 1931
rect 22609 1897 22621 1931
rect 22563 1891 22621 1897
rect 22681 2039 22739 2045
rect 22681 2005 22693 2039
rect 22693 2005 22727 2039
rect 22727 2005 22739 2039
rect 22681 1931 22739 2005
rect 22681 1897 22693 1931
rect 22693 1897 22727 1931
rect 22727 1897 22739 1931
rect 22681 1891 22739 1897
rect 22799 2039 22857 2045
rect 22799 2005 22811 2039
rect 22811 2005 22845 2039
rect 22845 2005 22857 2039
rect 22799 1931 22857 2005
rect 22799 1897 22811 1931
rect 22811 1897 22845 1931
rect 22845 1897 22857 1931
rect 22799 1891 22857 1897
rect 22917 2039 22975 2045
rect 22917 2005 22929 2039
rect 22929 2005 22963 2039
rect 22963 2005 22975 2039
rect 22917 1931 22975 2005
rect 22917 1897 22929 1931
rect 22929 1897 22963 1931
rect 22963 1897 22975 1931
rect 22917 1891 22975 1897
rect 23035 2039 23093 2045
rect 23035 2005 23047 2039
rect 23047 2005 23081 2039
rect 23081 2005 23093 2039
rect 23035 1931 23093 2005
rect 23035 1897 23047 1931
rect 23047 1897 23081 1931
rect 23081 1897 23093 1931
rect 23035 1891 23093 1897
rect 23153 2039 23211 2045
rect 23153 2005 23165 2039
rect 23165 2005 23199 2039
rect 23199 2005 23211 2039
rect 23153 1931 23211 2005
rect 23153 1897 23165 1931
rect 23165 1897 23199 1931
rect 23199 1897 23211 1931
rect 23153 1891 23211 1897
rect 23271 2039 23329 2045
rect 23271 2005 23283 2039
rect 23283 2005 23317 2039
rect 23317 2005 23329 2039
rect 23271 1931 23329 2005
rect 23271 1897 23283 1931
rect 23283 1897 23317 1931
rect 23317 1897 23329 1931
rect 23271 1891 23329 1897
rect 23389 2039 23447 2045
rect 23389 2005 23401 2039
rect 23401 2005 23435 2039
rect 23435 2005 23447 2039
rect 23389 1931 23447 2005
rect 23389 1897 23401 1931
rect 23401 1897 23435 1931
rect 23435 1897 23447 1931
rect 23389 1891 23447 1897
rect 23507 2039 23565 2045
rect 23507 2005 23519 2039
rect 23519 2005 23553 2039
rect 23553 2005 23565 2039
rect 23507 1931 23565 2005
rect 23507 1897 23519 1931
rect 23519 1897 23553 1931
rect 23553 1897 23565 1931
rect 23507 1891 23565 1897
rect 23625 2039 23683 2045
rect 23625 2005 23637 2039
rect 23637 2005 23671 2039
rect 23671 2005 23683 2039
rect 23625 1931 23683 2005
rect 23625 1897 23637 1931
rect 23637 1897 23671 1931
rect 23671 1897 23683 1931
rect 23625 1891 23683 1897
rect 23895 2061 23905 2093
rect 23905 2061 23939 2093
rect 23939 2061 23947 2093
rect 23895 2041 23947 2061
rect 23975 2061 23977 2093
rect 23977 2061 24011 2093
rect 24011 2061 24027 2093
rect 24055 2061 24083 2093
rect 24083 2061 24107 2093
rect 24135 2061 24155 2093
rect 24155 2061 24187 2093
rect 24215 2061 24227 2093
rect 24227 2061 24265 2093
rect 24265 2061 24267 2093
rect 24295 2061 24299 2093
rect 24299 2061 24337 2093
rect 24337 2061 24347 2093
rect 24375 2061 24409 2093
rect 24409 2061 24427 2093
rect 24455 2061 24481 2093
rect 24481 2061 24507 2093
rect 24535 2061 24553 2093
rect 24553 2061 24587 2093
rect 23975 2041 24027 2061
rect 24055 2041 24107 2061
rect 24135 2041 24187 2061
rect 24215 2041 24267 2061
rect 24295 2041 24347 2061
rect 24375 2041 24427 2061
rect 24455 2041 24507 2061
rect 24535 2041 24587 2061
rect 24615 2061 24625 2093
rect 24625 2061 24659 2093
rect 24659 2061 24667 2093
rect 24615 2041 24667 2061
rect 24695 2041 24747 2093
rect 24775 2041 24827 2093
rect 24855 2041 24907 2093
rect 24935 2041 24987 2093
rect 25015 2041 25067 2093
rect 23895 1987 23905 2013
rect 23905 1987 23939 2013
rect 23939 1987 23947 2013
rect 23895 1961 23947 1987
rect 23975 1987 23977 2013
rect 23977 1987 24011 2013
rect 24011 1987 24027 2013
rect 24055 1987 24083 2013
rect 24083 1987 24107 2013
rect 24135 1987 24155 2013
rect 24155 1987 24187 2013
rect 24215 1987 24227 2013
rect 24227 1987 24265 2013
rect 24265 1987 24267 2013
rect 24295 1987 24299 2013
rect 24299 1987 24337 2013
rect 24337 1987 24347 2013
rect 24375 1987 24409 2013
rect 24409 1987 24427 2013
rect 24455 1987 24481 2013
rect 24481 1987 24507 2013
rect 24535 1987 24553 2013
rect 24553 1987 24587 2013
rect 23975 1961 24027 1987
rect 24055 1961 24107 1987
rect 24135 1961 24187 1987
rect 24215 1961 24267 1987
rect 24295 1961 24347 1987
rect 24375 1961 24427 1987
rect 24455 1961 24507 1987
rect 24535 1961 24587 1987
rect 24615 1987 24625 2013
rect 24625 1987 24659 2013
rect 24659 1987 24667 2013
rect 24615 1961 24667 1987
rect 24695 1961 24747 2013
rect 24775 1961 24827 2013
rect 24855 1961 24907 2013
rect 24935 1961 24987 2013
rect 25015 1961 25067 2013
rect 4801 1319 4853 1569
rect 5037 1319 5089 1569
rect 5273 1319 5325 1569
rect 5509 1319 5561 1569
rect 5745 1319 5797 1569
rect 5981 1319 6033 1569
rect 6217 1319 6269 1569
rect 6453 1319 6505 1569
rect 6689 1319 6741 1569
rect 6925 1319 6977 1569
rect 7161 1319 7213 1569
rect 7397 1319 7449 1569
rect 7633 1319 7685 1569
rect 7869 1319 7921 1569
rect 8105 1319 8157 1569
rect 8341 1319 8393 1569
rect 8577 1319 8629 1569
rect 8813 1319 8865 1569
rect 9049 1319 9101 1569
rect 9285 1319 9337 1569
rect 9521 1319 9573 1569
rect 9757 1319 9809 1569
rect 9993 1319 10045 1569
rect 10229 1319 10281 1569
rect 10465 1319 10517 1569
rect 10701 1319 10753 1569
rect 12491 1270 12500 1830
rect 12500 1270 12534 1830
rect 12534 1270 12543 1830
rect 12609 1270 12618 1830
rect 12618 1270 12652 1830
rect 12652 1270 12661 1830
rect 12727 1270 12736 1830
rect 12736 1270 12770 1830
rect 12770 1270 12779 1830
rect 12845 1270 12854 1830
rect 12854 1270 12888 1830
rect 12888 1270 12897 1830
rect 12963 1270 12972 1830
rect 12972 1270 13006 1830
rect 13006 1270 13015 1830
rect 13081 1270 13090 1830
rect 13090 1270 13124 1830
rect 13124 1270 13133 1830
rect 13199 1270 13208 1830
rect 13208 1270 13242 1830
rect 13242 1270 13251 1830
rect 13317 1270 13326 1830
rect 13326 1270 13360 1830
rect 13360 1270 13369 1830
rect 13435 1270 13444 1830
rect 13444 1270 13478 1830
rect 13478 1270 13487 1830
rect 13553 1270 13562 1830
rect 13562 1270 13596 1830
rect 13596 1270 13605 1830
rect 13671 1270 13680 1830
rect 13680 1270 13714 1830
rect 13714 1270 13723 1830
rect 13789 1270 13798 1830
rect 13798 1270 13832 1830
rect 13832 1270 13841 1830
rect 13907 1270 13916 1830
rect 13916 1270 13950 1830
rect 13950 1270 13959 1830
rect 14025 1270 14034 1830
rect 14034 1270 14068 1830
rect 14068 1270 14077 1830
rect 14143 1270 14152 1830
rect 14152 1270 14186 1830
rect 14186 1270 14195 1830
rect 14261 1270 14270 1830
rect 14270 1270 14304 1830
rect 14304 1270 14313 1830
rect 14379 1270 14388 1830
rect 14388 1270 14422 1830
rect 14422 1270 14431 1830
rect 14497 1270 14506 1830
rect 14506 1270 14540 1830
rect 14540 1270 14549 1830
rect 14615 1270 14624 1830
rect 14624 1270 14658 1830
rect 14658 1270 14667 1830
rect 14733 1270 14742 1830
rect 14742 1270 14776 1830
rect 14776 1270 14785 1830
rect 14851 1270 14860 1830
rect 14860 1270 14894 1830
rect 14894 1270 14903 1830
rect 14969 1270 14978 1830
rect 14978 1270 15012 1830
rect 15012 1270 15021 1830
rect 15087 1270 15096 1830
rect 15096 1270 15130 1830
rect 15130 1270 15139 1830
rect 15205 1270 15214 1830
rect 15214 1270 15248 1830
rect 15248 1270 15257 1830
rect 15323 1270 15332 1830
rect 15332 1270 15366 1830
rect 15366 1270 15375 1830
rect 15441 1270 15450 1830
rect 15450 1270 15484 1830
rect 15484 1270 15493 1830
rect 23895 1913 23905 1933
rect 23905 1913 23939 1933
rect 23939 1913 23947 1933
rect 23895 1881 23947 1913
rect 23975 1913 23977 1933
rect 23977 1913 24011 1933
rect 24011 1913 24027 1933
rect 24055 1913 24083 1933
rect 24083 1913 24107 1933
rect 24135 1913 24155 1933
rect 24155 1913 24187 1933
rect 24215 1913 24227 1933
rect 24227 1913 24265 1933
rect 24265 1913 24267 1933
rect 24295 1913 24299 1933
rect 24299 1913 24337 1933
rect 24337 1913 24347 1933
rect 24375 1913 24409 1933
rect 24409 1913 24427 1933
rect 24455 1913 24481 1933
rect 24481 1913 24507 1933
rect 24535 1913 24553 1933
rect 24553 1913 24587 1933
rect 23975 1881 24027 1913
rect 24055 1881 24107 1913
rect 24135 1881 24187 1913
rect 24215 1881 24267 1913
rect 24295 1881 24347 1913
rect 24375 1881 24427 1913
rect 24455 1881 24507 1913
rect 24535 1881 24587 1913
rect 24615 1913 24625 1933
rect 24625 1913 24659 1933
rect 24659 1913 24667 1933
rect 24615 1881 24667 1913
rect 24695 1881 24747 1933
rect 24775 1881 24827 1933
rect 24855 1881 24907 1933
rect 24935 1881 24987 1933
rect 25015 1881 25067 1933
rect 16614 1270 16623 1830
rect 16623 1270 16657 1830
rect 16657 1270 16666 1830
rect 16732 1270 16741 1830
rect 16741 1270 16775 1830
rect 16775 1270 16784 1830
rect 16850 1270 16859 1830
rect 16859 1270 16893 1830
rect 16893 1270 16902 1830
rect 16968 1270 16977 1830
rect 16977 1270 17011 1830
rect 17011 1270 17020 1830
rect 17086 1270 17095 1830
rect 17095 1270 17129 1830
rect 17129 1270 17138 1830
rect 17204 1270 17213 1830
rect 17213 1270 17247 1830
rect 17247 1270 17256 1830
rect 17322 1270 17331 1830
rect 17331 1270 17365 1830
rect 17365 1270 17374 1830
rect 17440 1270 17449 1830
rect 17449 1270 17483 1830
rect 17483 1270 17492 1830
rect 17558 1270 17567 1830
rect 17567 1270 17601 1830
rect 17601 1270 17610 1830
rect 17676 1270 17685 1830
rect 17685 1270 17719 1830
rect 17719 1270 17728 1830
rect 17794 1270 17803 1830
rect 17803 1270 17837 1830
rect 17837 1270 17846 1830
rect 17912 1270 17921 1830
rect 17921 1270 17955 1830
rect 17955 1270 17964 1830
rect 18030 1270 18039 1830
rect 18039 1270 18073 1830
rect 18073 1270 18082 1830
rect 18148 1270 18157 1830
rect 18157 1270 18191 1830
rect 18191 1270 18200 1830
rect 18266 1270 18275 1830
rect 18275 1270 18309 1830
rect 18309 1270 18318 1830
rect 18384 1270 18393 1830
rect 18393 1270 18427 1830
rect 18427 1270 18436 1830
rect 18502 1270 18511 1830
rect 18511 1270 18545 1830
rect 18545 1270 18554 1830
rect 18620 1270 18629 1830
rect 18629 1270 18663 1830
rect 18663 1270 18672 1830
rect 18738 1270 18747 1830
rect 18747 1270 18781 1830
rect 18781 1270 18790 1830
rect 18856 1270 18865 1830
rect 18865 1270 18899 1830
rect 18899 1270 18908 1830
rect 18974 1270 18983 1830
rect 18983 1270 19017 1830
rect 19017 1270 19026 1830
rect 19092 1270 19101 1830
rect 19101 1270 19135 1830
rect 19135 1270 19144 1830
rect 19210 1270 19219 1830
rect 19219 1270 19253 1830
rect 19253 1270 19262 1830
rect 19328 1270 19337 1830
rect 19337 1270 19371 1830
rect 19371 1270 19380 1830
rect 19446 1270 19455 1830
rect 19455 1270 19489 1830
rect 19489 1270 19498 1830
rect 19564 1270 19573 1830
rect 19573 1270 19607 1830
rect 19607 1270 19616 1830
rect 4801 610 4810 1170
rect 4810 610 4844 1170
rect 4844 610 4853 1170
rect 4917 610 4928 1170
rect 4928 610 4962 1170
rect 4962 610 4969 1170
rect 5037 610 5046 1170
rect 5046 610 5080 1170
rect 5080 610 5089 1170
rect 5153 610 5164 1170
rect 5164 610 5198 1170
rect 5198 610 5205 1170
rect 5273 610 5282 1170
rect 5282 610 5316 1170
rect 5316 610 5325 1170
rect 5389 610 5400 1170
rect 5400 610 5434 1170
rect 5434 610 5441 1170
rect 5509 610 5518 1170
rect 5518 610 5552 1170
rect 5552 610 5561 1170
rect 5625 610 5636 1170
rect 5636 610 5670 1170
rect 5670 610 5677 1170
rect 5745 610 5754 1170
rect 5754 610 5788 1170
rect 5788 610 5797 1170
rect 5861 610 5872 1170
rect 5872 610 5906 1170
rect 5906 610 5913 1170
rect 5981 610 5990 1170
rect 5990 610 6024 1170
rect 6024 610 6033 1170
rect 6097 610 6108 1170
rect 6108 610 6142 1170
rect 6142 610 6149 1170
rect 6217 610 6226 1170
rect 6226 610 6260 1170
rect 6260 610 6269 1170
rect 6333 610 6344 1170
rect 6344 610 6378 1170
rect 6378 610 6385 1170
rect 6453 610 6462 1170
rect 6462 610 6496 1170
rect 6496 610 6505 1170
rect 6569 610 6580 1170
rect 6580 610 6614 1170
rect 6614 610 6621 1170
rect 6689 610 6698 1170
rect 6698 610 6732 1170
rect 6732 610 6741 1170
rect 6805 610 6816 1170
rect 6816 610 6850 1170
rect 6850 610 6857 1170
rect 6925 610 6934 1170
rect 6934 610 6968 1170
rect 6968 610 6977 1170
rect 7041 610 7052 1170
rect 7052 610 7086 1170
rect 7086 610 7093 1170
rect 7161 610 7170 1170
rect 7170 610 7204 1170
rect 7204 610 7213 1170
rect 7277 610 7288 1170
rect 7288 610 7322 1170
rect 7322 610 7329 1170
rect 7397 610 7406 1170
rect 7406 610 7440 1170
rect 7440 610 7449 1170
rect 7513 610 7524 1170
rect 7524 610 7558 1170
rect 7558 610 7565 1170
rect 7633 610 7642 1170
rect 7642 610 7676 1170
rect 7676 610 7685 1170
rect 7749 610 7760 1170
rect 7760 610 7794 1170
rect 7794 610 7801 1170
rect 7869 610 7878 1170
rect 7878 610 7912 1170
rect 7912 610 7921 1170
rect 7985 610 7996 1170
rect 7996 610 8030 1170
rect 8030 610 8037 1170
rect 8105 610 8114 1170
rect 8114 610 8148 1170
rect 8148 610 8157 1170
rect 8221 610 8232 1170
rect 8232 610 8266 1170
rect 8266 610 8273 1170
rect 8341 610 8350 1170
rect 8350 610 8384 1170
rect 8384 610 8393 1170
rect 8457 610 8468 1170
rect 8468 610 8502 1170
rect 8502 610 8509 1170
rect 8577 610 8586 1170
rect 8586 610 8620 1170
rect 8620 610 8629 1170
rect 8693 610 8704 1170
rect 8704 610 8738 1170
rect 8738 610 8745 1170
rect 8813 610 8822 1170
rect 8822 610 8856 1170
rect 8856 610 8865 1170
rect 8929 610 8940 1170
rect 8940 610 8974 1170
rect 8974 610 8981 1170
rect 9049 610 9058 1170
rect 9058 610 9092 1170
rect 9092 610 9101 1170
rect 9165 610 9176 1170
rect 9176 610 9210 1170
rect 9210 610 9217 1170
rect 9285 610 9294 1170
rect 9294 610 9328 1170
rect 9328 610 9337 1170
rect 9401 610 9412 1170
rect 9412 610 9446 1170
rect 9446 610 9453 1170
rect 9521 610 9530 1170
rect 9530 610 9564 1170
rect 9564 610 9573 1170
rect 9637 610 9648 1170
rect 9648 610 9682 1170
rect 9682 610 9689 1170
rect 9757 610 9766 1170
rect 9766 610 9800 1170
rect 9800 610 9809 1170
rect 9873 610 9884 1170
rect 9884 610 9918 1170
rect 9918 610 9925 1170
rect 9993 610 10002 1170
rect 10002 610 10036 1170
rect 10036 610 10045 1170
rect 10109 610 10120 1170
rect 10120 610 10154 1170
rect 10154 610 10161 1170
rect 10229 610 10238 1170
rect 10238 610 10272 1170
rect 10272 610 10281 1170
rect 10345 610 10356 1170
rect 10356 610 10390 1170
rect 10390 610 10397 1170
rect 10465 610 10474 1170
rect 10474 610 10508 1170
rect 10508 610 10517 1170
rect 10581 610 10592 1170
rect 10592 610 10626 1170
rect 10626 610 10633 1170
rect 10701 610 10710 1170
rect 10710 610 10744 1170
rect 10744 610 10753 1170
rect 20737 1270 20746 1830
rect 20746 1270 20780 1830
rect 20780 1270 20789 1830
rect 20855 1270 20864 1830
rect 20864 1270 20898 1830
rect 20898 1270 20907 1830
rect 20973 1270 20982 1830
rect 20982 1270 21016 1830
rect 21016 1270 21025 1830
rect 21091 1270 21100 1830
rect 21100 1270 21134 1830
rect 21134 1270 21143 1830
rect 21209 1270 21218 1830
rect 21218 1270 21252 1830
rect 21252 1270 21261 1830
rect 21327 1270 21336 1830
rect 21336 1270 21370 1830
rect 21370 1270 21379 1830
rect 21445 1270 21454 1830
rect 21454 1270 21488 1830
rect 21488 1270 21497 1830
rect 21563 1270 21572 1830
rect 21572 1270 21606 1830
rect 21606 1270 21615 1830
rect 21681 1270 21690 1830
rect 21690 1270 21724 1830
rect 21724 1270 21733 1830
rect 21799 1270 21808 1830
rect 21808 1270 21842 1830
rect 21842 1270 21851 1830
rect 21917 1270 21926 1830
rect 21926 1270 21960 1830
rect 21960 1270 21969 1830
rect 22035 1270 22044 1830
rect 22044 1270 22078 1830
rect 22078 1270 22087 1830
rect 22153 1270 22162 1830
rect 22162 1270 22196 1830
rect 22196 1270 22205 1830
rect 22271 1270 22280 1830
rect 22280 1270 22314 1830
rect 22314 1270 22323 1830
rect 22389 1270 22398 1830
rect 22398 1270 22432 1830
rect 22432 1270 22441 1830
rect 22507 1270 22516 1830
rect 22516 1270 22550 1830
rect 22550 1270 22559 1830
rect 22625 1270 22634 1830
rect 22634 1270 22668 1830
rect 22668 1270 22677 1830
rect 22743 1270 22752 1830
rect 22752 1270 22786 1830
rect 22786 1270 22795 1830
rect 22861 1270 22870 1830
rect 22870 1270 22904 1830
rect 22904 1270 22913 1830
rect 22979 1270 22988 1830
rect 22988 1270 23022 1830
rect 23022 1270 23031 1830
rect 23097 1270 23106 1830
rect 23106 1270 23140 1830
rect 23140 1270 23149 1830
rect 23215 1270 23224 1830
rect 23224 1270 23258 1830
rect 23258 1270 23267 1830
rect 23333 1270 23342 1830
rect 23342 1270 23376 1830
rect 23376 1270 23385 1830
rect 23451 1270 23460 1830
rect 23460 1270 23494 1830
rect 23494 1270 23503 1830
rect 23569 1270 23578 1830
rect 23578 1270 23612 1830
rect 23612 1270 23621 1830
rect 23687 1270 23696 1830
rect 23696 1270 23730 1830
rect 23730 1270 23739 1830
rect 23895 1839 23905 1853
rect 23905 1839 23939 1853
rect 23939 1839 23947 1853
rect 23895 1801 23947 1839
rect 23975 1839 23977 1853
rect 23977 1839 24011 1853
rect 24011 1839 24027 1853
rect 24055 1839 24083 1853
rect 24083 1839 24107 1853
rect 24135 1839 24155 1853
rect 24155 1839 24187 1853
rect 24215 1839 24227 1853
rect 24227 1839 24265 1853
rect 24265 1839 24267 1853
rect 24295 1839 24299 1853
rect 24299 1839 24337 1853
rect 24337 1839 24347 1853
rect 24375 1839 24409 1853
rect 24409 1839 24427 1853
rect 24455 1839 24481 1853
rect 24481 1839 24507 1853
rect 24535 1839 24553 1853
rect 24553 1839 24587 1853
rect 23975 1801 24027 1839
rect 24055 1801 24107 1839
rect 24135 1801 24187 1839
rect 24215 1801 24267 1839
rect 24295 1801 24347 1839
rect 24375 1801 24427 1839
rect 24455 1801 24507 1839
rect 24535 1801 24587 1839
rect 24615 1839 24625 1853
rect 24625 1839 24659 1853
rect 24659 1839 24667 1853
rect 24615 1801 24667 1839
rect 24695 1801 24747 1853
rect 24775 1801 24827 1853
rect 24855 1801 24907 1853
rect 24935 1801 24987 1853
rect 25015 1801 25067 1853
rect 23895 1765 23905 1773
rect 23905 1765 23939 1773
rect 23939 1765 23947 1773
rect 23895 1725 23947 1765
rect 23895 1721 23905 1725
rect 23905 1721 23939 1725
rect 23939 1721 23947 1725
rect 23975 1765 23977 1773
rect 23977 1765 24011 1773
rect 24011 1765 24027 1773
rect 24055 1765 24083 1773
rect 24083 1765 24107 1773
rect 24135 1765 24155 1773
rect 24155 1765 24187 1773
rect 24215 1765 24227 1773
rect 24227 1765 24265 1773
rect 24265 1765 24267 1773
rect 24295 1765 24299 1773
rect 24299 1765 24337 1773
rect 24337 1765 24347 1773
rect 24375 1765 24409 1773
rect 24409 1765 24427 1773
rect 24455 1765 24481 1773
rect 24481 1765 24507 1773
rect 24535 1765 24553 1773
rect 24553 1765 24587 1773
rect 23975 1725 24027 1765
rect 24055 1725 24107 1765
rect 24135 1725 24187 1765
rect 24215 1725 24267 1765
rect 24295 1725 24347 1765
rect 24375 1725 24427 1765
rect 24455 1725 24507 1765
rect 24535 1725 24587 1765
rect 23975 1721 23977 1725
rect 23977 1721 24011 1725
rect 24011 1721 24027 1725
rect 24055 1721 24083 1725
rect 24083 1721 24107 1725
rect 24135 1721 24155 1725
rect 24155 1721 24187 1725
rect 24215 1721 24227 1725
rect 24227 1721 24265 1725
rect 24265 1721 24267 1725
rect 24295 1721 24299 1725
rect 24299 1721 24337 1725
rect 24337 1721 24347 1725
rect 24375 1721 24409 1725
rect 24409 1721 24427 1725
rect 24455 1721 24481 1725
rect 24481 1721 24507 1725
rect 24535 1721 24553 1725
rect 24553 1721 24587 1725
rect 24615 1765 24625 1773
rect 24625 1765 24659 1773
rect 24659 1765 24667 1773
rect 24615 1725 24667 1765
rect 24615 1721 24625 1725
rect 24625 1721 24659 1725
rect 24659 1721 24667 1725
rect 24695 1721 24747 1773
rect 24775 1721 24827 1773
rect 24855 1721 24907 1773
rect 24935 1721 24987 1773
rect 25015 1721 25067 1773
rect 23895 1691 23905 1693
rect 23905 1691 23939 1693
rect 23939 1691 23947 1693
rect 23895 1651 23947 1691
rect 23895 1641 23905 1651
rect 23905 1641 23939 1651
rect 23939 1641 23947 1651
rect 23975 1691 23977 1693
rect 23977 1691 24011 1693
rect 24011 1691 24027 1693
rect 24055 1691 24083 1693
rect 24083 1691 24107 1693
rect 24135 1691 24155 1693
rect 24155 1691 24187 1693
rect 24215 1691 24227 1693
rect 24227 1691 24265 1693
rect 24265 1691 24267 1693
rect 24295 1691 24299 1693
rect 24299 1691 24337 1693
rect 24337 1691 24347 1693
rect 24375 1691 24409 1693
rect 24409 1691 24427 1693
rect 24455 1691 24481 1693
rect 24481 1691 24507 1693
rect 24535 1691 24553 1693
rect 24553 1691 24587 1693
rect 23975 1651 24027 1691
rect 24055 1651 24107 1691
rect 24135 1651 24187 1691
rect 24215 1651 24267 1691
rect 24295 1651 24347 1691
rect 24375 1651 24427 1691
rect 24455 1651 24507 1691
rect 24535 1651 24587 1691
rect 23975 1641 23977 1651
rect 23977 1641 24011 1651
rect 24011 1641 24027 1651
rect 24055 1641 24083 1651
rect 24083 1641 24107 1651
rect 24135 1641 24155 1651
rect 24155 1641 24187 1651
rect 24215 1641 24227 1651
rect 24227 1641 24265 1651
rect 24265 1641 24267 1651
rect 24295 1641 24299 1651
rect 24299 1641 24337 1651
rect 24337 1641 24347 1651
rect 24375 1641 24409 1651
rect 24409 1641 24427 1651
rect 24455 1641 24481 1651
rect 24481 1641 24507 1651
rect 24535 1641 24553 1651
rect 24553 1641 24587 1651
rect 24615 1691 24625 1693
rect 24625 1691 24659 1693
rect 24659 1691 24667 1693
rect 24615 1651 24667 1691
rect 24615 1641 24625 1651
rect 24625 1641 24659 1651
rect 24659 1641 24667 1651
rect 24695 1641 24747 1693
rect 24775 1641 24827 1693
rect 24855 1641 24907 1693
rect 24935 1641 24987 1693
rect 25015 1641 25067 1693
rect 23895 1577 23947 1613
rect 23895 1561 23905 1577
rect 23905 1561 23939 1577
rect 23939 1561 23947 1577
rect 23975 1577 24027 1613
rect 24055 1577 24107 1613
rect 24135 1577 24187 1613
rect 24215 1577 24267 1613
rect 24295 1577 24347 1613
rect 24375 1577 24427 1613
rect 24455 1577 24507 1613
rect 24535 1577 24587 1613
rect 23975 1561 23977 1577
rect 23977 1561 24011 1577
rect 24011 1561 24027 1577
rect 24055 1561 24083 1577
rect 24083 1561 24107 1577
rect 24135 1561 24155 1577
rect 24155 1561 24187 1577
rect 24215 1561 24227 1577
rect 24227 1561 24265 1577
rect 24265 1561 24267 1577
rect 24295 1561 24299 1577
rect 24299 1561 24337 1577
rect 24337 1561 24347 1577
rect 24375 1561 24409 1577
rect 24409 1561 24427 1577
rect 24455 1561 24481 1577
rect 24481 1561 24507 1577
rect 24535 1561 24553 1577
rect 24553 1561 24587 1577
rect 24615 1577 24667 1613
rect 24615 1561 24625 1577
rect 24625 1561 24659 1577
rect 24659 1561 24667 1577
rect 24695 1561 24747 1613
rect 24775 1561 24827 1613
rect 24855 1561 24907 1613
rect 24935 1561 24987 1613
rect 25015 1561 25067 1613
rect 23895 1503 23947 1533
rect 23895 1481 23905 1503
rect 23905 1481 23939 1503
rect 23939 1481 23947 1503
rect 23975 1503 24027 1533
rect 24055 1503 24107 1533
rect 24135 1503 24187 1533
rect 24215 1503 24267 1533
rect 24295 1503 24347 1533
rect 24375 1503 24427 1533
rect 24455 1503 24507 1533
rect 24535 1503 24587 1533
rect 23975 1481 23977 1503
rect 23977 1481 24011 1503
rect 24011 1481 24027 1503
rect 24055 1481 24083 1503
rect 24083 1481 24107 1503
rect 24135 1481 24155 1503
rect 24155 1481 24187 1503
rect 24215 1481 24227 1503
rect 24227 1481 24265 1503
rect 24265 1481 24267 1503
rect 24295 1481 24299 1503
rect 24299 1481 24337 1503
rect 24337 1481 24347 1503
rect 24375 1481 24409 1503
rect 24409 1481 24427 1503
rect 24455 1481 24481 1503
rect 24481 1481 24507 1503
rect 24535 1481 24553 1503
rect 24553 1481 24587 1503
rect 24615 1503 24667 1533
rect 24615 1481 24625 1503
rect 24625 1481 24659 1503
rect 24659 1481 24667 1503
rect 24695 1481 24747 1533
rect 24775 1481 24827 1533
rect 24855 1481 24907 1533
rect 24935 1481 24987 1533
rect 25015 1481 25067 1533
rect 23895 1429 23947 1453
rect 23895 1401 23905 1429
rect 23905 1401 23939 1429
rect 23939 1401 23947 1429
rect 23975 1429 24027 1453
rect 24055 1429 24107 1453
rect 24135 1429 24187 1453
rect 24215 1429 24267 1453
rect 24295 1429 24347 1453
rect 24375 1429 24427 1453
rect 24455 1429 24507 1453
rect 24535 1429 24587 1453
rect 23975 1401 23977 1429
rect 23977 1401 24011 1429
rect 24011 1401 24027 1429
rect 24055 1401 24083 1429
rect 24083 1401 24107 1429
rect 24135 1401 24155 1429
rect 24155 1401 24187 1429
rect 24215 1401 24227 1429
rect 24227 1401 24265 1429
rect 24265 1401 24267 1429
rect 24295 1401 24299 1429
rect 24299 1401 24337 1429
rect 24337 1401 24347 1429
rect 24375 1401 24409 1429
rect 24409 1401 24427 1429
rect 24455 1401 24481 1429
rect 24481 1401 24507 1429
rect 24535 1401 24553 1429
rect 24553 1401 24587 1429
rect 24615 1429 24667 1453
rect 24615 1401 24625 1429
rect 24625 1401 24659 1429
rect 24659 1401 24667 1429
rect 24695 1401 24747 1453
rect 24775 1401 24827 1453
rect 24855 1401 24907 1453
rect 24935 1401 24987 1453
rect 25015 1401 25067 1453
rect 23895 1355 23947 1373
rect 23895 1321 23905 1355
rect 23905 1321 23939 1355
rect 23939 1321 23947 1355
rect 23975 1355 24027 1373
rect 24055 1355 24107 1373
rect 24135 1355 24187 1373
rect 24215 1355 24267 1373
rect 24295 1355 24347 1373
rect 24375 1355 24427 1373
rect 24455 1355 24507 1373
rect 24535 1355 24587 1373
rect 23975 1321 23977 1355
rect 23977 1321 24011 1355
rect 24011 1321 24027 1355
rect 24055 1321 24083 1355
rect 24083 1321 24107 1355
rect 24135 1321 24155 1355
rect 24155 1321 24187 1355
rect 24215 1321 24227 1355
rect 24227 1321 24265 1355
rect 24265 1321 24267 1355
rect 24295 1321 24299 1355
rect 24299 1321 24337 1355
rect 24337 1321 24347 1355
rect 24375 1321 24409 1355
rect 24409 1321 24427 1355
rect 24455 1321 24481 1355
rect 24481 1321 24507 1355
rect 24535 1321 24553 1355
rect 24553 1321 24587 1355
rect 24615 1355 24667 1373
rect 24615 1321 24625 1355
rect 24625 1321 24659 1355
rect 24659 1321 24667 1355
rect 24695 1321 24747 1373
rect 24775 1321 24827 1373
rect 24855 1321 24907 1373
rect 24935 1321 24987 1373
rect 25015 1321 25067 1373
rect 23895 1281 23947 1293
rect 23895 1247 23905 1281
rect 23905 1247 23939 1281
rect 23939 1247 23947 1281
rect 23895 1241 23947 1247
rect 23975 1281 24027 1293
rect 24055 1281 24107 1293
rect 24135 1281 24187 1293
rect 24215 1281 24267 1293
rect 24295 1281 24347 1293
rect 24375 1281 24427 1293
rect 24455 1281 24507 1293
rect 24535 1281 24587 1293
rect 23975 1247 23977 1281
rect 23977 1247 24011 1281
rect 24011 1247 24027 1281
rect 24055 1247 24083 1281
rect 24083 1247 24107 1281
rect 24135 1247 24155 1281
rect 24155 1247 24187 1281
rect 24215 1247 24227 1281
rect 24227 1247 24265 1281
rect 24265 1247 24267 1281
rect 24295 1247 24299 1281
rect 24299 1247 24337 1281
rect 24337 1247 24347 1281
rect 24375 1247 24409 1281
rect 24409 1247 24427 1281
rect 24455 1247 24481 1281
rect 24481 1247 24507 1281
rect 24535 1247 24553 1281
rect 24553 1247 24587 1281
rect 23975 1241 24027 1247
rect 24055 1241 24107 1247
rect 24135 1241 24187 1247
rect 24215 1241 24267 1247
rect 24295 1241 24347 1247
rect 24375 1241 24427 1247
rect 24455 1241 24507 1247
rect 24535 1241 24587 1247
rect 24615 1281 24667 1293
rect 24615 1247 24625 1281
rect 24625 1247 24659 1281
rect 24659 1247 24667 1281
rect 24615 1241 24667 1247
rect 24695 1241 24747 1293
rect 24775 1241 24827 1293
rect 24855 1241 24907 1293
rect 24935 1241 24987 1293
rect 25015 1241 25067 1293
rect 12485 1101 12537 1149
rect 12485 1097 12513 1101
rect 12513 1097 12537 1101
rect 12565 1097 12617 1149
rect 12645 1097 12697 1149
rect 12725 1097 12777 1149
rect 12805 1097 12857 1149
rect 12885 1097 12937 1149
rect 12965 1097 13017 1149
rect 13045 1097 13097 1149
rect 13125 1097 13177 1149
rect 13205 1097 13257 1149
rect 13285 1097 13337 1149
rect 13365 1097 13417 1149
rect 13445 1097 13497 1149
rect 13525 1097 13577 1149
rect 13605 1097 13657 1149
rect 13685 1097 13737 1149
rect 13765 1097 13817 1149
rect 13845 1097 13897 1149
rect 13925 1097 13977 1149
rect 14005 1097 14057 1149
rect 14085 1097 14137 1149
rect 14165 1097 14217 1149
rect 14245 1097 14297 1149
rect 14325 1097 14377 1149
rect 14405 1097 14457 1149
rect 14485 1097 14537 1149
rect 14565 1097 14617 1149
rect 14645 1097 14697 1149
rect 14725 1097 14777 1149
rect 14805 1097 14857 1149
rect 14885 1097 14937 1149
rect 14965 1097 15017 1149
rect 15045 1097 15097 1149
rect 15125 1097 15177 1149
rect 15205 1097 15257 1149
rect 15285 1097 15337 1149
rect 15365 1097 15417 1149
rect 15445 1097 15497 1149
rect 15525 1097 15577 1149
rect 15605 1097 15657 1149
rect 15685 1097 15737 1149
rect 15765 1097 15817 1149
rect 15845 1097 15897 1149
rect 15925 1097 15977 1149
rect 16005 1097 16057 1149
rect 16085 1097 16137 1149
rect 16165 1097 16217 1149
rect 16245 1097 16297 1149
rect 16325 1097 16377 1149
rect 16405 1097 16457 1149
rect 16485 1097 16537 1149
rect 16565 1097 16617 1149
rect 16645 1097 16697 1149
rect 16725 1097 16777 1149
rect 16805 1097 16857 1149
rect 16885 1097 16937 1149
rect 16965 1097 17017 1149
rect 17045 1097 17097 1149
rect 17125 1097 17177 1149
rect 17205 1097 17257 1149
rect 17285 1097 17337 1149
rect 17365 1097 17417 1149
rect 17445 1097 17497 1149
rect 17525 1097 17577 1149
rect 17605 1097 17657 1149
rect 17685 1097 17737 1149
rect 17765 1097 17817 1149
rect 17845 1097 17897 1149
rect 17925 1097 17977 1149
rect 18005 1097 18057 1149
rect 18085 1097 18137 1149
rect 18165 1097 18217 1149
rect 18245 1097 18297 1149
rect 18325 1097 18377 1149
rect 18405 1097 18457 1149
rect 18485 1097 18537 1149
rect 18565 1097 18617 1149
rect 18645 1097 18697 1149
rect 18725 1097 18777 1149
rect 18805 1097 18857 1149
rect 18885 1097 18937 1149
rect 18965 1097 19017 1149
rect 19045 1097 19097 1149
rect 19125 1097 19177 1149
rect 19205 1097 19257 1149
rect 19285 1097 19337 1149
rect 19365 1097 19417 1149
rect 19445 1097 19497 1149
rect 19525 1097 19577 1149
rect 19605 1097 19657 1149
rect 19685 1097 19737 1149
rect 19765 1097 19817 1149
rect 19845 1097 19897 1149
rect 19925 1097 19977 1149
rect 20005 1097 20057 1149
rect 20085 1097 20137 1149
rect 20165 1097 20217 1149
rect 20245 1097 20297 1149
rect 20325 1097 20377 1149
rect 20405 1097 20457 1149
rect 20485 1097 20537 1149
rect 20565 1097 20617 1149
rect 20645 1097 20697 1149
rect 20725 1097 20777 1149
rect 20805 1097 20857 1149
rect 20885 1097 20937 1149
rect 20965 1097 21017 1149
rect 21045 1097 21097 1149
rect 21125 1097 21177 1149
rect 21205 1097 21257 1149
rect 21285 1097 21337 1149
rect 21365 1097 21417 1149
rect 21445 1097 21497 1149
rect 21525 1097 21577 1149
rect 21605 1097 21657 1149
rect 21685 1097 21737 1149
rect 21765 1097 21817 1149
rect 21845 1097 21897 1149
rect 21925 1097 21977 1149
rect 22005 1097 22057 1149
rect 22085 1097 22137 1149
rect 22165 1097 22217 1149
rect 22245 1097 22297 1149
rect 22325 1097 22377 1149
rect 22405 1097 22457 1149
rect 22485 1097 22537 1149
rect 22565 1097 22617 1149
rect 22645 1097 22697 1149
rect 22725 1097 22777 1149
rect 22805 1097 22857 1149
rect 22885 1097 22937 1149
rect 22965 1097 23017 1149
rect 23045 1097 23097 1149
rect 23125 1097 23177 1149
rect 23205 1097 23257 1149
rect 23285 1097 23337 1149
rect 23365 1097 23417 1149
rect 23445 1097 23497 1149
rect 23525 1097 23577 1149
rect 23605 1097 23657 1149
rect 23685 1097 23737 1149
rect 23765 1097 23817 1149
rect 23845 1097 23897 1149
rect 23925 1097 23977 1149
rect 24005 1097 24057 1149
rect 24085 1097 24137 1149
rect 24165 1097 24217 1149
rect 24245 1097 24297 1149
rect 24325 1097 24377 1149
rect 24405 1097 24457 1149
rect 12485 1067 12513 1069
rect 12513 1067 12537 1069
rect 12485 1017 12537 1067
rect 12565 1017 12617 1069
rect 12645 1017 12697 1069
rect 12725 1017 12777 1069
rect 12805 1017 12857 1069
rect 12885 1017 12937 1069
rect 12965 1017 13017 1069
rect 13045 1017 13097 1069
rect 13125 1017 13177 1069
rect 13205 1017 13257 1069
rect 13285 1017 13337 1069
rect 13365 1017 13417 1069
rect 13445 1017 13497 1069
rect 13525 1017 13577 1069
rect 13605 1017 13657 1069
rect 13685 1017 13737 1069
rect 13765 1017 13817 1069
rect 13845 1017 13897 1069
rect 13925 1017 13977 1069
rect 14005 1017 14057 1069
rect 14085 1017 14137 1069
rect 14165 1017 14217 1069
rect 14245 1017 14297 1069
rect 14325 1017 14377 1069
rect 14405 1017 14457 1069
rect 14485 1017 14537 1069
rect 14565 1017 14617 1069
rect 14645 1017 14697 1069
rect 14725 1017 14777 1069
rect 14805 1017 14857 1069
rect 14885 1017 14937 1069
rect 14965 1017 15017 1069
rect 15045 1017 15097 1069
rect 15125 1017 15177 1069
rect 15205 1017 15257 1069
rect 15285 1017 15337 1069
rect 15365 1017 15417 1069
rect 15445 1017 15497 1069
rect 15525 1017 15577 1069
rect 15605 1017 15657 1069
rect 15685 1017 15737 1069
rect 15765 1017 15817 1069
rect 15845 1017 15897 1069
rect 15925 1017 15977 1069
rect 16005 1017 16057 1069
rect 16085 1017 16137 1069
rect 16165 1017 16217 1069
rect 16245 1017 16297 1069
rect 16325 1017 16377 1069
rect 16405 1017 16457 1069
rect 16485 1017 16537 1069
rect 16565 1017 16617 1069
rect 16645 1017 16697 1069
rect 16725 1017 16777 1069
rect 16805 1017 16857 1069
rect 16885 1017 16937 1069
rect 16965 1017 17017 1069
rect 17045 1017 17097 1069
rect 17125 1017 17177 1069
rect 17205 1017 17257 1069
rect 17285 1017 17337 1069
rect 17365 1017 17417 1069
rect 17445 1017 17497 1069
rect 17525 1017 17577 1069
rect 17605 1017 17657 1069
rect 17685 1017 17737 1069
rect 17765 1017 17817 1069
rect 17845 1017 17897 1069
rect 17925 1017 17977 1069
rect 18005 1017 18057 1069
rect 18085 1017 18137 1069
rect 18165 1017 18217 1069
rect 18245 1017 18297 1069
rect 18325 1017 18377 1069
rect 18405 1017 18457 1069
rect 18485 1017 18537 1069
rect 18565 1017 18617 1069
rect 18645 1017 18697 1069
rect 18725 1017 18777 1069
rect 18805 1017 18857 1069
rect 18885 1017 18937 1069
rect 18965 1017 19017 1069
rect 19045 1017 19097 1069
rect 19125 1017 19177 1069
rect 19205 1017 19257 1069
rect 19285 1017 19337 1069
rect 19365 1017 19417 1069
rect 19445 1017 19497 1069
rect 19525 1017 19577 1069
rect 19605 1017 19657 1069
rect 19685 1017 19737 1069
rect 19765 1017 19817 1069
rect 19845 1017 19897 1069
rect 19925 1017 19977 1069
rect 20005 1017 20057 1069
rect 20085 1017 20137 1069
rect 20165 1017 20217 1069
rect 20245 1017 20297 1069
rect 20325 1017 20377 1069
rect 20405 1017 20457 1069
rect 20485 1017 20537 1069
rect 20565 1017 20617 1069
rect 20645 1017 20697 1069
rect 20725 1017 20777 1069
rect 20805 1017 20857 1069
rect 20885 1017 20937 1069
rect 20965 1017 21017 1069
rect 21045 1017 21097 1069
rect 21125 1017 21177 1069
rect 21205 1017 21257 1069
rect 21285 1017 21337 1069
rect 21365 1017 21417 1069
rect 21445 1017 21497 1069
rect 21525 1017 21577 1069
rect 21605 1017 21657 1069
rect 21685 1017 21737 1069
rect 21765 1017 21817 1069
rect 21845 1017 21897 1069
rect 21925 1017 21977 1069
rect 22005 1017 22057 1069
rect 22085 1017 22137 1069
rect 22165 1017 22217 1069
rect 22245 1017 22297 1069
rect 22325 1017 22377 1069
rect 22405 1017 22457 1069
rect 22485 1017 22537 1069
rect 22565 1017 22617 1069
rect 22645 1017 22697 1069
rect 22725 1017 22777 1069
rect 22805 1017 22857 1069
rect 22885 1017 22937 1069
rect 22965 1017 23017 1069
rect 23045 1017 23097 1069
rect 23125 1017 23177 1069
rect 23205 1017 23257 1069
rect 23285 1017 23337 1069
rect 23365 1017 23417 1069
rect 23445 1017 23497 1069
rect 23525 1017 23577 1069
rect 23605 1017 23657 1069
rect 23685 1017 23737 1069
rect 23765 1017 23817 1069
rect 23845 1017 23897 1069
rect 23925 1017 23977 1069
rect 24005 1017 24057 1069
rect 24085 1017 24137 1069
rect 24165 1017 24217 1069
rect 24245 1017 24297 1069
rect 24325 1017 24377 1069
rect 24405 1017 24457 1069
rect 4857 543 4915 549
rect 4857 509 4869 543
rect 4869 509 4903 543
rect 4903 509 4915 543
rect 4857 435 4915 509
rect 4857 401 4869 435
rect 4869 401 4903 435
rect 4903 401 4915 435
rect 4857 395 4915 401
rect 4975 543 5033 549
rect 4975 509 4987 543
rect 4987 509 5021 543
rect 5021 509 5033 543
rect 4975 435 5033 509
rect 4975 401 4987 435
rect 4987 401 5021 435
rect 5021 401 5033 435
rect 4975 395 5033 401
rect 5093 543 5151 549
rect 5093 509 5105 543
rect 5105 509 5139 543
rect 5139 509 5151 543
rect 5093 435 5151 509
rect 5093 401 5105 435
rect 5105 401 5139 435
rect 5139 401 5151 435
rect 5093 395 5151 401
rect 5211 543 5269 549
rect 5211 509 5223 543
rect 5223 509 5257 543
rect 5257 509 5269 543
rect 5211 435 5269 509
rect 5211 401 5223 435
rect 5223 401 5257 435
rect 5257 401 5269 435
rect 5211 395 5269 401
rect 5329 543 5387 549
rect 5329 509 5341 543
rect 5341 509 5375 543
rect 5375 509 5387 543
rect 5329 435 5387 509
rect 5329 401 5341 435
rect 5341 401 5375 435
rect 5375 401 5387 435
rect 5329 395 5387 401
rect 5447 543 5505 549
rect 5447 509 5459 543
rect 5459 509 5493 543
rect 5493 509 5505 543
rect 5447 435 5505 509
rect 5447 401 5459 435
rect 5459 401 5493 435
rect 5493 401 5505 435
rect 5447 395 5505 401
rect 5565 543 5623 549
rect 5565 509 5577 543
rect 5577 509 5611 543
rect 5611 509 5623 543
rect 5565 435 5623 509
rect 5565 401 5577 435
rect 5577 401 5611 435
rect 5611 401 5623 435
rect 5565 395 5623 401
rect 5683 543 5741 549
rect 5683 509 5695 543
rect 5695 509 5729 543
rect 5729 509 5741 543
rect 5683 435 5741 509
rect 5683 401 5695 435
rect 5695 401 5729 435
rect 5729 401 5741 435
rect 5683 395 5741 401
rect 5801 543 5859 549
rect 5801 509 5813 543
rect 5813 509 5847 543
rect 5847 509 5859 543
rect 5801 435 5859 509
rect 5801 401 5813 435
rect 5813 401 5847 435
rect 5847 401 5859 435
rect 5801 395 5859 401
rect 5919 543 5977 549
rect 5919 509 5931 543
rect 5931 509 5965 543
rect 5965 509 5977 543
rect 5919 435 5977 509
rect 5919 401 5931 435
rect 5931 401 5965 435
rect 5965 401 5977 435
rect 5919 395 5977 401
rect 6037 543 6095 549
rect 6037 509 6049 543
rect 6049 509 6083 543
rect 6083 509 6095 543
rect 6037 435 6095 509
rect 6037 401 6049 435
rect 6049 401 6083 435
rect 6083 401 6095 435
rect 6037 395 6095 401
rect 6155 543 6213 549
rect 6155 509 6167 543
rect 6167 509 6201 543
rect 6201 509 6213 543
rect 6155 435 6213 509
rect 6155 401 6167 435
rect 6167 401 6201 435
rect 6201 401 6213 435
rect 6155 395 6213 401
rect 6273 543 6331 549
rect 6273 509 6285 543
rect 6285 509 6319 543
rect 6319 509 6331 543
rect 6273 435 6331 509
rect 6273 401 6285 435
rect 6285 401 6319 435
rect 6319 401 6331 435
rect 6273 395 6331 401
rect 6391 543 6449 549
rect 6391 509 6403 543
rect 6403 509 6437 543
rect 6437 509 6449 543
rect 6391 435 6449 509
rect 6391 401 6403 435
rect 6403 401 6437 435
rect 6437 401 6449 435
rect 6391 395 6449 401
rect 6509 543 6567 549
rect 6509 509 6521 543
rect 6521 509 6555 543
rect 6555 509 6567 543
rect 6509 435 6567 509
rect 6509 401 6521 435
rect 6521 401 6555 435
rect 6555 401 6567 435
rect 6509 395 6567 401
rect 6627 543 6685 549
rect 6627 509 6639 543
rect 6639 509 6673 543
rect 6673 509 6685 543
rect 6627 435 6685 509
rect 6627 401 6639 435
rect 6639 401 6673 435
rect 6673 401 6685 435
rect 6627 395 6685 401
rect 6745 543 6803 549
rect 6745 509 6757 543
rect 6757 509 6791 543
rect 6791 509 6803 543
rect 6745 435 6803 509
rect 6745 401 6757 435
rect 6757 401 6791 435
rect 6791 401 6803 435
rect 6745 395 6803 401
rect 6863 543 6921 549
rect 6863 509 6875 543
rect 6875 509 6909 543
rect 6909 509 6921 543
rect 6863 435 6921 509
rect 6863 401 6875 435
rect 6875 401 6909 435
rect 6909 401 6921 435
rect 6863 395 6921 401
rect 6981 543 7039 549
rect 6981 509 6993 543
rect 6993 509 7027 543
rect 7027 509 7039 543
rect 6981 435 7039 509
rect 6981 401 6993 435
rect 6993 401 7027 435
rect 7027 401 7039 435
rect 6981 395 7039 401
rect 7099 543 7157 549
rect 7099 509 7111 543
rect 7111 509 7145 543
rect 7145 509 7157 543
rect 7099 435 7157 509
rect 7099 401 7111 435
rect 7111 401 7145 435
rect 7145 401 7157 435
rect 7099 395 7157 401
rect 7217 543 7275 549
rect 7217 509 7229 543
rect 7229 509 7263 543
rect 7263 509 7275 543
rect 7217 435 7275 509
rect 7217 401 7229 435
rect 7229 401 7263 435
rect 7263 401 7275 435
rect 7217 395 7275 401
rect 7335 543 7393 549
rect 7335 509 7347 543
rect 7347 509 7381 543
rect 7381 509 7393 543
rect 7335 435 7393 509
rect 7335 401 7347 435
rect 7347 401 7381 435
rect 7381 401 7393 435
rect 7335 395 7393 401
rect 7453 543 7511 549
rect 7453 509 7465 543
rect 7465 509 7499 543
rect 7499 509 7511 543
rect 7453 435 7511 509
rect 7453 401 7465 435
rect 7465 401 7499 435
rect 7499 401 7511 435
rect 7453 395 7511 401
rect 7571 543 7629 549
rect 7571 509 7583 543
rect 7583 509 7617 543
rect 7617 509 7629 543
rect 7571 435 7629 509
rect 7571 401 7583 435
rect 7583 401 7617 435
rect 7617 401 7629 435
rect 7571 395 7629 401
rect 7689 543 7747 549
rect 7689 509 7701 543
rect 7701 509 7735 543
rect 7735 509 7747 543
rect 7689 435 7747 509
rect 7689 401 7701 435
rect 7701 401 7735 435
rect 7735 401 7747 435
rect 7689 395 7747 401
rect 7807 543 7865 549
rect 7807 509 7819 543
rect 7819 509 7853 543
rect 7853 509 7865 543
rect 7807 435 7865 509
rect 7807 401 7819 435
rect 7819 401 7853 435
rect 7853 401 7865 435
rect 7807 395 7865 401
rect 7925 543 7983 549
rect 7925 509 7937 543
rect 7937 509 7971 543
rect 7971 509 7983 543
rect 7925 435 7983 509
rect 7925 401 7937 435
rect 7937 401 7971 435
rect 7971 401 7983 435
rect 7925 395 7983 401
rect 8043 543 8101 549
rect 8043 509 8055 543
rect 8055 509 8089 543
rect 8089 509 8101 543
rect 8043 435 8101 509
rect 8043 401 8055 435
rect 8055 401 8089 435
rect 8089 401 8101 435
rect 8043 395 8101 401
rect 8161 543 8219 549
rect 8161 509 8173 543
rect 8173 509 8207 543
rect 8207 509 8219 543
rect 8161 435 8219 509
rect 8161 401 8173 435
rect 8173 401 8207 435
rect 8207 401 8219 435
rect 8161 395 8219 401
rect 8279 543 8337 549
rect 8279 509 8291 543
rect 8291 509 8325 543
rect 8325 509 8337 543
rect 8279 435 8337 509
rect 8279 401 8291 435
rect 8291 401 8325 435
rect 8325 401 8337 435
rect 8279 395 8337 401
rect 8397 543 8455 549
rect 8397 509 8409 543
rect 8409 509 8443 543
rect 8443 509 8455 543
rect 8397 435 8455 509
rect 8397 401 8409 435
rect 8409 401 8443 435
rect 8443 401 8455 435
rect 8397 395 8455 401
rect 8515 543 8573 549
rect 8515 509 8527 543
rect 8527 509 8561 543
rect 8561 509 8573 543
rect 8515 435 8573 509
rect 8515 401 8527 435
rect 8527 401 8561 435
rect 8561 401 8573 435
rect 8515 395 8573 401
rect 8633 543 8691 549
rect 8633 509 8645 543
rect 8645 509 8679 543
rect 8679 509 8691 543
rect 8633 435 8691 509
rect 8633 401 8645 435
rect 8645 401 8679 435
rect 8679 401 8691 435
rect 8633 395 8691 401
rect 8751 543 8809 549
rect 8751 509 8763 543
rect 8763 509 8797 543
rect 8797 509 8809 543
rect 8751 435 8809 509
rect 8751 401 8763 435
rect 8763 401 8797 435
rect 8797 401 8809 435
rect 8751 395 8809 401
rect 8869 543 8927 549
rect 8869 509 8881 543
rect 8881 509 8915 543
rect 8915 509 8927 543
rect 8869 435 8927 509
rect 8869 401 8881 435
rect 8881 401 8915 435
rect 8915 401 8927 435
rect 8869 395 8927 401
rect 8987 543 9045 549
rect 8987 509 8999 543
rect 8999 509 9033 543
rect 9033 509 9045 543
rect 8987 435 9045 509
rect 8987 401 8999 435
rect 8999 401 9033 435
rect 9033 401 9045 435
rect 8987 395 9045 401
rect 9105 543 9163 549
rect 9105 509 9117 543
rect 9117 509 9151 543
rect 9151 509 9163 543
rect 9105 435 9163 509
rect 9105 401 9117 435
rect 9117 401 9151 435
rect 9151 401 9163 435
rect 9105 395 9163 401
rect 9223 543 9281 549
rect 9223 509 9235 543
rect 9235 509 9269 543
rect 9269 509 9281 543
rect 9223 435 9281 509
rect 9223 401 9235 435
rect 9235 401 9269 435
rect 9269 401 9281 435
rect 9223 395 9281 401
rect 9341 543 9399 549
rect 9341 509 9353 543
rect 9353 509 9387 543
rect 9387 509 9399 543
rect 9341 435 9399 509
rect 9341 401 9353 435
rect 9353 401 9387 435
rect 9387 401 9399 435
rect 9341 395 9399 401
rect 9459 543 9517 549
rect 9459 509 9471 543
rect 9471 509 9505 543
rect 9505 509 9517 543
rect 9459 435 9517 509
rect 9459 401 9471 435
rect 9471 401 9505 435
rect 9505 401 9517 435
rect 9459 395 9517 401
rect 9577 543 9635 549
rect 9577 509 9589 543
rect 9589 509 9623 543
rect 9623 509 9635 543
rect 9577 435 9635 509
rect 9577 401 9589 435
rect 9589 401 9623 435
rect 9623 401 9635 435
rect 9577 395 9635 401
rect 9695 543 9753 549
rect 9695 509 9707 543
rect 9707 509 9741 543
rect 9741 509 9753 543
rect 9695 435 9753 509
rect 9695 401 9707 435
rect 9707 401 9741 435
rect 9741 401 9753 435
rect 9695 395 9753 401
rect 9813 543 9871 549
rect 9813 509 9825 543
rect 9825 509 9859 543
rect 9859 509 9871 543
rect 9813 435 9871 509
rect 9813 401 9825 435
rect 9825 401 9859 435
rect 9859 401 9871 435
rect 9813 395 9871 401
rect 9931 543 9989 549
rect 9931 509 9943 543
rect 9943 509 9977 543
rect 9977 509 9989 543
rect 9931 435 9989 509
rect 9931 401 9943 435
rect 9943 401 9977 435
rect 9977 401 9989 435
rect 9931 395 9989 401
rect 10049 543 10107 549
rect 10049 509 10061 543
rect 10061 509 10095 543
rect 10095 509 10107 543
rect 10049 435 10107 509
rect 10049 401 10061 435
rect 10061 401 10095 435
rect 10095 401 10107 435
rect 10049 395 10107 401
rect 10167 543 10225 549
rect 10167 509 10179 543
rect 10179 509 10213 543
rect 10213 509 10225 543
rect 10167 435 10225 509
rect 10167 401 10179 435
rect 10179 401 10213 435
rect 10213 401 10225 435
rect 10167 395 10225 401
rect 10285 543 10343 549
rect 10285 509 10297 543
rect 10297 509 10331 543
rect 10331 509 10343 543
rect 10285 435 10343 509
rect 10285 401 10297 435
rect 10297 401 10331 435
rect 10331 401 10343 435
rect 10285 395 10343 401
rect 10403 543 10461 549
rect 10403 509 10415 543
rect 10415 509 10449 543
rect 10449 509 10461 543
rect 10403 435 10461 509
rect 10403 401 10415 435
rect 10415 401 10449 435
rect 10449 401 10461 435
rect 10403 395 10461 401
rect 10521 543 10579 549
rect 10521 509 10533 543
rect 10533 509 10567 543
rect 10567 509 10579 543
rect 10521 435 10579 509
rect 10521 401 10533 435
rect 10533 401 10567 435
rect 10567 401 10579 435
rect 10521 395 10579 401
rect 10639 543 10697 549
rect 10639 509 10651 543
rect 10651 509 10685 543
rect 10685 509 10697 543
rect 10639 435 10697 509
rect 10639 401 10651 435
rect 10651 401 10685 435
rect 10685 401 10697 435
rect 10639 395 10697 401
rect 4801 -226 4810 334
rect 4810 -226 4844 334
rect 4844 -226 4853 334
rect 4917 -226 4928 334
rect 4928 -226 4962 334
rect 4962 -226 4969 334
rect 5037 -226 5046 334
rect 5046 -226 5080 334
rect 5080 -226 5089 334
rect 5153 -226 5164 334
rect 5164 -226 5198 334
rect 5198 -226 5205 334
rect 5273 -226 5282 334
rect 5282 -226 5316 334
rect 5316 -226 5325 334
rect 5389 -226 5400 334
rect 5400 -226 5434 334
rect 5434 -226 5441 334
rect 5509 -226 5518 334
rect 5518 -226 5552 334
rect 5552 -226 5561 334
rect 5625 -226 5636 334
rect 5636 -226 5670 334
rect 5670 -226 5677 334
rect 5745 -226 5754 334
rect 5754 -226 5788 334
rect 5788 -226 5797 334
rect 5861 -226 5872 334
rect 5872 -226 5906 334
rect 5906 -226 5913 334
rect 5981 -226 5990 334
rect 5990 -226 6024 334
rect 6024 -226 6033 334
rect 6097 -226 6108 334
rect 6108 -226 6142 334
rect 6142 -226 6149 334
rect 6217 -226 6226 334
rect 6226 -226 6260 334
rect 6260 -226 6269 334
rect 6333 -226 6344 334
rect 6344 -226 6378 334
rect 6378 -226 6385 334
rect 6453 -226 6462 334
rect 6462 -226 6496 334
rect 6496 -226 6505 334
rect 6569 -226 6580 334
rect 6580 -226 6614 334
rect 6614 -226 6621 334
rect 6689 -226 6698 334
rect 6698 -226 6732 334
rect 6732 -226 6741 334
rect 6805 -226 6816 334
rect 6816 -226 6850 334
rect 6850 -226 6857 334
rect 6925 -226 6934 334
rect 6934 -226 6968 334
rect 6968 -226 6977 334
rect 7041 -226 7052 334
rect 7052 -226 7086 334
rect 7086 -226 7093 334
rect 7161 -226 7170 334
rect 7170 -226 7204 334
rect 7204 -226 7213 334
rect 7277 -226 7288 334
rect 7288 -226 7322 334
rect 7322 -226 7329 334
rect 7397 -226 7406 334
rect 7406 -226 7440 334
rect 7440 -226 7449 334
rect 7513 -226 7524 334
rect 7524 -226 7558 334
rect 7558 -226 7565 334
rect 7633 -226 7642 334
rect 7642 -226 7676 334
rect 7676 -226 7685 334
rect 7749 -226 7760 334
rect 7760 -226 7794 334
rect 7794 -226 7801 334
rect 7869 -226 7878 334
rect 7878 -226 7912 334
rect 7912 -226 7921 334
rect 7985 -226 7996 334
rect 7996 -226 8030 334
rect 8030 -226 8037 334
rect 8105 -226 8114 334
rect 8114 -226 8148 334
rect 8148 -226 8157 334
rect 8221 -226 8232 334
rect 8232 -226 8266 334
rect 8266 -226 8273 334
rect 8341 -226 8350 334
rect 8350 -226 8384 334
rect 8384 -226 8393 334
rect 8457 -226 8468 334
rect 8468 -226 8502 334
rect 8502 -226 8509 334
rect 8577 -226 8586 334
rect 8586 -226 8620 334
rect 8620 -226 8629 334
rect 8693 -226 8704 334
rect 8704 -226 8738 334
rect 8738 -226 8745 334
rect 8813 -226 8822 334
rect 8822 -226 8856 334
rect 8856 -226 8865 334
rect 8929 -226 8940 334
rect 8940 -226 8974 334
rect 8974 -226 8981 334
rect 9049 -226 9058 334
rect 9058 -226 9092 334
rect 9092 -226 9101 334
rect 9165 -226 9176 334
rect 9176 -226 9210 334
rect 9210 -226 9217 334
rect 9285 -226 9294 334
rect 9294 -226 9328 334
rect 9328 -226 9337 334
rect 9401 -226 9412 334
rect 9412 -226 9446 334
rect 9446 -226 9453 334
rect 9521 -226 9530 334
rect 9530 -226 9564 334
rect 9564 -226 9573 334
rect 9637 -226 9648 334
rect 9648 -226 9682 334
rect 9682 -226 9689 334
rect 9757 -226 9766 334
rect 9766 -226 9800 334
rect 9800 -226 9809 334
rect 9873 -226 9884 334
rect 9884 -226 9918 334
rect 9918 -226 9925 334
rect 9993 -226 10002 334
rect 10002 -226 10036 334
rect 10036 -226 10045 334
rect 10109 -226 10120 334
rect 10120 -226 10154 334
rect 10154 -226 10161 334
rect 10229 -226 10238 334
rect 10238 -226 10272 334
rect 10272 -226 10281 334
rect 10345 -226 10356 334
rect 10356 -226 10390 334
rect 10390 -226 10397 334
rect 10465 -226 10474 334
rect 10474 -226 10508 334
rect 10508 -226 10517 334
rect 10581 -226 10592 334
rect 10592 -226 10626 334
rect 10626 -226 10633 334
rect 10701 -226 10710 334
rect 10710 -226 10744 334
rect 10744 -226 10753 334
rect 4801 -395 4853 -375
rect 5037 -395 5089 -375
rect 5273 -395 5325 -375
rect 5509 -395 5561 -375
rect 5745 -395 5797 -375
rect 5981 -395 6033 -375
rect 6217 -395 6269 -375
rect 6453 -395 6505 -375
rect 6689 -395 6741 -375
rect 6925 -395 6977 -375
rect 7161 -395 7213 -375
rect 7397 -395 7449 -375
rect 7633 -395 7685 -375
rect 7869 -395 7921 -375
rect 8105 -395 8157 -375
rect 8341 -395 8393 -375
rect 8577 -395 8629 -375
rect 8813 -395 8865 -375
rect 9049 -395 9101 -375
rect 9285 -395 9337 -375
rect 9521 -395 9573 -375
rect 9757 -395 9809 -375
rect 9993 -395 10045 -375
rect 10229 -395 10281 -375
rect 10465 -395 10517 -375
rect 10701 -395 10753 -375
rect 4801 -429 4810 -395
rect 4810 -429 4848 -395
rect 4848 -429 4853 -395
rect 5037 -429 5064 -395
rect 5064 -429 5089 -395
rect 5273 -429 5280 -395
rect 5280 -429 5314 -395
rect 5314 -429 5325 -395
rect 5509 -429 5530 -395
rect 5530 -429 5561 -395
rect 5745 -429 5746 -395
rect 5746 -429 5784 -395
rect 5784 -429 5797 -395
rect 5981 -429 6000 -395
rect 6000 -429 6033 -395
rect 6217 -429 6250 -395
rect 6250 -429 6269 -395
rect 6453 -429 6466 -395
rect 6466 -429 6504 -395
rect 6504 -429 6505 -395
rect 6689 -429 6720 -395
rect 6720 -429 6741 -395
rect 6925 -429 6936 -395
rect 6936 -429 6970 -395
rect 6970 -429 6977 -395
rect 7161 -429 7186 -395
rect 7186 -429 7213 -395
rect 7397 -429 7402 -395
rect 7402 -429 7440 -395
rect 7440 -429 7449 -395
rect 7633 -429 7656 -395
rect 7656 -429 7685 -395
rect 7869 -429 7872 -395
rect 7872 -429 7906 -395
rect 7906 -429 7921 -395
rect 8105 -429 8122 -395
rect 8122 -429 8157 -395
rect 8341 -429 8376 -395
rect 8376 -429 8393 -395
rect 8577 -429 8592 -395
rect 8592 -429 8626 -395
rect 8626 -429 8629 -395
rect 8813 -429 8842 -395
rect 8842 -429 8865 -395
rect 9049 -429 9058 -395
rect 9058 -429 9096 -395
rect 9096 -429 9101 -395
rect 9285 -429 9312 -395
rect 9312 -429 9337 -395
rect 9521 -429 9528 -395
rect 9528 -429 9562 -395
rect 9562 -429 9573 -395
rect 9757 -429 9778 -395
rect 9778 -429 9809 -395
rect 9993 -429 9994 -395
rect 9994 -429 10032 -395
rect 10032 -429 10045 -395
rect 10229 -429 10248 -395
rect 10248 -429 10281 -395
rect 10465 -429 10498 -395
rect 10498 -429 10517 -395
rect 10701 -429 10714 -395
rect 10714 -429 10752 -395
rect 10752 -429 10753 -395
rect 4801 -483 4853 -429
rect 5037 -483 5089 -429
rect 5273 -483 5325 -429
rect 5509 -483 5561 -429
rect 5745 -483 5797 -429
rect 5981 -483 6033 -429
rect 6217 -483 6269 -429
rect 6453 -483 6505 -429
rect 6689 -483 6741 -429
rect 6925 -483 6977 -429
rect 7161 -483 7213 -429
rect 7397 -483 7449 -429
rect 7633 -483 7685 -429
rect 7869 -483 7921 -429
rect 8105 -483 8157 -429
rect 8341 -483 8393 -429
rect 8577 -483 8629 -429
rect 8813 -483 8865 -429
rect 9049 -483 9101 -429
rect 9285 -483 9337 -429
rect 9521 -483 9573 -429
rect 9757 -483 9809 -429
rect 9993 -483 10045 -429
rect 10229 -483 10281 -429
rect 10465 -483 10517 -429
rect 10701 -483 10753 -429
rect 4801 -517 4810 -483
rect 4810 -517 4848 -483
rect 4848 -517 4853 -483
rect 5037 -517 5064 -483
rect 5064 -517 5089 -483
rect 5273 -517 5280 -483
rect 5280 -517 5314 -483
rect 5314 -517 5325 -483
rect 5509 -517 5530 -483
rect 5530 -517 5561 -483
rect 5745 -517 5746 -483
rect 5746 -517 5784 -483
rect 5784 -517 5797 -483
rect 5981 -517 6000 -483
rect 6000 -517 6033 -483
rect 6217 -517 6250 -483
rect 6250 -517 6269 -483
rect 6453 -517 6466 -483
rect 6466 -517 6504 -483
rect 6504 -517 6505 -483
rect 6689 -517 6720 -483
rect 6720 -517 6741 -483
rect 6925 -517 6936 -483
rect 6936 -517 6970 -483
rect 6970 -517 6977 -483
rect 7161 -517 7186 -483
rect 7186 -517 7213 -483
rect 7397 -517 7402 -483
rect 7402 -517 7440 -483
rect 7440 -517 7449 -483
rect 7633 -517 7656 -483
rect 7656 -517 7685 -483
rect 7869 -517 7872 -483
rect 7872 -517 7906 -483
rect 7906 -517 7921 -483
rect 8105 -517 8122 -483
rect 8122 -517 8157 -483
rect 8341 -517 8376 -483
rect 8376 -517 8393 -483
rect 8577 -517 8592 -483
rect 8592 -517 8626 -483
rect 8626 -517 8629 -483
rect 8813 -517 8842 -483
rect 8842 -517 8865 -483
rect 9049 -517 9058 -483
rect 9058 -517 9096 -483
rect 9096 -517 9101 -483
rect 9285 -517 9312 -483
rect 9312 -517 9337 -483
rect 9521 -517 9528 -483
rect 9528 -517 9562 -483
rect 9562 -517 9573 -483
rect 9757 -517 9778 -483
rect 9778 -517 9809 -483
rect 9993 -517 9994 -483
rect 9994 -517 10032 -483
rect 10032 -517 10045 -483
rect 10229 -517 10248 -483
rect 10248 -517 10281 -483
rect 10465 -517 10498 -483
rect 10498 -517 10517 -483
rect 10701 -517 10714 -483
rect 10714 -517 10752 -483
rect 10752 -517 10753 -483
rect 4801 -571 4853 -517
rect 5037 -571 5089 -517
rect 5273 -571 5325 -517
rect 5509 -571 5561 -517
rect 5745 -571 5797 -517
rect 5981 -571 6033 -517
rect 6217 -571 6269 -517
rect 6453 -571 6505 -517
rect 6689 -571 6741 -517
rect 6925 -571 6977 -517
rect 7161 -571 7213 -517
rect 7397 -571 7449 -517
rect 7633 -571 7685 -517
rect 7869 -571 7921 -517
rect 8105 -571 8157 -517
rect 8341 -571 8393 -517
rect 8577 -571 8629 -517
rect 8813 -571 8865 -517
rect 9049 -571 9101 -517
rect 9285 -571 9337 -517
rect 9521 -571 9573 -517
rect 9757 -571 9809 -517
rect 9993 -571 10045 -517
rect 10229 -571 10281 -517
rect 10465 -571 10517 -517
rect 10701 -571 10753 -517
rect 4801 -605 4810 -571
rect 4810 -605 4848 -571
rect 4848 -605 4853 -571
rect 5037 -605 5064 -571
rect 5064 -605 5089 -571
rect 5273 -605 5280 -571
rect 5280 -605 5314 -571
rect 5314 -605 5325 -571
rect 5509 -605 5530 -571
rect 5530 -605 5561 -571
rect 5745 -605 5746 -571
rect 5746 -605 5784 -571
rect 5784 -605 5797 -571
rect 5981 -605 6000 -571
rect 6000 -605 6033 -571
rect 6217 -605 6250 -571
rect 6250 -605 6269 -571
rect 6453 -605 6466 -571
rect 6466 -605 6504 -571
rect 6504 -605 6505 -571
rect 6689 -605 6720 -571
rect 6720 -605 6741 -571
rect 6925 -605 6936 -571
rect 6936 -605 6970 -571
rect 6970 -605 6977 -571
rect 7161 -605 7186 -571
rect 7186 -605 7213 -571
rect 7397 -605 7402 -571
rect 7402 -605 7440 -571
rect 7440 -605 7449 -571
rect 7633 -605 7656 -571
rect 7656 -605 7685 -571
rect 7869 -605 7872 -571
rect 7872 -605 7906 -571
rect 7906 -605 7921 -571
rect 8105 -605 8122 -571
rect 8122 -605 8157 -571
rect 8341 -605 8376 -571
rect 8376 -605 8393 -571
rect 8577 -605 8592 -571
rect 8592 -605 8626 -571
rect 8626 -605 8629 -571
rect 8813 -605 8842 -571
rect 8842 -605 8865 -571
rect 9049 -605 9058 -571
rect 9058 -605 9096 -571
rect 9096 -605 9101 -571
rect 9285 -605 9312 -571
rect 9312 -605 9337 -571
rect 9521 -605 9528 -571
rect 9528 -605 9562 -571
rect 9562 -605 9573 -571
rect 9757 -605 9778 -571
rect 9778 -605 9809 -571
rect 9993 -605 9994 -571
rect 9994 -605 10032 -571
rect 10032 -605 10045 -571
rect 10229 -605 10248 -571
rect 10248 -605 10281 -571
rect 10465 -605 10498 -571
rect 10498 -605 10517 -571
rect 10701 -605 10714 -571
rect 10714 -605 10752 -571
rect 10752 -605 10753 -571
rect 4801 -625 4853 -605
rect 5037 -625 5089 -605
rect 5273 -625 5325 -605
rect 5509 -625 5561 -605
rect 5745 -625 5797 -605
rect 5981 -625 6033 -605
rect 6217 -625 6269 -605
rect 6453 -625 6505 -605
rect 6689 -625 6741 -605
rect 6925 -625 6977 -605
rect 7161 -625 7213 -605
rect 7397 -625 7449 -605
rect 7633 -625 7685 -605
rect 7869 -625 7921 -605
rect 8105 -625 8157 -605
rect 8341 -625 8393 -605
rect 8577 -625 8629 -605
rect 8813 -625 8865 -605
rect 9049 -625 9101 -605
rect 9285 -625 9337 -605
rect 9521 -625 9573 -605
rect 9757 -625 9809 -605
rect 9993 -625 10045 -605
rect 10229 -625 10281 -605
rect 10465 -625 10517 -605
rect 10701 -625 10753 -605
rect 4801 -1440 4810 -880
rect 4810 -1440 4844 -880
rect 4844 -1440 4853 -880
rect 4917 -1440 4928 -880
rect 4928 -1440 4962 -880
rect 4962 -1440 4969 -880
rect 5037 -1440 5046 -880
rect 5046 -1440 5080 -880
rect 5080 -1440 5089 -880
rect 5153 -1440 5164 -880
rect 5164 -1440 5198 -880
rect 5198 -1440 5205 -880
rect 5273 -1440 5282 -880
rect 5282 -1440 5316 -880
rect 5316 -1440 5325 -880
rect 5389 -1440 5400 -880
rect 5400 -1440 5434 -880
rect 5434 -1440 5441 -880
rect 5509 -1440 5518 -880
rect 5518 -1440 5552 -880
rect 5552 -1440 5561 -880
rect 5625 -1440 5636 -880
rect 5636 -1440 5670 -880
rect 5670 -1440 5677 -880
rect 5745 -1440 5754 -880
rect 5754 -1440 5788 -880
rect 5788 -1440 5797 -880
rect 5861 -1440 5872 -880
rect 5872 -1440 5906 -880
rect 5906 -1440 5913 -880
rect 5981 -1440 5990 -880
rect 5990 -1440 6024 -880
rect 6024 -1440 6033 -880
rect 6097 -1440 6108 -880
rect 6108 -1440 6142 -880
rect 6142 -1440 6149 -880
rect 6217 -1440 6226 -880
rect 6226 -1440 6260 -880
rect 6260 -1440 6269 -880
rect 6333 -1440 6344 -880
rect 6344 -1440 6378 -880
rect 6378 -1440 6385 -880
rect 6453 -1440 6462 -880
rect 6462 -1440 6496 -880
rect 6496 -1440 6505 -880
rect 6569 -1440 6580 -880
rect 6580 -1440 6614 -880
rect 6614 -1440 6621 -880
rect 6689 -1440 6698 -880
rect 6698 -1440 6732 -880
rect 6732 -1440 6741 -880
rect 6805 -1440 6816 -880
rect 6816 -1440 6850 -880
rect 6850 -1440 6857 -880
rect 6925 -1440 6934 -880
rect 6934 -1440 6968 -880
rect 6968 -1440 6977 -880
rect 7041 -1440 7052 -880
rect 7052 -1440 7086 -880
rect 7086 -1440 7093 -880
rect 7161 -1440 7170 -880
rect 7170 -1440 7204 -880
rect 7204 -1440 7213 -880
rect 7277 -1440 7288 -880
rect 7288 -1440 7322 -880
rect 7322 -1440 7329 -880
rect 7397 -1440 7406 -880
rect 7406 -1440 7440 -880
rect 7440 -1440 7449 -880
rect 7513 -1440 7524 -880
rect 7524 -1440 7558 -880
rect 7558 -1440 7565 -880
rect 7633 -1440 7642 -880
rect 7642 -1440 7676 -880
rect 7676 -1440 7685 -880
rect 7749 -1440 7760 -880
rect 7760 -1440 7794 -880
rect 7794 -1440 7801 -880
rect 7869 -1440 7878 -880
rect 7878 -1440 7912 -880
rect 7912 -1440 7921 -880
rect 7985 -1440 7996 -880
rect 7996 -1440 8030 -880
rect 8030 -1440 8037 -880
rect 8105 -1440 8114 -880
rect 8114 -1440 8148 -880
rect 8148 -1440 8157 -880
rect 8221 -1440 8232 -880
rect 8232 -1440 8266 -880
rect 8266 -1440 8273 -880
rect 8341 -1440 8350 -880
rect 8350 -1440 8384 -880
rect 8384 -1440 8393 -880
rect 8457 -1440 8468 -880
rect 8468 -1440 8502 -880
rect 8502 -1440 8509 -880
rect 8577 -1440 8586 -880
rect 8586 -1440 8620 -880
rect 8620 -1440 8629 -880
rect 8693 -1440 8704 -880
rect 8704 -1440 8738 -880
rect 8738 -1440 8745 -880
rect 8813 -1440 8822 -880
rect 8822 -1440 8856 -880
rect 8856 -1440 8865 -880
rect 8929 -1440 8940 -880
rect 8940 -1440 8974 -880
rect 8974 -1440 8981 -880
rect 9049 -1440 9058 -880
rect 9058 -1440 9092 -880
rect 9092 -1440 9101 -880
rect 9165 -1440 9176 -880
rect 9176 -1440 9210 -880
rect 9210 -1440 9217 -880
rect 9285 -1440 9294 -880
rect 9294 -1440 9328 -880
rect 9328 -1440 9337 -880
rect 9401 -1440 9412 -880
rect 9412 -1440 9446 -880
rect 9446 -1440 9453 -880
rect 9521 -1440 9530 -880
rect 9530 -1440 9564 -880
rect 9564 -1440 9573 -880
rect 9637 -1440 9648 -880
rect 9648 -1440 9682 -880
rect 9682 -1440 9689 -880
rect 9757 -1440 9766 -880
rect 9766 -1440 9800 -880
rect 9800 -1440 9809 -880
rect 9873 -1440 9884 -880
rect 9884 -1440 9918 -880
rect 9918 -1440 9925 -880
rect 9993 -1440 10002 -880
rect 10002 -1440 10036 -880
rect 10036 -1440 10045 -880
rect 10109 -1440 10120 -880
rect 10120 -1440 10154 -880
rect 10154 -1440 10161 -880
rect 10229 -1440 10238 -880
rect 10238 -1440 10272 -880
rect 10272 -1440 10281 -880
rect 10345 -1440 10356 -880
rect 10356 -1440 10390 -880
rect 10390 -1440 10397 -880
rect 10465 -1440 10474 -880
rect 10474 -1440 10508 -880
rect 10508 -1440 10517 -880
rect 10581 -1440 10592 -880
rect 10592 -1440 10626 -880
rect 10626 -1440 10633 -880
rect 10701 -1440 10710 -880
rect 10710 -1440 10744 -880
rect 10744 -1440 10753 -880
rect 4857 -1507 4915 -1501
rect 4857 -1541 4869 -1507
rect 4869 -1541 4903 -1507
rect 4903 -1541 4915 -1507
rect 4857 -1615 4915 -1541
rect 4857 -1649 4869 -1615
rect 4869 -1649 4903 -1615
rect 4903 -1649 4915 -1615
rect 4857 -1655 4915 -1649
rect 4975 -1507 5033 -1501
rect 4975 -1541 4987 -1507
rect 4987 -1541 5021 -1507
rect 5021 -1541 5033 -1507
rect 4975 -1615 5033 -1541
rect 4975 -1649 4987 -1615
rect 4987 -1649 5021 -1615
rect 5021 -1649 5033 -1615
rect 4975 -1655 5033 -1649
rect 5093 -1507 5151 -1501
rect 5093 -1541 5105 -1507
rect 5105 -1541 5139 -1507
rect 5139 -1541 5151 -1507
rect 5093 -1615 5151 -1541
rect 5093 -1649 5105 -1615
rect 5105 -1649 5139 -1615
rect 5139 -1649 5151 -1615
rect 5093 -1655 5151 -1649
rect 5211 -1507 5269 -1501
rect 5211 -1541 5223 -1507
rect 5223 -1541 5257 -1507
rect 5257 -1541 5269 -1507
rect 5211 -1615 5269 -1541
rect 5211 -1649 5223 -1615
rect 5223 -1649 5257 -1615
rect 5257 -1649 5269 -1615
rect 5211 -1655 5269 -1649
rect 5329 -1507 5387 -1501
rect 5329 -1541 5341 -1507
rect 5341 -1541 5375 -1507
rect 5375 -1541 5387 -1507
rect 5329 -1615 5387 -1541
rect 5329 -1649 5341 -1615
rect 5341 -1649 5375 -1615
rect 5375 -1649 5387 -1615
rect 5329 -1655 5387 -1649
rect 5447 -1507 5505 -1501
rect 5447 -1541 5459 -1507
rect 5459 -1541 5493 -1507
rect 5493 -1541 5505 -1507
rect 5447 -1615 5505 -1541
rect 5447 -1649 5459 -1615
rect 5459 -1649 5493 -1615
rect 5493 -1649 5505 -1615
rect 5447 -1655 5505 -1649
rect 5565 -1507 5623 -1501
rect 5565 -1541 5577 -1507
rect 5577 -1541 5611 -1507
rect 5611 -1541 5623 -1507
rect 5565 -1615 5623 -1541
rect 5565 -1649 5577 -1615
rect 5577 -1649 5611 -1615
rect 5611 -1649 5623 -1615
rect 5565 -1655 5623 -1649
rect 5683 -1507 5741 -1501
rect 5683 -1541 5695 -1507
rect 5695 -1541 5729 -1507
rect 5729 -1541 5741 -1507
rect 5683 -1615 5741 -1541
rect 5683 -1649 5695 -1615
rect 5695 -1649 5729 -1615
rect 5729 -1649 5741 -1615
rect 5683 -1655 5741 -1649
rect 5801 -1507 5859 -1501
rect 5801 -1541 5813 -1507
rect 5813 -1541 5847 -1507
rect 5847 -1541 5859 -1507
rect 5801 -1615 5859 -1541
rect 5801 -1649 5813 -1615
rect 5813 -1649 5847 -1615
rect 5847 -1649 5859 -1615
rect 5801 -1655 5859 -1649
rect 5919 -1507 5977 -1501
rect 5919 -1541 5931 -1507
rect 5931 -1541 5965 -1507
rect 5965 -1541 5977 -1507
rect 5919 -1615 5977 -1541
rect 5919 -1649 5931 -1615
rect 5931 -1649 5965 -1615
rect 5965 -1649 5977 -1615
rect 5919 -1655 5977 -1649
rect 6037 -1507 6095 -1501
rect 6037 -1541 6049 -1507
rect 6049 -1541 6083 -1507
rect 6083 -1541 6095 -1507
rect 6037 -1615 6095 -1541
rect 6037 -1649 6049 -1615
rect 6049 -1649 6083 -1615
rect 6083 -1649 6095 -1615
rect 6037 -1655 6095 -1649
rect 6155 -1507 6213 -1501
rect 6155 -1541 6167 -1507
rect 6167 -1541 6201 -1507
rect 6201 -1541 6213 -1507
rect 6155 -1615 6213 -1541
rect 6155 -1649 6167 -1615
rect 6167 -1649 6201 -1615
rect 6201 -1649 6213 -1615
rect 6155 -1655 6213 -1649
rect 6273 -1507 6331 -1501
rect 6273 -1541 6285 -1507
rect 6285 -1541 6319 -1507
rect 6319 -1541 6331 -1507
rect 6273 -1615 6331 -1541
rect 6273 -1649 6285 -1615
rect 6285 -1649 6319 -1615
rect 6319 -1649 6331 -1615
rect 6273 -1655 6331 -1649
rect 6391 -1507 6449 -1501
rect 6391 -1541 6403 -1507
rect 6403 -1541 6437 -1507
rect 6437 -1541 6449 -1507
rect 6391 -1615 6449 -1541
rect 6391 -1649 6403 -1615
rect 6403 -1649 6437 -1615
rect 6437 -1649 6449 -1615
rect 6391 -1655 6449 -1649
rect 6509 -1507 6567 -1501
rect 6509 -1541 6521 -1507
rect 6521 -1541 6555 -1507
rect 6555 -1541 6567 -1507
rect 6509 -1615 6567 -1541
rect 6509 -1649 6521 -1615
rect 6521 -1649 6555 -1615
rect 6555 -1649 6567 -1615
rect 6509 -1655 6567 -1649
rect 6627 -1507 6685 -1501
rect 6627 -1541 6639 -1507
rect 6639 -1541 6673 -1507
rect 6673 -1541 6685 -1507
rect 6627 -1615 6685 -1541
rect 6627 -1649 6639 -1615
rect 6639 -1649 6673 -1615
rect 6673 -1649 6685 -1615
rect 6627 -1655 6685 -1649
rect 6745 -1507 6803 -1501
rect 6745 -1541 6757 -1507
rect 6757 -1541 6791 -1507
rect 6791 -1541 6803 -1507
rect 6745 -1615 6803 -1541
rect 6745 -1649 6757 -1615
rect 6757 -1649 6791 -1615
rect 6791 -1649 6803 -1615
rect 6745 -1655 6803 -1649
rect 6863 -1507 6921 -1501
rect 6863 -1541 6875 -1507
rect 6875 -1541 6909 -1507
rect 6909 -1541 6921 -1507
rect 6863 -1615 6921 -1541
rect 6863 -1649 6875 -1615
rect 6875 -1649 6909 -1615
rect 6909 -1649 6921 -1615
rect 6863 -1655 6921 -1649
rect 6981 -1507 7039 -1501
rect 6981 -1541 6993 -1507
rect 6993 -1541 7027 -1507
rect 7027 -1541 7039 -1507
rect 6981 -1615 7039 -1541
rect 6981 -1649 6993 -1615
rect 6993 -1649 7027 -1615
rect 7027 -1649 7039 -1615
rect 6981 -1655 7039 -1649
rect 7099 -1507 7157 -1501
rect 7099 -1541 7111 -1507
rect 7111 -1541 7145 -1507
rect 7145 -1541 7157 -1507
rect 7099 -1615 7157 -1541
rect 7099 -1649 7111 -1615
rect 7111 -1649 7145 -1615
rect 7145 -1649 7157 -1615
rect 7099 -1655 7157 -1649
rect 7217 -1507 7275 -1501
rect 7217 -1541 7229 -1507
rect 7229 -1541 7263 -1507
rect 7263 -1541 7275 -1507
rect 7217 -1615 7275 -1541
rect 7217 -1649 7229 -1615
rect 7229 -1649 7263 -1615
rect 7263 -1649 7275 -1615
rect 7217 -1655 7275 -1649
rect 7335 -1507 7393 -1501
rect 7335 -1541 7347 -1507
rect 7347 -1541 7381 -1507
rect 7381 -1541 7393 -1507
rect 7335 -1615 7393 -1541
rect 7335 -1649 7347 -1615
rect 7347 -1649 7381 -1615
rect 7381 -1649 7393 -1615
rect 7335 -1655 7393 -1649
rect 7453 -1507 7511 -1501
rect 7453 -1541 7465 -1507
rect 7465 -1541 7499 -1507
rect 7499 -1541 7511 -1507
rect 7453 -1615 7511 -1541
rect 7453 -1649 7465 -1615
rect 7465 -1649 7499 -1615
rect 7499 -1649 7511 -1615
rect 7453 -1655 7511 -1649
rect 7571 -1507 7629 -1501
rect 7571 -1541 7583 -1507
rect 7583 -1541 7617 -1507
rect 7617 -1541 7629 -1507
rect 7571 -1615 7629 -1541
rect 7571 -1649 7583 -1615
rect 7583 -1649 7617 -1615
rect 7617 -1649 7629 -1615
rect 7571 -1655 7629 -1649
rect 7689 -1507 7747 -1501
rect 7689 -1541 7701 -1507
rect 7701 -1541 7735 -1507
rect 7735 -1541 7747 -1507
rect 7689 -1615 7747 -1541
rect 7689 -1649 7701 -1615
rect 7701 -1649 7735 -1615
rect 7735 -1649 7747 -1615
rect 7689 -1655 7747 -1649
rect 7807 -1507 7865 -1501
rect 7807 -1541 7819 -1507
rect 7819 -1541 7853 -1507
rect 7853 -1541 7865 -1507
rect 7807 -1615 7865 -1541
rect 7807 -1649 7819 -1615
rect 7819 -1649 7853 -1615
rect 7853 -1649 7865 -1615
rect 7807 -1655 7865 -1649
rect 7925 -1507 7983 -1501
rect 7925 -1541 7937 -1507
rect 7937 -1541 7971 -1507
rect 7971 -1541 7983 -1507
rect 7925 -1615 7983 -1541
rect 7925 -1649 7937 -1615
rect 7937 -1649 7971 -1615
rect 7971 -1649 7983 -1615
rect 7925 -1655 7983 -1649
rect 8043 -1507 8101 -1501
rect 8043 -1541 8055 -1507
rect 8055 -1541 8089 -1507
rect 8089 -1541 8101 -1507
rect 8043 -1615 8101 -1541
rect 8043 -1649 8055 -1615
rect 8055 -1649 8089 -1615
rect 8089 -1649 8101 -1615
rect 8043 -1655 8101 -1649
rect 8161 -1507 8219 -1501
rect 8161 -1541 8173 -1507
rect 8173 -1541 8207 -1507
rect 8207 -1541 8219 -1507
rect 8161 -1615 8219 -1541
rect 8161 -1649 8173 -1615
rect 8173 -1649 8207 -1615
rect 8207 -1649 8219 -1615
rect 8161 -1655 8219 -1649
rect 8279 -1507 8337 -1501
rect 8279 -1541 8291 -1507
rect 8291 -1541 8325 -1507
rect 8325 -1541 8337 -1507
rect 8279 -1615 8337 -1541
rect 8279 -1649 8291 -1615
rect 8291 -1649 8325 -1615
rect 8325 -1649 8337 -1615
rect 8279 -1655 8337 -1649
rect 8397 -1507 8455 -1501
rect 8397 -1541 8409 -1507
rect 8409 -1541 8443 -1507
rect 8443 -1541 8455 -1507
rect 8397 -1615 8455 -1541
rect 8397 -1649 8409 -1615
rect 8409 -1649 8443 -1615
rect 8443 -1649 8455 -1615
rect 8397 -1655 8455 -1649
rect 8515 -1507 8573 -1501
rect 8515 -1541 8527 -1507
rect 8527 -1541 8561 -1507
rect 8561 -1541 8573 -1507
rect 8515 -1615 8573 -1541
rect 8515 -1649 8527 -1615
rect 8527 -1649 8561 -1615
rect 8561 -1649 8573 -1615
rect 8515 -1655 8573 -1649
rect 8633 -1507 8691 -1501
rect 8633 -1541 8645 -1507
rect 8645 -1541 8679 -1507
rect 8679 -1541 8691 -1507
rect 8633 -1615 8691 -1541
rect 8633 -1649 8645 -1615
rect 8645 -1649 8679 -1615
rect 8679 -1649 8691 -1615
rect 8633 -1655 8691 -1649
rect 8751 -1507 8809 -1501
rect 8751 -1541 8763 -1507
rect 8763 -1541 8797 -1507
rect 8797 -1541 8809 -1507
rect 8751 -1615 8809 -1541
rect 8751 -1649 8763 -1615
rect 8763 -1649 8797 -1615
rect 8797 -1649 8809 -1615
rect 8751 -1655 8809 -1649
rect 8869 -1507 8927 -1501
rect 8869 -1541 8881 -1507
rect 8881 -1541 8915 -1507
rect 8915 -1541 8927 -1507
rect 8869 -1615 8927 -1541
rect 8869 -1649 8881 -1615
rect 8881 -1649 8915 -1615
rect 8915 -1649 8927 -1615
rect 8869 -1655 8927 -1649
rect 8987 -1507 9045 -1501
rect 8987 -1541 8999 -1507
rect 8999 -1541 9033 -1507
rect 9033 -1541 9045 -1507
rect 8987 -1615 9045 -1541
rect 8987 -1649 8999 -1615
rect 8999 -1649 9033 -1615
rect 9033 -1649 9045 -1615
rect 8987 -1655 9045 -1649
rect 9105 -1507 9163 -1501
rect 9105 -1541 9117 -1507
rect 9117 -1541 9151 -1507
rect 9151 -1541 9163 -1507
rect 9105 -1615 9163 -1541
rect 9105 -1649 9117 -1615
rect 9117 -1649 9151 -1615
rect 9151 -1649 9163 -1615
rect 9105 -1655 9163 -1649
rect 9223 -1507 9281 -1501
rect 9223 -1541 9235 -1507
rect 9235 -1541 9269 -1507
rect 9269 -1541 9281 -1507
rect 9223 -1615 9281 -1541
rect 9223 -1649 9235 -1615
rect 9235 -1649 9269 -1615
rect 9269 -1649 9281 -1615
rect 9223 -1655 9281 -1649
rect 9341 -1507 9399 -1501
rect 9341 -1541 9353 -1507
rect 9353 -1541 9387 -1507
rect 9387 -1541 9399 -1507
rect 9341 -1615 9399 -1541
rect 9341 -1649 9353 -1615
rect 9353 -1649 9387 -1615
rect 9387 -1649 9399 -1615
rect 9341 -1655 9399 -1649
rect 9459 -1507 9517 -1501
rect 9459 -1541 9471 -1507
rect 9471 -1541 9505 -1507
rect 9505 -1541 9517 -1507
rect 9459 -1615 9517 -1541
rect 9459 -1649 9471 -1615
rect 9471 -1649 9505 -1615
rect 9505 -1649 9517 -1615
rect 9459 -1655 9517 -1649
rect 9577 -1507 9635 -1501
rect 9577 -1541 9589 -1507
rect 9589 -1541 9623 -1507
rect 9623 -1541 9635 -1507
rect 9577 -1615 9635 -1541
rect 9577 -1649 9589 -1615
rect 9589 -1649 9623 -1615
rect 9623 -1649 9635 -1615
rect 9577 -1655 9635 -1649
rect 9695 -1507 9753 -1501
rect 9695 -1541 9707 -1507
rect 9707 -1541 9741 -1507
rect 9741 -1541 9753 -1507
rect 9695 -1615 9753 -1541
rect 9695 -1649 9707 -1615
rect 9707 -1649 9741 -1615
rect 9741 -1649 9753 -1615
rect 9695 -1655 9753 -1649
rect 9813 -1507 9871 -1501
rect 9813 -1541 9825 -1507
rect 9825 -1541 9859 -1507
rect 9859 -1541 9871 -1507
rect 9813 -1615 9871 -1541
rect 9813 -1649 9825 -1615
rect 9825 -1649 9859 -1615
rect 9859 -1649 9871 -1615
rect 9813 -1655 9871 -1649
rect 9931 -1507 9989 -1501
rect 9931 -1541 9943 -1507
rect 9943 -1541 9977 -1507
rect 9977 -1541 9989 -1507
rect 9931 -1615 9989 -1541
rect 9931 -1649 9943 -1615
rect 9943 -1649 9977 -1615
rect 9977 -1649 9989 -1615
rect 9931 -1655 9989 -1649
rect 10049 -1507 10107 -1501
rect 10049 -1541 10061 -1507
rect 10061 -1541 10095 -1507
rect 10095 -1541 10107 -1507
rect 10049 -1615 10107 -1541
rect 10049 -1649 10061 -1615
rect 10061 -1649 10095 -1615
rect 10095 -1649 10107 -1615
rect 10049 -1655 10107 -1649
rect 10167 -1507 10225 -1501
rect 10167 -1541 10179 -1507
rect 10179 -1541 10213 -1507
rect 10213 -1541 10225 -1507
rect 10167 -1615 10225 -1541
rect 10167 -1649 10179 -1615
rect 10179 -1649 10213 -1615
rect 10213 -1649 10225 -1615
rect 10167 -1655 10225 -1649
rect 10285 -1507 10343 -1501
rect 10285 -1541 10297 -1507
rect 10297 -1541 10331 -1507
rect 10331 -1541 10343 -1507
rect 10285 -1615 10343 -1541
rect 10285 -1649 10297 -1615
rect 10297 -1649 10331 -1615
rect 10331 -1649 10343 -1615
rect 10285 -1655 10343 -1649
rect 10403 -1507 10461 -1501
rect 10403 -1541 10415 -1507
rect 10415 -1541 10449 -1507
rect 10449 -1541 10461 -1507
rect 10403 -1615 10461 -1541
rect 10403 -1649 10415 -1615
rect 10415 -1649 10449 -1615
rect 10449 -1649 10461 -1615
rect 10403 -1655 10461 -1649
rect 10521 -1507 10579 -1501
rect 10521 -1541 10533 -1507
rect 10533 -1541 10567 -1507
rect 10567 -1541 10579 -1507
rect 10521 -1615 10579 -1541
rect 10521 -1649 10533 -1615
rect 10533 -1649 10567 -1615
rect 10567 -1649 10579 -1615
rect 10521 -1655 10579 -1649
rect 10639 -1507 10697 -1501
rect 10639 -1541 10651 -1507
rect 10651 -1541 10685 -1507
rect 10685 -1541 10697 -1507
rect 10639 -1615 10697 -1541
rect 10639 -1649 10651 -1615
rect 10651 -1649 10685 -1615
rect 10685 -1649 10697 -1615
rect 10639 -1655 10697 -1649
rect 4801 -2276 4810 -1716
rect 4810 -2276 4844 -1716
rect 4844 -2276 4853 -1716
rect 4917 -2276 4928 -1716
rect 4928 -2276 4962 -1716
rect 4962 -2276 4969 -1716
rect 5037 -2276 5046 -1716
rect 5046 -2276 5080 -1716
rect 5080 -2276 5089 -1716
rect 5153 -2276 5164 -1716
rect 5164 -2276 5198 -1716
rect 5198 -2276 5205 -1716
rect 5273 -2276 5282 -1716
rect 5282 -2276 5316 -1716
rect 5316 -2276 5325 -1716
rect 5389 -2276 5400 -1716
rect 5400 -2276 5434 -1716
rect 5434 -2276 5441 -1716
rect 5509 -2276 5518 -1716
rect 5518 -2276 5552 -1716
rect 5552 -2276 5561 -1716
rect 5625 -2276 5636 -1716
rect 5636 -2276 5670 -1716
rect 5670 -2276 5677 -1716
rect 5745 -2276 5754 -1716
rect 5754 -2276 5788 -1716
rect 5788 -2276 5797 -1716
rect 5861 -2276 5872 -1716
rect 5872 -2276 5906 -1716
rect 5906 -2276 5913 -1716
rect 5981 -2276 5990 -1716
rect 5990 -2276 6024 -1716
rect 6024 -2276 6033 -1716
rect 6097 -2276 6108 -1716
rect 6108 -2276 6142 -1716
rect 6142 -2276 6149 -1716
rect 6217 -2276 6226 -1716
rect 6226 -2276 6260 -1716
rect 6260 -2276 6269 -1716
rect 6333 -2276 6344 -1716
rect 6344 -2276 6378 -1716
rect 6378 -2276 6385 -1716
rect 6453 -2276 6462 -1716
rect 6462 -2276 6496 -1716
rect 6496 -2276 6505 -1716
rect 6569 -2276 6580 -1716
rect 6580 -2276 6614 -1716
rect 6614 -2276 6621 -1716
rect 6689 -2276 6698 -1716
rect 6698 -2276 6732 -1716
rect 6732 -2276 6741 -1716
rect 6805 -2276 6816 -1716
rect 6816 -2276 6850 -1716
rect 6850 -2276 6857 -1716
rect 6925 -2276 6934 -1716
rect 6934 -2276 6968 -1716
rect 6968 -2276 6977 -1716
rect 7041 -2276 7052 -1716
rect 7052 -2276 7086 -1716
rect 7086 -2276 7093 -1716
rect 7161 -2276 7170 -1716
rect 7170 -2276 7204 -1716
rect 7204 -2276 7213 -1716
rect 7277 -2276 7288 -1716
rect 7288 -2276 7322 -1716
rect 7322 -2276 7329 -1716
rect 7397 -2276 7406 -1716
rect 7406 -2276 7440 -1716
rect 7440 -2276 7449 -1716
rect 7513 -2276 7524 -1716
rect 7524 -2276 7558 -1716
rect 7558 -2276 7565 -1716
rect 7633 -2276 7642 -1716
rect 7642 -2276 7676 -1716
rect 7676 -2276 7685 -1716
rect 7749 -2276 7760 -1716
rect 7760 -2276 7794 -1716
rect 7794 -2276 7801 -1716
rect 7869 -2276 7878 -1716
rect 7878 -2276 7912 -1716
rect 7912 -2276 7921 -1716
rect 7985 -2276 7996 -1716
rect 7996 -2276 8030 -1716
rect 8030 -2276 8037 -1716
rect 8105 -2276 8114 -1716
rect 8114 -2276 8148 -1716
rect 8148 -2276 8157 -1716
rect 8221 -2276 8232 -1716
rect 8232 -2276 8266 -1716
rect 8266 -2276 8273 -1716
rect 8341 -2276 8350 -1716
rect 8350 -2276 8384 -1716
rect 8384 -2276 8393 -1716
rect 8457 -2276 8468 -1716
rect 8468 -2276 8502 -1716
rect 8502 -2276 8509 -1716
rect 8577 -2276 8586 -1716
rect 8586 -2276 8620 -1716
rect 8620 -2276 8629 -1716
rect 8693 -2276 8704 -1716
rect 8704 -2276 8738 -1716
rect 8738 -2276 8745 -1716
rect 8813 -2276 8822 -1716
rect 8822 -2276 8856 -1716
rect 8856 -2276 8865 -1716
rect 8929 -2276 8940 -1716
rect 8940 -2276 8974 -1716
rect 8974 -2276 8981 -1716
rect 9049 -2276 9058 -1716
rect 9058 -2276 9092 -1716
rect 9092 -2276 9101 -1716
rect 9165 -2276 9176 -1716
rect 9176 -2276 9210 -1716
rect 9210 -2276 9217 -1716
rect 9285 -2276 9294 -1716
rect 9294 -2276 9328 -1716
rect 9328 -2276 9337 -1716
rect 9401 -2276 9412 -1716
rect 9412 -2276 9446 -1716
rect 9446 -2276 9453 -1716
rect 9521 -2276 9530 -1716
rect 9530 -2276 9564 -1716
rect 9564 -2276 9573 -1716
rect 9637 -2276 9648 -1716
rect 9648 -2276 9682 -1716
rect 9682 -2276 9689 -1716
rect 9757 -2276 9766 -1716
rect 9766 -2276 9800 -1716
rect 9800 -2276 9809 -1716
rect 9873 -2276 9884 -1716
rect 9884 -2276 9918 -1716
rect 9918 -2276 9925 -1716
rect 9993 -2276 10002 -1716
rect 10002 -2276 10036 -1716
rect 10036 -2276 10045 -1716
rect 10109 -2276 10120 -1716
rect 10120 -2276 10154 -1716
rect 10154 -2276 10161 -1716
rect 10229 -2276 10238 -1716
rect 10238 -2276 10272 -1716
rect 10272 -2276 10281 -1716
rect 10345 -2276 10356 -1716
rect 10356 -2276 10390 -1716
rect 10390 -2276 10397 -1716
rect 10465 -2276 10474 -1716
rect 10474 -2276 10508 -1716
rect 10508 -2276 10517 -1716
rect 10581 -2276 10592 -1716
rect 10592 -2276 10626 -1716
rect 10626 -2276 10633 -1716
rect 10701 -2276 10710 -1716
rect 10710 -2276 10744 -1716
rect 10744 -2276 10753 -1716
rect 4801 -2445 4853 -2425
rect 5037 -2445 5089 -2425
rect 5273 -2445 5325 -2425
rect 5509 -2445 5561 -2425
rect 5745 -2445 5797 -2425
rect 5981 -2445 6033 -2425
rect 6217 -2445 6269 -2425
rect 6453 -2445 6505 -2425
rect 6689 -2445 6741 -2425
rect 6925 -2445 6977 -2425
rect 7161 -2445 7213 -2425
rect 7397 -2445 7449 -2425
rect 7633 -2445 7685 -2425
rect 7869 -2445 7921 -2425
rect 8105 -2445 8157 -2425
rect 8341 -2445 8393 -2425
rect 8577 -2445 8629 -2425
rect 8813 -2445 8865 -2425
rect 9049 -2445 9101 -2425
rect 9285 -2445 9337 -2425
rect 9521 -2445 9573 -2425
rect 9757 -2445 9809 -2425
rect 9993 -2445 10045 -2425
rect 10229 -2445 10281 -2425
rect 10465 -2445 10517 -2425
rect 10701 -2445 10753 -2425
rect 4801 -2479 4810 -2445
rect 4810 -2479 4848 -2445
rect 4848 -2479 4853 -2445
rect 5037 -2479 5064 -2445
rect 5064 -2479 5089 -2445
rect 5273 -2479 5280 -2445
rect 5280 -2479 5314 -2445
rect 5314 -2479 5325 -2445
rect 5509 -2479 5530 -2445
rect 5530 -2479 5561 -2445
rect 5745 -2479 5746 -2445
rect 5746 -2479 5784 -2445
rect 5784 -2479 5797 -2445
rect 5981 -2479 6000 -2445
rect 6000 -2479 6033 -2445
rect 6217 -2479 6250 -2445
rect 6250 -2479 6269 -2445
rect 6453 -2479 6466 -2445
rect 6466 -2479 6504 -2445
rect 6504 -2479 6505 -2445
rect 6689 -2479 6720 -2445
rect 6720 -2479 6741 -2445
rect 6925 -2479 6936 -2445
rect 6936 -2479 6970 -2445
rect 6970 -2479 6977 -2445
rect 7161 -2479 7186 -2445
rect 7186 -2479 7213 -2445
rect 7397 -2479 7402 -2445
rect 7402 -2479 7440 -2445
rect 7440 -2479 7449 -2445
rect 7633 -2479 7656 -2445
rect 7656 -2479 7685 -2445
rect 7869 -2479 7872 -2445
rect 7872 -2479 7906 -2445
rect 7906 -2479 7921 -2445
rect 8105 -2479 8122 -2445
rect 8122 -2479 8157 -2445
rect 8341 -2479 8376 -2445
rect 8376 -2479 8393 -2445
rect 8577 -2479 8592 -2445
rect 8592 -2479 8626 -2445
rect 8626 -2479 8629 -2445
rect 8813 -2479 8842 -2445
rect 8842 -2479 8865 -2445
rect 9049 -2479 9058 -2445
rect 9058 -2479 9096 -2445
rect 9096 -2479 9101 -2445
rect 9285 -2479 9312 -2445
rect 9312 -2479 9337 -2445
rect 9521 -2479 9528 -2445
rect 9528 -2479 9562 -2445
rect 9562 -2479 9573 -2445
rect 9757 -2479 9778 -2445
rect 9778 -2479 9809 -2445
rect 9993 -2479 9994 -2445
rect 9994 -2479 10032 -2445
rect 10032 -2479 10045 -2445
rect 10229 -2479 10248 -2445
rect 10248 -2479 10281 -2445
rect 10465 -2479 10498 -2445
rect 10498 -2479 10517 -2445
rect 10701 -2479 10714 -2445
rect 10714 -2479 10752 -2445
rect 10752 -2479 10753 -2445
rect 4801 -2533 4853 -2479
rect 5037 -2533 5089 -2479
rect 5273 -2533 5325 -2479
rect 5509 -2533 5561 -2479
rect 5745 -2533 5797 -2479
rect 5981 -2533 6033 -2479
rect 6217 -2533 6269 -2479
rect 6453 -2533 6505 -2479
rect 6689 -2533 6741 -2479
rect 6925 -2533 6977 -2479
rect 7161 -2533 7213 -2479
rect 7397 -2533 7449 -2479
rect 7633 -2533 7685 -2479
rect 7869 -2533 7921 -2479
rect 8105 -2533 8157 -2479
rect 8341 -2533 8393 -2479
rect 8577 -2533 8629 -2479
rect 8813 -2533 8865 -2479
rect 9049 -2533 9101 -2479
rect 9285 -2533 9337 -2479
rect 9521 -2533 9573 -2479
rect 9757 -2533 9809 -2479
rect 9993 -2533 10045 -2479
rect 10229 -2533 10281 -2479
rect 10465 -2533 10517 -2479
rect 10701 -2533 10753 -2479
rect 4801 -2567 4810 -2533
rect 4810 -2567 4848 -2533
rect 4848 -2567 4853 -2533
rect 5037 -2567 5064 -2533
rect 5064 -2567 5089 -2533
rect 5273 -2567 5280 -2533
rect 5280 -2567 5314 -2533
rect 5314 -2567 5325 -2533
rect 5509 -2567 5530 -2533
rect 5530 -2567 5561 -2533
rect 5745 -2567 5746 -2533
rect 5746 -2567 5784 -2533
rect 5784 -2567 5797 -2533
rect 5981 -2567 6000 -2533
rect 6000 -2567 6033 -2533
rect 6217 -2567 6250 -2533
rect 6250 -2567 6269 -2533
rect 6453 -2567 6466 -2533
rect 6466 -2567 6504 -2533
rect 6504 -2567 6505 -2533
rect 6689 -2567 6720 -2533
rect 6720 -2567 6741 -2533
rect 6925 -2567 6936 -2533
rect 6936 -2567 6970 -2533
rect 6970 -2567 6977 -2533
rect 7161 -2567 7186 -2533
rect 7186 -2567 7213 -2533
rect 7397 -2567 7402 -2533
rect 7402 -2567 7440 -2533
rect 7440 -2567 7449 -2533
rect 7633 -2567 7656 -2533
rect 7656 -2567 7685 -2533
rect 7869 -2567 7872 -2533
rect 7872 -2567 7906 -2533
rect 7906 -2567 7921 -2533
rect 8105 -2567 8122 -2533
rect 8122 -2567 8157 -2533
rect 8341 -2567 8376 -2533
rect 8376 -2567 8393 -2533
rect 8577 -2567 8592 -2533
rect 8592 -2567 8626 -2533
rect 8626 -2567 8629 -2533
rect 8813 -2567 8842 -2533
rect 8842 -2567 8865 -2533
rect 9049 -2567 9058 -2533
rect 9058 -2567 9096 -2533
rect 9096 -2567 9101 -2533
rect 9285 -2567 9312 -2533
rect 9312 -2567 9337 -2533
rect 9521 -2567 9528 -2533
rect 9528 -2567 9562 -2533
rect 9562 -2567 9573 -2533
rect 9757 -2567 9778 -2533
rect 9778 -2567 9809 -2533
rect 9993 -2567 9994 -2533
rect 9994 -2567 10032 -2533
rect 10032 -2567 10045 -2533
rect 10229 -2567 10248 -2533
rect 10248 -2567 10281 -2533
rect 10465 -2567 10498 -2533
rect 10498 -2567 10517 -2533
rect 10701 -2567 10714 -2533
rect 10714 -2567 10752 -2533
rect 10752 -2567 10753 -2533
rect 4801 -2621 4853 -2567
rect 5037 -2621 5089 -2567
rect 5273 -2621 5325 -2567
rect 5509 -2621 5561 -2567
rect 5745 -2621 5797 -2567
rect 5981 -2621 6033 -2567
rect 6217 -2621 6269 -2567
rect 6453 -2621 6505 -2567
rect 6689 -2621 6741 -2567
rect 6925 -2621 6977 -2567
rect 7161 -2621 7213 -2567
rect 7397 -2621 7449 -2567
rect 7633 -2621 7685 -2567
rect 7869 -2621 7921 -2567
rect 8105 -2621 8157 -2567
rect 8341 -2621 8393 -2567
rect 8577 -2621 8629 -2567
rect 8813 -2621 8865 -2567
rect 9049 -2621 9101 -2567
rect 9285 -2621 9337 -2567
rect 9521 -2621 9573 -2567
rect 9757 -2621 9809 -2567
rect 9993 -2621 10045 -2567
rect 10229 -2621 10281 -2567
rect 10465 -2621 10517 -2567
rect 10701 -2621 10753 -2567
rect 4801 -2655 4810 -2621
rect 4810 -2655 4848 -2621
rect 4848 -2655 4853 -2621
rect 5037 -2655 5064 -2621
rect 5064 -2655 5089 -2621
rect 5273 -2655 5280 -2621
rect 5280 -2655 5314 -2621
rect 5314 -2655 5325 -2621
rect 5509 -2655 5530 -2621
rect 5530 -2655 5561 -2621
rect 5745 -2655 5746 -2621
rect 5746 -2655 5784 -2621
rect 5784 -2655 5797 -2621
rect 5981 -2655 6000 -2621
rect 6000 -2655 6033 -2621
rect 6217 -2655 6250 -2621
rect 6250 -2655 6269 -2621
rect 6453 -2655 6466 -2621
rect 6466 -2655 6504 -2621
rect 6504 -2655 6505 -2621
rect 6689 -2655 6720 -2621
rect 6720 -2655 6741 -2621
rect 6925 -2655 6936 -2621
rect 6936 -2655 6970 -2621
rect 6970 -2655 6977 -2621
rect 7161 -2655 7186 -2621
rect 7186 -2655 7213 -2621
rect 7397 -2655 7402 -2621
rect 7402 -2655 7440 -2621
rect 7440 -2655 7449 -2621
rect 7633 -2655 7656 -2621
rect 7656 -2655 7685 -2621
rect 7869 -2655 7872 -2621
rect 7872 -2655 7906 -2621
rect 7906 -2655 7921 -2621
rect 8105 -2655 8122 -2621
rect 8122 -2655 8157 -2621
rect 8341 -2655 8376 -2621
rect 8376 -2655 8393 -2621
rect 8577 -2655 8592 -2621
rect 8592 -2655 8626 -2621
rect 8626 -2655 8629 -2621
rect 8813 -2655 8842 -2621
rect 8842 -2655 8865 -2621
rect 9049 -2655 9058 -2621
rect 9058 -2655 9096 -2621
rect 9096 -2655 9101 -2621
rect 9285 -2655 9312 -2621
rect 9312 -2655 9337 -2621
rect 9521 -2655 9528 -2621
rect 9528 -2655 9562 -2621
rect 9562 -2655 9573 -2621
rect 9757 -2655 9778 -2621
rect 9778 -2655 9809 -2621
rect 9993 -2655 9994 -2621
rect 9994 -2655 10032 -2621
rect 10032 -2655 10045 -2621
rect 10229 -2655 10248 -2621
rect 10248 -2655 10281 -2621
rect 10465 -2655 10498 -2621
rect 10498 -2655 10517 -2621
rect 10701 -2655 10714 -2621
rect 10714 -2655 10752 -2621
rect 10752 -2655 10753 -2621
rect 4801 -2675 4853 -2655
rect 5037 -2675 5089 -2655
rect 5273 -2675 5325 -2655
rect 5509 -2675 5561 -2655
rect 5745 -2675 5797 -2655
rect 5981 -2675 6033 -2655
rect 6217 -2675 6269 -2655
rect 6453 -2675 6505 -2655
rect 6689 -2675 6741 -2655
rect 6925 -2675 6977 -2655
rect 7161 -2675 7213 -2655
rect 7397 -2675 7449 -2655
rect 7633 -2675 7685 -2655
rect 7869 -2675 7921 -2655
rect 8105 -2675 8157 -2655
rect 8341 -2675 8393 -2655
rect 8577 -2675 8629 -2655
rect 8813 -2675 8865 -2655
rect 9049 -2675 9101 -2655
rect 9285 -2675 9337 -2655
rect 9521 -2675 9573 -2655
rect 9757 -2675 9809 -2655
rect 9993 -2675 10045 -2655
rect 10229 -2675 10281 -2655
rect 10465 -2675 10517 -2655
rect 10701 -2675 10753 -2655
rect 4801 -3490 4810 -2930
rect 4810 -3490 4844 -2930
rect 4844 -3490 4853 -2930
rect 4921 -3490 4928 -2930
rect 4928 -3490 4962 -2930
rect 4962 -3490 4973 -2930
rect 5037 -3490 5046 -2930
rect 5046 -3490 5080 -2930
rect 5080 -3490 5089 -2930
rect 5157 -3490 5164 -2930
rect 5164 -3490 5198 -2930
rect 5198 -3490 5209 -2930
rect 5273 -3490 5282 -2930
rect 5282 -3490 5316 -2930
rect 5316 -3490 5325 -2930
rect 5393 -3490 5400 -2930
rect 5400 -3490 5434 -2930
rect 5434 -3490 5445 -2930
rect 5509 -3490 5518 -2930
rect 5518 -3490 5552 -2930
rect 5552 -3490 5561 -2930
rect 5629 -3490 5636 -2930
rect 5636 -3490 5670 -2930
rect 5670 -3490 5681 -2930
rect 5745 -3490 5754 -2930
rect 5754 -3490 5788 -2930
rect 5788 -3490 5797 -2930
rect 5865 -3490 5872 -2930
rect 5872 -3490 5906 -2930
rect 5906 -3490 5917 -2930
rect 5981 -3490 5990 -2930
rect 5990 -3490 6024 -2930
rect 6024 -3490 6033 -2930
rect 6101 -3490 6108 -2930
rect 6108 -3490 6142 -2930
rect 6142 -3490 6153 -2930
rect 6217 -3490 6226 -2930
rect 6226 -3490 6260 -2930
rect 6260 -3490 6269 -2930
rect 6337 -3490 6344 -2930
rect 6344 -3490 6378 -2930
rect 6378 -3490 6389 -2930
rect 6453 -3490 6462 -2930
rect 6462 -3490 6496 -2930
rect 6496 -3490 6505 -2930
rect 6573 -3490 6580 -2930
rect 6580 -3490 6614 -2930
rect 6614 -3490 6625 -2930
rect 6689 -3490 6698 -2930
rect 6698 -3490 6732 -2930
rect 6732 -3490 6741 -2930
rect 6809 -3490 6816 -2930
rect 6816 -3490 6850 -2930
rect 6850 -3490 6861 -2930
rect 6925 -3490 6934 -2930
rect 6934 -3490 6968 -2930
rect 6968 -3490 6977 -2930
rect 7045 -3490 7052 -2930
rect 7052 -3490 7086 -2930
rect 7086 -3490 7097 -2930
rect 7161 -3490 7170 -2930
rect 7170 -3490 7204 -2930
rect 7204 -3490 7213 -2930
rect 7281 -3490 7288 -2930
rect 7288 -3490 7322 -2930
rect 7322 -3490 7333 -2930
rect 7397 -3490 7406 -2930
rect 7406 -3490 7440 -2930
rect 7440 -3490 7449 -2930
rect 7517 -3490 7524 -2930
rect 7524 -3490 7558 -2930
rect 7558 -3490 7569 -2930
rect 7633 -3490 7642 -2930
rect 7642 -3490 7676 -2930
rect 7676 -3490 7685 -2930
rect 7753 -3490 7760 -2930
rect 7760 -3490 7794 -2930
rect 7794 -3490 7805 -2930
rect 7869 -3490 7878 -2930
rect 7878 -3490 7912 -2930
rect 7912 -3490 7921 -2930
rect 7989 -3490 7996 -2930
rect 7996 -3490 8030 -2930
rect 8030 -3490 8041 -2930
rect 8105 -3490 8114 -2930
rect 8114 -3490 8148 -2930
rect 8148 -3490 8157 -2930
rect 8225 -3490 8232 -2930
rect 8232 -3490 8266 -2930
rect 8266 -3490 8277 -2930
rect 8341 -3490 8350 -2930
rect 8350 -3490 8384 -2930
rect 8384 -3490 8393 -2930
rect 8461 -3490 8468 -2930
rect 8468 -3490 8502 -2930
rect 8502 -3490 8513 -2930
rect 8577 -3490 8586 -2930
rect 8586 -3490 8620 -2930
rect 8620 -3490 8629 -2930
rect 8697 -3490 8704 -2930
rect 8704 -3490 8738 -2930
rect 8738 -3490 8749 -2930
rect 8813 -3490 8822 -2930
rect 8822 -3490 8856 -2930
rect 8856 -3490 8865 -2930
rect 8933 -3490 8940 -2930
rect 8940 -3490 8974 -2930
rect 8974 -3490 8985 -2930
rect 9049 -3490 9058 -2930
rect 9058 -3490 9092 -2930
rect 9092 -3490 9101 -2930
rect 9169 -3490 9176 -2930
rect 9176 -3490 9210 -2930
rect 9210 -3490 9221 -2930
rect 9285 -3490 9294 -2930
rect 9294 -3490 9328 -2930
rect 9328 -3490 9337 -2930
rect 9405 -3490 9412 -2930
rect 9412 -3490 9446 -2930
rect 9446 -3490 9457 -2930
rect 9521 -3490 9530 -2930
rect 9530 -3490 9564 -2930
rect 9564 -3490 9573 -2930
rect 9641 -3490 9648 -2930
rect 9648 -3490 9682 -2930
rect 9682 -3490 9693 -2930
rect 9757 -3490 9766 -2930
rect 9766 -3490 9800 -2930
rect 9800 -3490 9809 -2930
rect 9877 -3490 9884 -2930
rect 9884 -3490 9918 -2930
rect 9918 -3490 9929 -2930
rect 9993 -3490 10002 -2930
rect 10002 -3490 10036 -2930
rect 10036 -3490 10045 -2930
rect 10113 -3490 10120 -2930
rect 10120 -3490 10154 -2930
rect 10154 -3490 10165 -2930
rect 10229 -3490 10238 -2930
rect 10238 -3490 10272 -2930
rect 10272 -3490 10281 -2930
rect 10349 -3490 10356 -2930
rect 10356 -3490 10390 -2930
rect 10390 -3490 10401 -2930
rect 10465 -3490 10474 -2930
rect 10474 -3490 10508 -2930
rect 10508 -3490 10517 -2930
rect 10585 -3490 10592 -2930
rect 10592 -3490 10626 -2930
rect 10626 -3490 10637 -2930
rect 10701 -3490 10710 -2930
rect 10710 -3490 10744 -2930
rect 10744 -3490 10753 -2930
rect 4857 -3557 4915 -3551
rect 4857 -3591 4869 -3557
rect 4869 -3591 4903 -3557
rect 4903 -3591 4915 -3557
rect 4857 -3665 4915 -3591
rect 4857 -3699 4869 -3665
rect 4869 -3699 4903 -3665
rect 4903 -3699 4915 -3665
rect 4857 -3705 4915 -3699
rect 4975 -3557 5033 -3551
rect 4975 -3591 4987 -3557
rect 4987 -3591 5021 -3557
rect 5021 -3591 5033 -3557
rect 4975 -3665 5033 -3591
rect 4975 -3699 4987 -3665
rect 4987 -3699 5021 -3665
rect 5021 -3699 5033 -3665
rect 4975 -3705 5033 -3699
rect 5093 -3557 5151 -3551
rect 5093 -3591 5105 -3557
rect 5105 -3591 5139 -3557
rect 5139 -3591 5151 -3557
rect 5093 -3665 5151 -3591
rect 5093 -3699 5105 -3665
rect 5105 -3699 5139 -3665
rect 5139 -3699 5151 -3665
rect 5093 -3705 5151 -3699
rect 5211 -3557 5269 -3551
rect 5211 -3591 5223 -3557
rect 5223 -3591 5257 -3557
rect 5257 -3591 5269 -3557
rect 5211 -3665 5269 -3591
rect 5211 -3699 5223 -3665
rect 5223 -3699 5257 -3665
rect 5257 -3699 5269 -3665
rect 5211 -3705 5269 -3699
rect 5329 -3557 5387 -3551
rect 5329 -3591 5341 -3557
rect 5341 -3591 5375 -3557
rect 5375 -3591 5387 -3557
rect 5329 -3665 5387 -3591
rect 5329 -3699 5341 -3665
rect 5341 -3699 5375 -3665
rect 5375 -3699 5387 -3665
rect 5329 -3705 5387 -3699
rect 5447 -3557 5505 -3551
rect 5447 -3591 5459 -3557
rect 5459 -3591 5493 -3557
rect 5493 -3591 5505 -3557
rect 5447 -3665 5505 -3591
rect 5447 -3699 5459 -3665
rect 5459 -3699 5493 -3665
rect 5493 -3699 5505 -3665
rect 5447 -3705 5505 -3699
rect 5565 -3557 5623 -3551
rect 5565 -3591 5577 -3557
rect 5577 -3591 5611 -3557
rect 5611 -3591 5623 -3557
rect 5565 -3665 5623 -3591
rect 5565 -3699 5577 -3665
rect 5577 -3699 5611 -3665
rect 5611 -3699 5623 -3665
rect 5565 -3705 5623 -3699
rect 5683 -3557 5741 -3551
rect 5683 -3591 5695 -3557
rect 5695 -3591 5729 -3557
rect 5729 -3591 5741 -3557
rect 5683 -3665 5741 -3591
rect 5683 -3699 5695 -3665
rect 5695 -3699 5729 -3665
rect 5729 -3699 5741 -3665
rect 5683 -3705 5741 -3699
rect 5801 -3557 5859 -3551
rect 5801 -3591 5813 -3557
rect 5813 -3591 5847 -3557
rect 5847 -3591 5859 -3557
rect 5801 -3665 5859 -3591
rect 5801 -3699 5813 -3665
rect 5813 -3699 5847 -3665
rect 5847 -3699 5859 -3665
rect 5801 -3705 5859 -3699
rect 5919 -3557 5977 -3551
rect 5919 -3591 5931 -3557
rect 5931 -3591 5965 -3557
rect 5965 -3591 5977 -3557
rect 5919 -3665 5977 -3591
rect 5919 -3699 5931 -3665
rect 5931 -3699 5965 -3665
rect 5965 -3699 5977 -3665
rect 5919 -3705 5977 -3699
rect 6037 -3557 6095 -3551
rect 6037 -3591 6049 -3557
rect 6049 -3591 6083 -3557
rect 6083 -3591 6095 -3557
rect 6037 -3665 6095 -3591
rect 6037 -3699 6049 -3665
rect 6049 -3699 6083 -3665
rect 6083 -3699 6095 -3665
rect 6037 -3705 6095 -3699
rect 6155 -3557 6213 -3551
rect 6155 -3591 6167 -3557
rect 6167 -3591 6201 -3557
rect 6201 -3591 6213 -3557
rect 6155 -3665 6213 -3591
rect 6155 -3699 6167 -3665
rect 6167 -3699 6201 -3665
rect 6201 -3699 6213 -3665
rect 6155 -3705 6213 -3699
rect 6273 -3557 6331 -3551
rect 6273 -3591 6285 -3557
rect 6285 -3591 6319 -3557
rect 6319 -3591 6331 -3557
rect 6273 -3665 6331 -3591
rect 6273 -3699 6285 -3665
rect 6285 -3699 6319 -3665
rect 6319 -3699 6331 -3665
rect 6273 -3705 6331 -3699
rect 6391 -3557 6449 -3551
rect 6391 -3591 6403 -3557
rect 6403 -3591 6437 -3557
rect 6437 -3591 6449 -3557
rect 6391 -3665 6449 -3591
rect 6391 -3699 6403 -3665
rect 6403 -3699 6437 -3665
rect 6437 -3699 6449 -3665
rect 6391 -3705 6449 -3699
rect 6509 -3557 6567 -3551
rect 6509 -3591 6521 -3557
rect 6521 -3591 6555 -3557
rect 6555 -3591 6567 -3557
rect 6509 -3665 6567 -3591
rect 6509 -3699 6521 -3665
rect 6521 -3699 6555 -3665
rect 6555 -3699 6567 -3665
rect 6509 -3705 6567 -3699
rect 6627 -3557 6685 -3551
rect 6627 -3591 6639 -3557
rect 6639 -3591 6673 -3557
rect 6673 -3591 6685 -3557
rect 6627 -3665 6685 -3591
rect 6627 -3699 6639 -3665
rect 6639 -3699 6673 -3665
rect 6673 -3699 6685 -3665
rect 6627 -3705 6685 -3699
rect 6745 -3557 6803 -3551
rect 6745 -3591 6757 -3557
rect 6757 -3591 6791 -3557
rect 6791 -3591 6803 -3557
rect 6745 -3665 6803 -3591
rect 6745 -3699 6757 -3665
rect 6757 -3699 6791 -3665
rect 6791 -3699 6803 -3665
rect 6745 -3705 6803 -3699
rect 6863 -3557 6921 -3551
rect 6863 -3591 6875 -3557
rect 6875 -3591 6909 -3557
rect 6909 -3591 6921 -3557
rect 6863 -3665 6921 -3591
rect 6863 -3699 6875 -3665
rect 6875 -3699 6909 -3665
rect 6909 -3699 6921 -3665
rect 6863 -3705 6921 -3699
rect 6981 -3557 7039 -3551
rect 6981 -3591 6993 -3557
rect 6993 -3591 7027 -3557
rect 7027 -3591 7039 -3557
rect 6981 -3665 7039 -3591
rect 6981 -3699 6993 -3665
rect 6993 -3699 7027 -3665
rect 7027 -3699 7039 -3665
rect 6981 -3705 7039 -3699
rect 7099 -3557 7157 -3551
rect 7099 -3591 7111 -3557
rect 7111 -3591 7145 -3557
rect 7145 -3591 7157 -3557
rect 7099 -3665 7157 -3591
rect 7099 -3699 7111 -3665
rect 7111 -3699 7145 -3665
rect 7145 -3699 7157 -3665
rect 7099 -3705 7157 -3699
rect 7217 -3557 7275 -3551
rect 7217 -3591 7229 -3557
rect 7229 -3591 7263 -3557
rect 7263 -3591 7275 -3557
rect 7217 -3665 7275 -3591
rect 7217 -3699 7229 -3665
rect 7229 -3699 7263 -3665
rect 7263 -3699 7275 -3665
rect 7217 -3705 7275 -3699
rect 7335 -3557 7393 -3551
rect 7335 -3591 7347 -3557
rect 7347 -3591 7381 -3557
rect 7381 -3591 7393 -3557
rect 7335 -3665 7393 -3591
rect 7335 -3699 7347 -3665
rect 7347 -3699 7381 -3665
rect 7381 -3699 7393 -3665
rect 7335 -3705 7393 -3699
rect 7453 -3557 7511 -3551
rect 7453 -3591 7465 -3557
rect 7465 -3591 7499 -3557
rect 7499 -3591 7511 -3557
rect 7453 -3665 7511 -3591
rect 7453 -3699 7465 -3665
rect 7465 -3699 7499 -3665
rect 7499 -3699 7511 -3665
rect 7453 -3705 7511 -3699
rect 7571 -3557 7629 -3551
rect 7571 -3591 7583 -3557
rect 7583 -3591 7617 -3557
rect 7617 -3591 7629 -3557
rect 7571 -3665 7629 -3591
rect 7571 -3699 7583 -3665
rect 7583 -3699 7617 -3665
rect 7617 -3699 7629 -3665
rect 7571 -3705 7629 -3699
rect 7689 -3557 7747 -3551
rect 7689 -3591 7701 -3557
rect 7701 -3591 7735 -3557
rect 7735 -3591 7747 -3557
rect 7689 -3665 7747 -3591
rect 7689 -3699 7701 -3665
rect 7701 -3699 7735 -3665
rect 7735 -3699 7747 -3665
rect 7689 -3705 7747 -3699
rect 7807 -3557 7865 -3551
rect 7807 -3591 7819 -3557
rect 7819 -3591 7853 -3557
rect 7853 -3591 7865 -3557
rect 7807 -3665 7865 -3591
rect 7807 -3699 7819 -3665
rect 7819 -3699 7853 -3665
rect 7853 -3699 7865 -3665
rect 7807 -3705 7865 -3699
rect 7925 -3557 7983 -3551
rect 7925 -3591 7937 -3557
rect 7937 -3591 7971 -3557
rect 7971 -3591 7983 -3557
rect 7925 -3665 7983 -3591
rect 7925 -3699 7937 -3665
rect 7937 -3699 7971 -3665
rect 7971 -3699 7983 -3665
rect 7925 -3705 7983 -3699
rect 8043 -3557 8101 -3551
rect 8043 -3591 8055 -3557
rect 8055 -3591 8089 -3557
rect 8089 -3591 8101 -3557
rect 8043 -3665 8101 -3591
rect 8043 -3699 8055 -3665
rect 8055 -3699 8089 -3665
rect 8089 -3699 8101 -3665
rect 8043 -3705 8101 -3699
rect 8161 -3557 8219 -3551
rect 8161 -3591 8173 -3557
rect 8173 -3591 8207 -3557
rect 8207 -3591 8219 -3557
rect 8161 -3665 8219 -3591
rect 8161 -3699 8173 -3665
rect 8173 -3699 8207 -3665
rect 8207 -3699 8219 -3665
rect 8161 -3705 8219 -3699
rect 8279 -3557 8337 -3551
rect 8279 -3591 8291 -3557
rect 8291 -3591 8325 -3557
rect 8325 -3591 8337 -3557
rect 8279 -3665 8337 -3591
rect 8279 -3699 8291 -3665
rect 8291 -3699 8325 -3665
rect 8325 -3699 8337 -3665
rect 8279 -3705 8337 -3699
rect 8397 -3557 8455 -3551
rect 8397 -3591 8409 -3557
rect 8409 -3591 8443 -3557
rect 8443 -3591 8455 -3557
rect 8397 -3665 8455 -3591
rect 8397 -3699 8409 -3665
rect 8409 -3699 8443 -3665
rect 8443 -3699 8455 -3665
rect 8397 -3705 8455 -3699
rect 8515 -3557 8573 -3551
rect 8515 -3591 8527 -3557
rect 8527 -3591 8561 -3557
rect 8561 -3591 8573 -3557
rect 8515 -3665 8573 -3591
rect 8515 -3699 8527 -3665
rect 8527 -3699 8561 -3665
rect 8561 -3699 8573 -3665
rect 8515 -3705 8573 -3699
rect 8633 -3557 8691 -3551
rect 8633 -3591 8645 -3557
rect 8645 -3591 8679 -3557
rect 8679 -3591 8691 -3557
rect 8633 -3665 8691 -3591
rect 8633 -3699 8645 -3665
rect 8645 -3699 8679 -3665
rect 8679 -3699 8691 -3665
rect 8633 -3705 8691 -3699
rect 8751 -3557 8809 -3551
rect 8751 -3591 8763 -3557
rect 8763 -3591 8797 -3557
rect 8797 -3591 8809 -3557
rect 8751 -3665 8809 -3591
rect 8751 -3699 8763 -3665
rect 8763 -3699 8797 -3665
rect 8797 -3699 8809 -3665
rect 8751 -3705 8809 -3699
rect 8869 -3557 8927 -3551
rect 8869 -3591 8881 -3557
rect 8881 -3591 8915 -3557
rect 8915 -3591 8927 -3557
rect 8869 -3665 8927 -3591
rect 8869 -3699 8881 -3665
rect 8881 -3699 8915 -3665
rect 8915 -3699 8927 -3665
rect 8869 -3705 8927 -3699
rect 8987 -3557 9045 -3551
rect 8987 -3591 8999 -3557
rect 8999 -3591 9033 -3557
rect 9033 -3591 9045 -3557
rect 8987 -3665 9045 -3591
rect 8987 -3699 8999 -3665
rect 8999 -3699 9033 -3665
rect 9033 -3699 9045 -3665
rect 8987 -3705 9045 -3699
rect 9105 -3557 9163 -3551
rect 9105 -3591 9117 -3557
rect 9117 -3591 9151 -3557
rect 9151 -3591 9163 -3557
rect 9105 -3665 9163 -3591
rect 9105 -3699 9117 -3665
rect 9117 -3699 9151 -3665
rect 9151 -3699 9163 -3665
rect 9105 -3705 9163 -3699
rect 9223 -3557 9281 -3551
rect 9223 -3591 9235 -3557
rect 9235 -3591 9269 -3557
rect 9269 -3591 9281 -3557
rect 9223 -3665 9281 -3591
rect 9223 -3699 9235 -3665
rect 9235 -3699 9269 -3665
rect 9269 -3699 9281 -3665
rect 9223 -3705 9281 -3699
rect 9341 -3557 9399 -3551
rect 9341 -3591 9353 -3557
rect 9353 -3591 9387 -3557
rect 9387 -3591 9399 -3557
rect 9341 -3665 9399 -3591
rect 9341 -3699 9353 -3665
rect 9353 -3699 9387 -3665
rect 9387 -3699 9399 -3665
rect 9341 -3705 9399 -3699
rect 9459 -3557 9517 -3551
rect 9459 -3591 9471 -3557
rect 9471 -3591 9505 -3557
rect 9505 -3591 9517 -3557
rect 9459 -3665 9517 -3591
rect 9459 -3699 9471 -3665
rect 9471 -3699 9505 -3665
rect 9505 -3699 9517 -3665
rect 9459 -3705 9517 -3699
rect 9577 -3557 9635 -3551
rect 9577 -3591 9589 -3557
rect 9589 -3591 9623 -3557
rect 9623 -3591 9635 -3557
rect 9577 -3665 9635 -3591
rect 9577 -3699 9589 -3665
rect 9589 -3699 9623 -3665
rect 9623 -3699 9635 -3665
rect 9577 -3705 9635 -3699
rect 9695 -3557 9753 -3551
rect 9695 -3591 9707 -3557
rect 9707 -3591 9741 -3557
rect 9741 -3591 9753 -3557
rect 9695 -3665 9753 -3591
rect 9695 -3699 9707 -3665
rect 9707 -3699 9741 -3665
rect 9741 -3699 9753 -3665
rect 9695 -3705 9753 -3699
rect 9813 -3557 9871 -3551
rect 9813 -3591 9825 -3557
rect 9825 -3591 9859 -3557
rect 9859 -3591 9871 -3557
rect 9813 -3665 9871 -3591
rect 9813 -3699 9825 -3665
rect 9825 -3699 9859 -3665
rect 9859 -3699 9871 -3665
rect 9813 -3705 9871 -3699
rect 9931 -3557 9989 -3551
rect 9931 -3591 9943 -3557
rect 9943 -3591 9977 -3557
rect 9977 -3591 9989 -3557
rect 9931 -3665 9989 -3591
rect 9931 -3699 9943 -3665
rect 9943 -3699 9977 -3665
rect 9977 -3699 9989 -3665
rect 9931 -3705 9989 -3699
rect 10049 -3557 10107 -3551
rect 10049 -3591 10061 -3557
rect 10061 -3591 10095 -3557
rect 10095 -3591 10107 -3557
rect 10049 -3665 10107 -3591
rect 10049 -3699 10061 -3665
rect 10061 -3699 10095 -3665
rect 10095 -3699 10107 -3665
rect 10049 -3705 10107 -3699
rect 10167 -3557 10225 -3551
rect 10167 -3591 10179 -3557
rect 10179 -3591 10213 -3557
rect 10213 -3591 10225 -3557
rect 10167 -3665 10225 -3591
rect 10167 -3699 10179 -3665
rect 10179 -3699 10213 -3665
rect 10213 -3699 10225 -3665
rect 10167 -3705 10225 -3699
rect 10285 -3557 10343 -3551
rect 10285 -3591 10297 -3557
rect 10297 -3591 10331 -3557
rect 10331 -3591 10343 -3557
rect 10285 -3665 10343 -3591
rect 10285 -3699 10297 -3665
rect 10297 -3699 10331 -3665
rect 10331 -3699 10343 -3665
rect 10285 -3705 10343 -3699
rect 10403 -3557 10461 -3551
rect 10403 -3591 10415 -3557
rect 10415 -3591 10449 -3557
rect 10449 -3591 10461 -3557
rect 10403 -3665 10461 -3591
rect 10403 -3699 10415 -3665
rect 10415 -3699 10449 -3665
rect 10449 -3699 10461 -3665
rect 10403 -3705 10461 -3699
rect 10521 -3557 10579 -3551
rect 10521 -3591 10533 -3557
rect 10533 -3591 10567 -3557
rect 10567 -3591 10579 -3557
rect 10521 -3665 10579 -3591
rect 10521 -3699 10533 -3665
rect 10533 -3699 10567 -3665
rect 10567 -3699 10579 -3665
rect 10521 -3705 10579 -3699
rect 10639 -3557 10697 -3551
rect 10639 -3591 10651 -3557
rect 10651 -3591 10685 -3557
rect 10685 -3591 10697 -3557
rect 10639 -3665 10697 -3591
rect 10639 -3699 10651 -3665
rect 10651 -3699 10685 -3665
rect 10685 -3699 10697 -3665
rect 10639 -3705 10697 -3699
rect 4801 -4326 4810 -3766
rect 4810 -4326 4844 -3766
rect 4844 -4326 4853 -3766
rect 4921 -4326 4928 -3766
rect 4928 -4326 4962 -3766
rect 4962 -4326 4973 -3766
rect 5037 -4326 5046 -3766
rect 5046 -4326 5080 -3766
rect 5080 -4326 5089 -3766
rect 5157 -4326 5164 -3766
rect 5164 -4326 5198 -3766
rect 5198 -4326 5209 -3766
rect 5273 -4326 5282 -3766
rect 5282 -4326 5316 -3766
rect 5316 -4326 5325 -3766
rect 5393 -4326 5400 -3766
rect 5400 -4326 5434 -3766
rect 5434 -4326 5445 -3766
rect 5509 -4326 5518 -3766
rect 5518 -4326 5552 -3766
rect 5552 -4326 5561 -3766
rect 5629 -4326 5636 -3766
rect 5636 -4326 5670 -3766
rect 5670 -4326 5681 -3766
rect 5745 -4326 5754 -3766
rect 5754 -4326 5788 -3766
rect 5788 -4326 5797 -3766
rect 5865 -4326 5872 -3766
rect 5872 -4326 5906 -3766
rect 5906 -4326 5917 -3766
rect 5981 -4326 5990 -3766
rect 5990 -4326 6024 -3766
rect 6024 -4326 6033 -3766
rect 6101 -4326 6108 -3766
rect 6108 -4326 6142 -3766
rect 6142 -4326 6153 -3766
rect 6217 -4326 6226 -3766
rect 6226 -4326 6260 -3766
rect 6260 -4326 6269 -3766
rect 6337 -4326 6344 -3766
rect 6344 -4326 6378 -3766
rect 6378 -4326 6389 -3766
rect 6453 -4326 6462 -3766
rect 6462 -4326 6496 -3766
rect 6496 -4326 6505 -3766
rect 6573 -4326 6580 -3766
rect 6580 -4326 6614 -3766
rect 6614 -4326 6625 -3766
rect 6689 -4326 6698 -3766
rect 6698 -4326 6732 -3766
rect 6732 -4326 6741 -3766
rect 6809 -4326 6816 -3766
rect 6816 -4326 6850 -3766
rect 6850 -4326 6861 -3766
rect 6925 -4326 6934 -3766
rect 6934 -4326 6968 -3766
rect 6968 -4326 6977 -3766
rect 7045 -4326 7052 -3766
rect 7052 -4326 7086 -3766
rect 7086 -4326 7097 -3766
rect 7161 -4326 7170 -3766
rect 7170 -4326 7204 -3766
rect 7204 -4326 7213 -3766
rect 7281 -4326 7288 -3766
rect 7288 -4326 7322 -3766
rect 7322 -4326 7333 -3766
rect 7397 -4326 7406 -3766
rect 7406 -4326 7440 -3766
rect 7440 -4326 7449 -3766
rect 7517 -4326 7524 -3766
rect 7524 -4326 7558 -3766
rect 7558 -4326 7569 -3766
rect 7633 -4326 7642 -3766
rect 7642 -4326 7676 -3766
rect 7676 -4326 7685 -3766
rect 7753 -4326 7760 -3766
rect 7760 -4326 7794 -3766
rect 7794 -4326 7805 -3766
rect 7869 -4326 7878 -3766
rect 7878 -4326 7912 -3766
rect 7912 -4326 7921 -3766
rect 7989 -4326 7996 -3766
rect 7996 -4326 8030 -3766
rect 8030 -4326 8041 -3766
rect 8105 -4326 8114 -3766
rect 8114 -4326 8148 -3766
rect 8148 -4326 8157 -3766
rect 8225 -4326 8232 -3766
rect 8232 -4326 8266 -3766
rect 8266 -4326 8277 -3766
rect 8341 -4326 8350 -3766
rect 8350 -4326 8384 -3766
rect 8384 -4326 8393 -3766
rect 8461 -4326 8468 -3766
rect 8468 -4326 8502 -3766
rect 8502 -4326 8513 -3766
rect 8577 -4326 8586 -3766
rect 8586 -4326 8620 -3766
rect 8620 -4326 8629 -3766
rect 8697 -4326 8704 -3766
rect 8704 -4326 8738 -3766
rect 8738 -4326 8749 -3766
rect 8813 -4326 8822 -3766
rect 8822 -4326 8856 -3766
rect 8856 -4326 8865 -3766
rect 8933 -4326 8940 -3766
rect 8940 -4326 8974 -3766
rect 8974 -4326 8985 -3766
rect 9049 -4326 9058 -3766
rect 9058 -4326 9092 -3766
rect 9092 -4326 9101 -3766
rect 9169 -4326 9176 -3766
rect 9176 -4326 9210 -3766
rect 9210 -4326 9221 -3766
rect 9285 -4326 9294 -3766
rect 9294 -4326 9328 -3766
rect 9328 -4326 9337 -3766
rect 9405 -4326 9412 -3766
rect 9412 -4326 9446 -3766
rect 9446 -4326 9457 -3766
rect 9521 -4326 9530 -3766
rect 9530 -4326 9564 -3766
rect 9564 -4326 9573 -3766
rect 9641 -4326 9648 -3766
rect 9648 -4326 9682 -3766
rect 9682 -4326 9693 -3766
rect 9757 -4326 9766 -3766
rect 9766 -4326 9800 -3766
rect 9800 -4326 9809 -3766
rect 9877 -4326 9884 -3766
rect 9884 -4326 9918 -3766
rect 9918 -4326 9929 -3766
rect 9993 -4326 10002 -3766
rect 10002 -4326 10036 -3766
rect 10036 -4326 10045 -3766
rect 10113 -4326 10120 -3766
rect 10120 -4326 10154 -3766
rect 10154 -4326 10165 -3766
rect 10229 -4326 10238 -3766
rect 10238 -4326 10272 -3766
rect 10272 -4326 10281 -3766
rect 10349 -4326 10356 -3766
rect 10356 -4326 10390 -3766
rect 10390 -4326 10401 -3766
rect 10465 -4326 10474 -3766
rect 10474 -4326 10508 -3766
rect 10508 -4326 10517 -3766
rect 10585 -4326 10592 -3766
rect 10592 -4326 10626 -3766
rect 10626 -4326 10637 -3766
rect 10701 -4326 10710 -3766
rect 10710 -4326 10744 -3766
rect 10744 -4326 10753 -3766
rect 4801 -4495 4853 -4475
rect 5037 -4495 5089 -4475
rect 5273 -4495 5325 -4475
rect 5509 -4495 5561 -4475
rect 5745 -4495 5797 -4475
rect 5981 -4495 6033 -4475
rect 6217 -4495 6269 -4475
rect 6453 -4495 6505 -4475
rect 6689 -4495 6741 -4475
rect 6925 -4495 6977 -4475
rect 7161 -4495 7213 -4475
rect 7397 -4495 7449 -4475
rect 7633 -4495 7685 -4475
rect 7869 -4495 7921 -4475
rect 8105 -4495 8157 -4475
rect 8341 -4495 8393 -4475
rect 8577 -4495 8629 -4475
rect 8813 -4495 8865 -4475
rect 9049 -4495 9101 -4475
rect 9285 -4495 9337 -4475
rect 9521 -4495 9573 -4475
rect 9757 -4495 9809 -4475
rect 9993 -4495 10045 -4475
rect 10229 -4495 10281 -4475
rect 10465 -4495 10517 -4475
rect 10701 -4495 10753 -4475
rect 4801 -4529 4802 -4495
rect 4802 -4529 4840 -4495
rect 4840 -4529 4853 -4495
rect 5037 -4529 5056 -4495
rect 5056 -4529 5089 -4495
rect 5273 -4529 5306 -4495
rect 5306 -4529 5325 -4495
rect 5509 -4529 5522 -4495
rect 5522 -4529 5560 -4495
rect 5560 -4529 5561 -4495
rect 5745 -4529 5776 -4495
rect 5776 -4529 5797 -4495
rect 5981 -4529 5992 -4495
rect 5992 -4529 6026 -4495
rect 6026 -4529 6033 -4495
rect 6217 -4529 6242 -4495
rect 6242 -4529 6269 -4495
rect 6453 -4529 6458 -4495
rect 6458 -4529 6496 -4495
rect 6496 -4529 6505 -4495
rect 6689 -4529 6712 -4495
rect 6712 -4529 6741 -4495
rect 6925 -4529 6928 -4495
rect 6928 -4529 6962 -4495
rect 6962 -4529 6977 -4495
rect 7161 -4529 7178 -4495
rect 7178 -4529 7213 -4495
rect 7397 -4529 7432 -4495
rect 7432 -4529 7449 -4495
rect 7633 -4529 7648 -4495
rect 7648 -4529 7682 -4495
rect 7682 -4529 7685 -4495
rect 7869 -4529 7898 -4495
rect 7898 -4529 7921 -4495
rect 8105 -4529 8114 -4495
rect 8114 -4529 8152 -4495
rect 8152 -4529 8157 -4495
rect 8341 -4529 8368 -4495
rect 8368 -4529 8393 -4495
rect 8577 -4529 8584 -4495
rect 8584 -4529 8618 -4495
rect 8618 -4529 8629 -4495
rect 8813 -4529 8834 -4495
rect 8834 -4529 8865 -4495
rect 9049 -4529 9050 -4495
rect 9050 -4529 9088 -4495
rect 9088 -4529 9101 -4495
rect 9285 -4529 9304 -4495
rect 9304 -4529 9337 -4495
rect 9521 -4529 9554 -4495
rect 9554 -4529 9573 -4495
rect 9757 -4529 9770 -4495
rect 9770 -4529 9808 -4495
rect 9808 -4529 9809 -4495
rect 9993 -4529 10024 -4495
rect 10024 -4529 10045 -4495
rect 10229 -4529 10240 -4495
rect 10240 -4529 10274 -4495
rect 10274 -4529 10281 -4495
rect 10465 -4529 10490 -4495
rect 10490 -4529 10517 -4495
rect 10701 -4529 10706 -4495
rect 10706 -4529 10744 -4495
rect 10744 -4529 10753 -4495
rect 4801 -4583 4853 -4529
rect 5037 -4583 5089 -4529
rect 5273 -4583 5325 -4529
rect 5509 -4583 5561 -4529
rect 5745 -4583 5797 -4529
rect 5981 -4583 6033 -4529
rect 6217 -4583 6269 -4529
rect 6453 -4583 6505 -4529
rect 6689 -4583 6741 -4529
rect 6925 -4583 6977 -4529
rect 7161 -4583 7213 -4529
rect 7397 -4583 7449 -4529
rect 7633 -4583 7685 -4529
rect 7869 -4583 7921 -4529
rect 8105 -4583 8157 -4529
rect 8341 -4583 8393 -4529
rect 8577 -4583 8629 -4529
rect 8813 -4583 8865 -4529
rect 9049 -4583 9101 -4529
rect 9285 -4583 9337 -4529
rect 9521 -4583 9573 -4529
rect 9757 -4583 9809 -4529
rect 9993 -4583 10045 -4529
rect 10229 -4583 10281 -4529
rect 10465 -4583 10517 -4529
rect 10701 -4583 10753 -4529
rect 4801 -4617 4802 -4583
rect 4802 -4617 4840 -4583
rect 4840 -4617 4853 -4583
rect 5037 -4617 5056 -4583
rect 5056 -4617 5089 -4583
rect 5273 -4617 5306 -4583
rect 5306 -4617 5325 -4583
rect 5509 -4617 5522 -4583
rect 5522 -4617 5560 -4583
rect 5560 -4617 5561 -4583
rect 5745 -4617 5776 -4583
rect 5776 -4617 5797 -4583
rect 5981 -4617 5992 -4583
rect 5992 -4617 6026 -4583
rect 6026 -4617 6033 -4583
rect 6217 -4617 6242 -4583
rect 6242 -4617 6269 -4583
rect 6453 -4617 6458 -4583
rect 6458 -4617 6496 -4583
rect 6496 -4617 6505 -4583
rect 6689 -4617 6712 -4583
rect 6712 -4617 6741 -4583
rect 6925 -4617 6928 -4583
rect 6928 -4617 6962 -4583
rect 6962 -4617 6977 -4583
rect 7161 -4617 7178 -4583
rect 7178 -4617 7213 -4583
rect 7397 -4617 7432 -4583
rect 7432 -4617 7449 -4583
rect 7633 -4617 7648 -4583
rect 7648 -4617 7682 -4583
rect 7682 -4617 7685 -4583
rect 7869 -4617 7898 -4583
rect 7898 -4617 7921 -4583
rect 8105 -4617 8114 -4583
rect 8114 -4617 8152 -4583
rect 8152 -4617 8157 -4583
rect 8341 -4617 8368 -4583
rect 8368 -4617 8393 -4583
rect 8577 -4617 8584 -4583
rect 8584 -4617 8618 -4583
rect 8618 -4617 8629 -4583
rect 8813 -4617 8834 -4583
rect 8834 -4617 8865 -4583
rect 9049 -4617 9050 -4583
rect 9050 -4617 9088 -4583
rect 9088 -4617 9101 -4583
rect 9285 -4617 9304 -4583
rect 9304 -4617 9337 -4583
rect 9521 -4617 9554 -4583
rect 9554 -4617 9573 -4583
rect 9757 -4617 9770 -4583
rect 9770 -4617 9808 -4583
rect 9808 -4617 9809 -4583
rect 9993 -4617 10024 -4583
rect 10024 -4617 10045 -4583
rect 10229 -4617 10240 -4583
rect 10240 -4617 10274 -4583
rect 10274 -4617 10281 -4583
rect 10465 -4617 10490 -4583
rect 10490 -4617 10517 -4583
rect 10701 -4617 10706 -4583
rect 10706 -4617 10744 -4583
rect 10744 -4617 10753 -4583
rect 4801 -4671 4853 -4617
rect 5037 -4671 5089 -4617
rect 5273 -4671 5325 -4617
rect 5509 -4671 5561 -4617
rect 5745 -4671 5797 -4617
rect 5981 -4671 6033 -4617
rect 6217 -4671 6269 -4617
rect 6453 -4671 6505 -4617
rect 6689 -4671 6741 -4617
rect 6925 -4671 6977 -4617
rect 7161 -4671 7213 -4617
rect 7397 -4671 7449 -4617
rect 7633 -4671 7685 -4617
rect 7869 -4671 7921 -4617
rect 8105 -4671 8157 -4617
rect 8341 -4671 8393 -4617
rect 8577 -4671 8629 -4617
rect 8813 -4671 8865 -4617
rect 9049 -4671 9101 -4617
rect 9285 -4671 9337 -4617
rect 9521 -4671 9573 -4617
rect 9757 -4671 9809 -4617
rect 9993 -4671 10045 -4617
rect 10229 -4671 10281 -4617
rect 10465 -4671 10517 -4617
rect 10701 -4671 10753 -4617
rect 4801 -4705 4802 -4671
rect 4802 -4705 4840 -4671
rect 4840 -4705 4853 -4671
rect 5037 -4705 5056 -4671
rect 5056 -4705 5089 -4671
rect 5273 -4705 5306 -4671
rect 5306 -4705 5325 -4671
rect 5509 -4705 5522 -4671
rect 5522 -4705 5560 -4671
rect 5560 -4705 5561 -4671
rect 5745 -4705 5776 -4671
rect 5776 -4705 5797 -4671
rect 5981 -4705 5992 -4671
rect 5992 -4705 6026 -4671
rect 6026 -4705 6033 -4671
rect 6217 -4705 6242 -4671
rect 6242 -4705 6269 -4671
rect 6453 -4705 6458 -4671
rect 6458 -4705 6496 -4671
rect 6496 -4705 6505 -4671
rect 6689 -4705 6712 -4671
rect 6712 -4705 6741 -4671
rect 6925 -4705 6928 -4671
rect 6928 -4705 6962 -4671
rect 6962 -4705 6977 -4671
rect 7161 -4705 7178 -4671
rect 7178 -4705 7213 -4671
rect 7397 -4705 7432 -4671
rect 7432 -4705 7449 -4671
rect 7633 -4705 7648 -4671
rect 7648 -4705 7682 -4671
rect 7682 -4705 7685 -4671
rect 7869 -4705 7898 -4671
rect 7898 -4705 7921 -4671
rect 8105 -4705 8114 -4671
rect 8114 -4705 8152 -4671
rect 8152 -4705 8157 -4671
rect 8341 -4705 8368 -4671
rect 8368 -4705 8393 -4671
rect 8577 -4705 8584 -4671
rect 8584 -4705 8618 -4671
rect 8618 -4705 8629 -4671
rect 8813 -4705 8834 -4671
rect 8834 -4705 8865 -4671
rect 9049 -4705 9050 -4671
rect 9050 -4705 9088 -4671
rect 9088 -4705 9101 -4671
rect 9285 -4705 9304 -4671
rect 9304 -4705 9337 -4671
rect 9521 -4705 9554 -4671
rect 9554 -4705 9573 -4671
rect 9757 -4705 9770 -4671
rect 9770 -4705 9808 -4671
rect 9808 -4705 9809 -4671
rect 9993 -4705 10024 -4671
rect 10024 -4705 10045 -4671
rect 10229 -4705 10240 -4671
rect 10240 -4705 10274 -4671
rect 10274 -4705 10281 -4671
rect 10465 -4705 10490 -4671
rect 10490 -4705 10517 -4671
rect 10701 -4705 10706 -4671
rect 10706 -4705 10744 -4671
rect 10744 -4705 10753 -4671
rect 4801 -4725 4853 -4705
rect 5037 -4725 5089 -4705
rect 5273 -4725 5325 -4705
rect 5509 -4725 5561 -4705
rect 5745 -4725 5797 -4705
rect 5981 -4725 6033 -4705
rect 6217 -4725 6269 -4705
rect 6453 -4725 6505 -4705
rect 6689 -4725 6741 -4705
rect 6925 -4725 6977 -4705
rect 7161 -4725 7213 -4705
rect 7397 -4725 7449 -4705
rect 7633 -4725 7685 -4705
rect 7869 -4725 7921 -4705
rect 8105 -4725 8157 -4705
rect 8341 -4725 8393 -4705
rect 8577 -4725 8629 -4705
rect 8813 -4725 8865 -4705
rect 9049 -4725 9101 -4705
rect 9285 -4725 9337 -4705
rect 9521 -4725 9573 -4705
rect 9757 -4725 9809 -4705
rect 9993 -4725 10045 -4705
rect 10229 -4725 10281 -4705
rect 10465 -4725 10517 -4705
rect 10701 -4725 10753 -4705
rect 4801 -5540 4853 -4980
rect 4921 -5540 4973 -4980
rect 5037 -5540 5046 -4980
rect 5046 -5540 5080 -4980
rect 5080 -5540 5089 -4980
rect 5157 -5540 5164 -4980
rect 5164 -5540 5198 -4980
rect 5198 -5540 5209 -4980
rect 5273 -5540 5282 -4980
rect 5282 -5540 5316 -4980
rect 5316 -5540 5325 -4980
rect 5393 -5540 5400 -4980
rect 5400 -5540 5434 -4980
rect 5434 -5540 5445 -4980
rect 5509 -5540 5518 -4980
rect 5518 -5540 5552 -4980
rect 5552 -5540 5561 -4980
rect 5629 -5540 5636 -4980
rect 5636 -5540 5670 -4980
rect 5670 -5540 5681 -4980
rect 5745 -5540 5754 -4980
rect 5754 -5540 5788 -4980
rect 5788 -5540 5797 -4980
rect 5865 -5540 5872 -4980
rect 5872 -5540 5906 -4980
rect 5906 -5540 5917 -4980
rect 5981 -5540 5990 -4980
rect 5990 -5540 6024 -4980
rect 6024 -5540 6033 -4980
rect 6101 -5540 6108 -4980
rect 6108 -5540 6142 -4980
rect 6142 -5540 6153 -4980
rect 6217 -5540 6226 -4980
rect 6226 -5540 6260 -4980
rect 6260 -5540 6269 -4980
rect 6337 -5540 6344 -4980
rect 6344 -5540 6378 -4980
rect 6378 -5540 6389 -4980
rect 6453 -5540 6462 -4980
rect 6462 -5540 6496 -4980
rect 6496 -5540 6505 -4980
rect 6573 -5540 6580 -4980
rect 6580 -5540 6614 -4980
rect 6614 -5540 6625 -4980
rect 6689 -5540 6698 -4980
rect 6698 -5540 6732 -4980
rect 6732 -5540 6741 -4980
rect 6809 -5540 6816 -4980
rect 6816 -5540 6850 -4980
rect 6850 -5540 6861 -4980
rect 6925 -5540 6934 -4980
rect 6934 -5540 6968 -4980
rect 6968 -5540 6977 -4980
rect 7045 -5540 7052 -4980
rect 7052 -5540 7086 -4980
rect 7086 -5540 7097 -4980
rect 7161 -5540 7170 -4980
rect 7170 -5540 7204 -4980
rect 7204 -5540 7213 -4980
rect 7281 -5540 7288 -4980
rect 7288 -5540 7322 -4980
rect 7322 -5540 7333 -4980
rect 7397 -5540 7406 -4980
rect 7406 -5540 7440 -4980
rect 7440 -5540 7449 -4980
rect 7517 -5540 7524 -4980
rect 7524 -5540 7558 -4980
rect 7558 -5540 7569 -4980
rect 7633 -5540 7642 -4980
rect 7642 -5540 7676 -4980
rect 7676 -5540 7685 -4980
rect 7753 -5540 7760 -4980
rect 7760 -5540 7794 -4980
rect 7794 -5540 7805 -4980
rect 7869 -5540 7878 -4980
rect 7878 -5540 7912 -4980
rect 7912 -5540 7921 -4980
rect 7989 -5540 7996 -4980
rect 7996 -5540 8030 -4980
rect 8030 -5540 8041 -4980
rect 8105 -5540 8114 -4980
rect 8114 -5540 8148 -4980
rect 8148 -5540 8157 -4980
rect 8225 -5540 8232 -4980
rect 8232 -5540 8266 -4980
rect 8266 -5540 8277 -4980
rect 8341 -5540 8350 -4980
rect 8350 -5540 8384 -4980
rect 8384 -5540 8393 -4980
rect 8461 -5540 8468 -4980
rect 8468 -5540 8502 -4980
rect 8502 -5540 8513 -4980
rect 8577 -5540 8586 -4980
rect 8586 -5540 8620 -4980
rect 8620 -5540 8629 -4980
rect 8697 -5540 8704 -4980
rect 8704 -5540 8738 -4980
rect 8738 -5540 8749 -4980
rect 8813 -5540 8822 -4980
rect 8822 -5540 8856 -4980
rect 8856 -5540 8865 -4980
rect 8933 -5540 8940 -4980
rect 8940 -5540 8974 -4980
rect 8974 -5540 8985 -4980
rect 9049 -5540 9058 -4980
rect 9058 -5540 9092 -4980
rect 9092 -5540 9101 -4980
rect 9169 -5540 9176 -4980
rect 9176 -5540 9210 -4980
rect 9210 -5540 9221 -4980
rect 9285 -5540 9294 -4980
rect 9294 -5540 9328 -4980
rect 9328 -5540 9337 -4980
rect 9405 -5540 9412 -4980
rect 9412 -5540 9446 -4980
rect 9446 -5540 9457 -4980
rect 9521 -5540 9530 -4980
rect 9530 -5540 9564 -4980
rect 9564 -5540 9573 -4980
rect 9641 -5540 9648 -4980
rect 9648 -5540 9682 -4980
rect 9682 -5540 9693 -4980
rect 9757 -5540 9766 -4980
rect 9766 -5540 9800 -4980
rect 9800 -5540 9809 -4980
rect 9877 -5540 9884 -4980
rect 9884 -5540 9918 -4980
rect 9918 -5540 9929 -4980
rect 9993 -5540 10002 -4980
rect 10002 -5540 10036 -4980
rect 10036 -5540 10045 -4980
rect 10113 -5540 10120 -4980
rect 10120 -5540 10154 -4980
rect 10154 -5540 10165 -4980
rect 10229 -5540 10238 -4980
rect 10238 -5540 10272 -4980
rect 10272 -5540 10281 -4980
rect 10349 -5540 10356 -4980
rect 10356 -5540 10390 -4980
rect 10390 -5540 10401 -4980
rect 10465 -5540 10474 -4980
rect 10474 -5540 10508 -4980
rect 10508 -5540 10517 -4980
rect 10585 -5540 10592 -4980
rect 10592 -5540 10626 -4980
rect 10626 -5540 10637 -4980
rect 10701 -5540 10710 -4980
rect 10710 -5540 10744 -4980
rect 10744 -5540 10753 -4980
rect 4857 -5607 4915 -5601
rect 4857 -5641 4869 -5607
rect 4869 -5641 4903 -5607
rect 4903 -5641 4915 -5607
rect 4857 -5715 4915 -5641
rect 4857 -5749 4869 -5715
rect 4869 -5749 4903 -5715
rect 4903 -5749 4915 -5715
rect 4857 -5755 4915 -5749
rect 4975 -5607 5033 -5601
rect 4975 -5641 4987 -5607
rect 4987 -5641 5021 -5607
rect 5021 -5641 5033 -5607
rect 4975 -5715 5033 -5641
rect 4975 -5749 4987 -5715
rect 4987 -5749 5021 -5715
rect 5021 -5749 5033 -5715
rect 4975 -5755 5033 -5749
rect 5093 -5607 5151 -5601
rect 5093 -5641 5105 -5607
rect 5105 -5641 5139 -5607
rect 5139 -5641 5151 -5607
rect 5093 -5715 5151 -5641
rect 5093 -5749 5105 -5715
rect 5105 -5749 5139 -5715
rect 5139 -5749 5151 -5715
rect 5093 -5755 5151 -5749
rect 5211 -5607 5269 -5601
rect 5211 -5641 5223 -5607
rect 5223 -5641 5257 -5607
rect 5257 -5641 5269 -5607
rect 5211 -5715 5269 -5641
rect 5211 -5749 5223 -5715
rect 5223 -5749 5257 -5715
rect 5257 -5749 5269 -5715
rect 5211 -5755 5269 -5749
rect 5329 -5607 5387 -5601
rect 5329 -5641 5341 -5607
rect 5341 -5641 5375 -5607
rect 5375 -5641 5387 -5607
rect 5329 -5715 5387 -5641
rect 5329 -5749 5341 -5715
rect 5341 -5749 5375 -5715
rect 5375 -5749 5387 -5715
rect 5329 -5755 5387 -5749
rect 5447 -5607 5505 -5601
rect 5447 -5641 5459 -5607
rect 5459 -5641 5493 -5607
rect 5493 -5641 5505 -5607
rect 5447 -5715 5505 -5641
rect 5447 -5749 5459 -5715
rect 5459 -5749 5493 -5715
rect 5493 -5749 5505 -5715
rect 5447 -5755 5505 -5749
rect 5565 -5607 5623 -5601
rect 5565 -5641 5577 -5607
rect 5577 -5641 5611 -5607
rect 5611 -5641 5623 -5607
rect 5565 -5715 5623 -5641
rect 5565 -5749 5577 -5715
rect 5577 -5749 5611 -5715
rect 5611 -5749 5623 -5715
rect 5565 -5755 5623 -5749
rect 5683 -5607 5741 -5601
rect 5683 -5641 5695 -5607
rect 5695 -5641 5729 -5607
rect 5729 -5641 5741 -5607
rect 5683 -5715 5741 -5641
rect 5683 -5749 5695 -5715
rect 5695 -5749 5729 -5715
rect 5729 -5749 5741 -5715
rect 5683 -5755 5741 -5749
rect 5801 -5607 5859 -5601
rect 5801 -5641 5813 -5607
rect 5813 -5641 5847 -5607
rect 5847 -5641 5859 -5607
rect 5801 -5715 5859 -5641
rect 5801 -5749 5813 -5715
rect 5813 -5749 5847 -5715
rect 5847 -5749 5859 -5715
rect 5801 -5755 5859 -5749
rect 5919 -5607 5977 -5601
rect 5919 -5641 5931 -5607
rect 5931 -5641 5965 -5607
rect 5965 -5641 5977 -5607
rect 5919 -5715 5977 -5641
rect 5919 -5749 5931 -5715
rect 5931 -5749 5965 -5715
rect 5965 -5749 5977 -5715
rect 5919 -5755 5977 -5749
rect 6037 -5607 6095 -5601
rect 6037 -5641 6049 -5607
rect 6049 -5641 6083 -5607
rect 6083 -5641 6095 -5607
rect 6037 -5715 6095 -5641
rect 6037 -5749 6049 -5715
rect 6049 -5749 6083 -5715
rect 6083 -5749 6095 -5715
rect 6037 -5755 6095 -5749
rect 6155 -5607 6213 -5601
rect 6155 -5641 6167 -5607
rect 6167 -5641 6201 -5607
rect 6201 -5641 6213 -5607
rect 6155 -5715 6213 -5641
rect 6155 -5749 6167 -5715
rect 6167 -5749 6201 -5715
rect 6201 -5749 6213 -5715
rect 6155 -5755 6213 -5749
rect 6273 -5607 6331 -5601
rect 6273 -5641 6285 -5607
rect 6285 -5641 6319 -5607
rect 6319 -5641 6331 -5607
rect 6273 -5715 6331 -5641
rect 6273 -5749 6285 -5715
rect 6285 -5749 6319 -5715
rect 6319 -5749 6331 -5715
rect 6273 -5755 6331 -5749
rect 6391 -5607 6449 -5601
rect 6391 -5641 6403 -5607
rect 6403 -5641 6437 -5607
rect 6437 -5641 6449 -5607
rect 6391 -5715 6449 -5641
rect 6391 -5749 6403 -5715
rect 6403 -5749 6437 -5715
rect 6437 -5749 6449 -5715
rect 6391 -5755 6449 -5749
rect 6509 -5607 6567 -5601
rect 6509 -5641 6521 -5607
rect 6521 -5641 6555 -5607
rect 6555 -5641 6567 -5607
rect 6509 -5715 6567 -5641
rect 6509 -5749 6521 -5715
rect 6521 -5749 6555 -5715
rect 6555 -5749 6567 -5715
rect 6509 -5755 6567 -5749
rect 6627 -5607 6685 -5601
rect 6627 -5641 6639 -5607
rect 6639 -5641 6673 -5607
rect 6673 -5641 6685 -5607
rect 6627 -5715 6685 -5641
rect 6627 -5749 6639 -5715
rect 6639 -5749 6673 -5715
rect 6673 -5749 6685 -5715
rect 6627 -5755 6685 -5749
rect 6745 -5607 6803 -5601
rect 6745 -5641 6757 -5607
rect 6757 -5641 6791 -5607
rect 6791 -5641 6803 -5607
rect 6745 -5715 6803 -5641
rect 6745 -5749 6757 -5715
rect 6757 -5749 6791 -5715
rect 6791 -5749 6803 -5715
rect 6745 -5755 6803 -5749
rect 6863 -5607 6921 -5601
rect 6863 -5641 6875 -5607
rect 6875 -5641 6909 -5607
rect 6909 -5641 6921 -5607
rect 6863 -5715 6921 -5641
rect 6863 -5749 6875 -5715
rect 6875 -5749 6909 -5715
rect 6909 -5749 6921 -5715
rect 6863 -5755 6921 -5749
rect 6981 -5607 7039 -5601
rect 6981 -5641 6993 -5607
rect 6993 -5641 7027 -5607
rect 7027 -5641 7039 -5607
rect 6981 -5715 7039 -5641
rect 6981 -5749 6993 -5715
rect 6993 -5749 7027 -5715
rect 7027 -5749 7039 -5715
rect 6981 -5755 7039 -5749
rect 7099 -5607 7157 -5601
rect 7099 -5641 7111 -5607
rect 7111 -5641 7145 -5607
rect 7145 -5641 7157 -5607
rect 7099 -5715 7157 -5641
rect 7099 -5749 7111 -5715
rect 7111 -5749 7145 -5715
rect 7145 -5749 7157 -5715
rect 7099 -5755 7157 -5749
rect 7217 -5607 7275 -5601
rect 7217 -5641 7229 -5607
rect 7229 -5641 7263 -5607
rect 7263 -5641 7275 -5607
rect 7217 -5715 7275 -5641
rect 7217 -5749 7229 -5715
rect 7229 -5749 7263 -5715
rect 7263 -5749 7275 -5715
rect 7217 -5755 7275 -5749
rect 7335 -5607 7393 -5601
rect 7335 -5641 7347 -5607
rect 7347 -5641 7381 -5607
rect 7381 -5641 7393 -5607
rect 7335 -5715 7393 -5641
rect 7335 -5749 7347 -5715
rect 7347 -5749 7381 -5715
rect 7381 -5749 7393 -5715
rect 7335 -5755 7393 -5749
rect 7453 -5607 7511 -5601
rect 7453 -5641 7465 -5607
rect 7465 -5641 7499 -5607
rect 7499 -5641 7511 -5607
rect 7453 -5715 7511 -5641
rect 7453 -5749 7465 -5715
rect 7465 -5749 7499 -5715
rect 7499 -5749 7511 -5715
rect 7453 -5755 7511 -5749
rect 7571 -5607 7629 -5601
rect 7571 -5641 7583 -5607
rect 7583 -5641 7617 -5607
rect 7617 -5641 7629 -5607
rect 7571 -5715 7629 -5641
rect 7571 -5749 7583 -5715
rect 7583 -5749 7617 -5715
rect 7617 -5749 7629 -5715
rect 7571 -5755 7629 -5749
rect 7689 -5607 7747 -5601
rect 7689 -5641 7701 -5607
rect 7701 -5641 7735 -5607
rect 7735 -5641 7747 -5607
rect 7689 -5715 7747 -5641
rect 7689 -5749 7701 -5715
rect 7701 -5749 7735 -5715
rect 7735 -5749 7747 -5715
rect 7689 -5755 7747 -5749
rect 7807 -5607 7865 -5601
rect 7807 -5641 7819 -5607
rect 7819 -5641 7853 -5607
rect 7853 -5641 7865 -5607
rect 7807 -5715 7865 -5641
rect 7807 -5749 7819 -5715
rect 7819 -5749 7853 -5715
rect 7853 -5749 7865 -5715
rect 7807 -5755 7865 -5749
rect 7925 -5607 7983 -5601
rect 7925 -5641 7937 -5607
rect 7937 -5641 7971 -5607
rect 7971 -5641 7983 -5607
rect 7925 -5715 7983 -5641
rect 7925 -5749 7937 -5715
rect 7937 -5749 7971 -5715
rect 7971 -5749 7983 -5715
rect 7925 -5755 7983 -5749
rect 8043 -5607 8101 -5601
rect 8043 -5641 8055 -5607
rect 8055 -5641 8089 -5607
rect 8089 -5641 8101 -5607
rect 8043 -5715 8101 -5641
rect 8043 -5749 8055 -5715
rect 8055 -5749 8089 -5715
rect 8089 -5749 8101 -5715
rect 8043 -5755 8101 -5749
rect 8161 -5607 8219 -5601
rect 8161 -5641 8173 -5607
rect 8173 -5641 8207 -5607
rect 8207 -5641 8219 -5607
rect 8161 -5715 8219 -5641
rect 8161 -5749 8173 -5715
rect 8173 -5749 8207 -5715
rect 8207 -5749 8219 -5715
rect 8161 -5755 8219 -5749
rect 8279 -5607 8337 -5601
rect 8279 -5641 8291 -5607
rect 8291 -5641 8325 -5607
rect 8325 -5641 8337 -5607
rect 8279 -5715 8337 -5641
rect 8279 -5749 8291 -5715
rect 8291 -5749 8325 -5715
rect 8325 -5749 8337 -5715
rect 8279 -5755 8337 -5749
rect 8397 -5607 8455 -5601
rect 8397 -5641 8409 -5607
rect 8409 -5641 8443 -5607
rect 8443 -5641 8455 -5607
rect 8397 -5715 8455 -5641
rect 8397 -5749 8409 -5715
rect 8409 -5749 8443 -5715
rect 8443 -5749 8455 -5715
rect 8397 -5755 8455 -5749
rect 8515 -5607 8573 -5601
rect 8515 -5641 8527 -5607
rect 8527 -5641 8561 -5607
rect 8561 -5641 8573 -5607
rect 8515 -5715 8573 -5641
rect 8515 -5749 8527 -5715
rect 8527 -5749 8561 -5715
rect 8561 -5749 8573 -5715
rect 8515 -5755 8573 -5749
rect 8633 -5607 8691 -5601
rect 8633 -5641 8645 -5607
rect 8645 -5641 8679 -5607
rect 8679 -5641 8691 -5607
rect 8633 -5715 8691 -5641
rect 8633 -5749 8645 -5715
rect 8645 -5749 8679 -5715
rect 8679 -5749 8691 -5715
rect 8633 -5755 8691 -5749
rect 8751 -5607 8809 -5601
rect 8751 -5641 8763 -5607
rect 8763 -5641 8797 -5607
rect 8797 -5641 8809 -5607
rect 8751 -5715 8809 -5641
rect 8751 -5749 8763 -5715
rect 8763 -5749 8797 -5715
rect 8797 -5749 8809 -5715
rect 8751 -5755 8809 -5749
rect 8869 -5607 8927 -5601
rect 8869 -5641 8881 -5607
rect 8881 -5641 8915 -5607
rect 8915 -5641 8927 -5607
rect 8869 -5715 8927 -5641
rect 8869 -5749 8881 -5715
rect 8881 -5749 8915 -5715
rect 8915 -5749 8927 -5715
rect 8869 -5755 8927 -5749
rect 8987 -5607 9045 -5601
rect 8987 -5641 8999 -5607
rect 8999 -5641 9033 -5607
rect 9033 -5641 9045 -5607
rect 8987 -5715 9045 -5641
rect 8987 -5749 8999 -5715
rect 8999 -5749 9033 -5715
rect 9033 -5749 9045 -5715
rect 8987 -5755 9045 -5749
rect 9105 -5607 9163 -5601
rect 9105 -5641 9117 -5607
rect 9117 -5641 9151 -5607
rect 9151 -5641 9163 -5607
rect 9105 -5715 9163 -5641
rect 9105 -5749 9117 -5715
rect 9117 -5749 9151 -5715
rect 9151 -5749 9163 -5715
rect 9105 -5755 9163 -5749
rect 9223 -5607 9281 -5601
rect 9223 -5641 9235 -5607
rect 9235 -5641 9269 -5607
rect 9269 -5641 9281 -5607
rect 9223 -5715 9281 -5641
rect 9223 -5749 9235 -5715
rect 9235 -5749 9269 -5715
rect 9269 -5749 9281 -5715
rect 9223 -5755 9281 -5749
rect 9341 -5607 9399 -5601
rect 9341 -5641 9353 -5607
rect 9353 -5641 9387 -5607
rect 9387 -5641 9399 -5607
rect 9341 -5715 9399 -5641
rect 9341 -5749 9353 -5715
rect 9353 -5749 9387 -5715
rect 9387 -5749 9399 -5715
rect 9341 -5755 9399 -5749
rect 9459 -5607 9517 -5601
rect 9459 -5641 9471 -5607
rect 9471 -5641 9505 -5607
rect 9505 -5641 9517 -5607
rect 9459 -5715 9517 -5641
rect 9459 -5749 9471 -5715
rect 9471 -5749 9505 -5715
rect 9505 -5749 9517 -5715
rect 9459 -5755 9517 -5749
rect 9577 -5607 9635 -5601
rect 9577 -5641 9589 -5607
rect 9589 -5641 9623 -5607
rect 9623 -5641 9635 -5607
rect 9577 -5715 9635 -5641
rect 9577 -5749 9589 -5715
rect 9589 -5749 9623 -5715
rect 9623 -5749 9635 -5715
rect 9577 -5755 9635 -5749
rect 9695 -5607 9753 -5601
rect 9695 -5641 9707 -5607
rect 9707 -5641 9741 -5607
rect 9741 -5641 9753 -5607
rect 9695 -5715 9753 -5641
rect 9695 -5749 9707 -5715
rect 9707 -5749 9741 -5715
rect 9741 -5749 9753 -5715
rect 9695 -5755 9753 -5749
rect 9813 -5607 9871 -5601
rect 9813 -5641 9825 -5607
rect 9825 -5641 9859 -5607
rect 9859 -5641 9871 -5607
rect 9813 -5715 9871 -5641
rect 9813 -5749 9825 -5715
rect 9825 -5749 9859 -5715
rect 9859 -5749 9871 -5715
rect 9813 -5755 9871 -5749
rect 9931 -5607 9989 -5601
rect 9931 -5641 9943 -5607
rect 9943 -5641 9977 -5607
rect 9977 -5641 9989 -5607
rect 9931 -5715 9989 -5641
rect 9931 -5749 9943 -5715
rect 9943 -5749 9977 -5715
rect 9977 -5749 9989 -5715
rect 9931 -5755 9989 -5749
rect 10049 -5607 10107 -5601
rect 10049 -5641 10061 -5607
rect 10061 -5641 10095 -5607
rect 10095 -5641 10107 -5607
rect 10049 -5715 10107 -5641
rect 10049 -5749 10061 -5715
rect 10061 -5749 10095 -5715
rect 10095 -5749 10107 -5715
rect 10049 -5755 10107 -5749
rect 10167 -5607 10225 -5601
rect 10167 -5641 10179 -5607
rect 10179 -5641 10213 -5607
rect 10213 -5641 10225 -5607
rect 10167 -5715 10225 -5641
rect 10167 -5749 10179 -5715
rect 10179 -5749 10213 -5715
rect 10213 -5749 10225 -5715
rect 10167 -5755 10225 -5749
rect 10285 -5607 10343 -5601
rect 10285 -5641 10297 -5607
rect 10297 -5641 10331 -5607
rect 10331 -5641 10343 -5607
rect 10285 -5715 10343 -5641
rect 10285 -5749 10297 -5715
rect 10297 -5749 10331 -5715
rect 10331 -5749 10343 -5715
rect 10285 -5755 10343 -5749
rect 10403 -5607 10461 -5601
rect 10403 -5641 10415 -5607
rect 10415 -5641 10449 -5607
rect 10449 -5641 10461 -5607
rect 10403 -5715 10461 -5641
rect 10403 -5749 10415 -5715
rect 10415 -5749 10449 -5715
rect 10449 -5749 10461 -5715
rect 10403 -5755 10461 -5749
rect 10521 -5607 10579 -5601
rect 10521 -5641 10533 -5607
rect 10533 -5641 10567 -5607
rect 10567 -5641 10579 -5607
rect 10521 -5715 10579 -5641
rect 10521 -5749 10533 -5715
rect 10533 -5749 10567 -5715
rect 10567 -5749 10579 -5715
rect 10521 -5755 10579 -5749
rect 10639 -5607 10697 -5601
rect 10639 -5641 10651 -5607
rect 10651 -5641 10685 -5607
rect 10685 -5641 10697 -5607
rect 10639 -5715 10697 -5641
rect 10639 -5749 10651 -5715
rect 10651 -5749 10685 -5715
rect 10685 -5749 10697 -5715
rect 10639 -5755 10697 -5749
rect 4801 -6376 4810 -5816
rect 4810 -6376 4844 -5816
rect 4844 -6376 4853 -5816
rect 4921 -6376 4928 -5816
rect 4928 -6376 4962 -5816
rect 4962 -6376 4973 -5816
rect 5037 -6376 5046 -5816
rect 5046 -6376 5080 -5816
rect 5080 -6376 5089 -5816
rect 5157 -6376 5164 -5816
rect 5164 -6376 5198 -5816
rect 5198 -6376 5209 -5816
rect 5273 -6376 5282 -5816
rect 5282 -6376 5316 -5816
rect 5316 -6376 5325 -5816
rect 5393 -6376 5400 -5816
rect 5400 -6376 5434 -5816
rect 5434 -6376 5445 -5816
rect 5509 -6376 5518 -5816
rect 5518 -6376 5552 -5816
rect 5552 -6376 5561 -5816
rect 5629 -6376 5636 -5816
rect 5636 -6376 5670 -5816
rect 5670 -6376 5681 -5816
rect 5745 -6376 5754 -5816
rect 5754 -6376 5788 -5816
rect 5788 -6376 5797 -5816
rect 5865 -6376 5872 -5816
rect 5872 -6376 5906 -5816
rect 5906 -6376 5917 -5816
rect 5981 -6376 5990 -5816
rect 5990 -6376 6024 -5816
rect 6024 -6376 6033 -5816
rect 6101 -6376 6108 -5816
rect 6108 -6376 6142 -5816
rect 6142 -6376 6153 -5816
rect 6217 -6376 6226 -5816
rect 6226 -6376 6260 -5816
rect 6260 -6376 6269 -5816
rect 6337 -6376 6344 -5816
rect 6344 -6376 6378 -5816
rect 6378 -6376 6389 -5816
rect 6453 -6376 6462 -5816
rect 6462 -6376 6496 -5816
rect 6496 -6376 6505 -5816
rect 6573 -6376 6580 -5816
rect 6580 -6376 6614 -5816
rect 6614 -6376 6625 -5816
rect 6689 -6376 6698 -5816
rect 6698 -6376 6732 -5816
rect 6732 -6376 6741 -5816
rect 6809 -6376 6816 -5816
rect 6816 -6376 6850 -5816
rect 6850 -6376 6861 -5816
rect 6925 -6376 6934 -5816
rect 6934 -6376 6968 -5816
rect 6968 -6376 6977 -5816
rect 7045 -6376 7052 -5816
rect 7052 -6376 7086 -5816
rect 7086 -6376 7097 -5816
rect 7161 -6376 7170 -5816
rect 7170 -6376 7204 -5816
rect 7204 -6376 7213 -5816
rect 7281 -6376 7288 -5816
rect 7288 -6376 7322 -5816
rect 7322 -6376 7333 -5816
rect 7397 -6376 7406 -5816
rect 7406 -6376 7440 -5816
rect 7440 -6376 7449 -5816
rect 7517 -6376 7524 -5816
rect 7524 -6376 7558 -5816
rect 7558 -6376 7569 -5816
rect 7633 -6376 7642 -5816
rect 7642 -6376 7676 -5816
rect 7676 -6376 7685 -5816
rect 7753 -6376 7760 -5816
rect 7760 -6376 7794 -5816
rect 7794 -6376 7805 -5816
rect 7869 -6376 7878 -5816
rect 7878 -6376 7912 -5816
rect 7912 -6376 7921 -5816
rect 7989 -6376 7996 -5816
rect 7996 -6376 8030 -5816
rect 8030 -6376 8041 -5816
rect 8105 -6376 8114 -5816
rect 8114 -6376 8148 -5816
rect 8148 -6376 8157 -5816
rect 8225 -6376 8232 -5816
rect 8232 -6376 8266 -5816
rect 8266 -6376 8277 -5816
rect 8341 -6376 8350 -5816
rect 8350 -6376 8384 -5816
rect 8384 -6376 8393 -5816
rect 8461 -6376 8468 -5816
rect 8468 -6376 8502 -5816
rect 8502 -6376 8513 -5816
rect 8577 -6376 8586 -5816
rect 8586 -6376 8620 -5816
rect 8620 -6376 8629 -5816
rect 8697 -6376 8704 -5816
rect 8704 -6376 8738 -5816
rect 8738 -6376 8749 -5816
rect 8813 -6376 8822 -5816
rect 8822 -6376 8856 -5816
rect 8856 -6376 8865 -5816
rect 8933 -6376 8940 -5816
rect 8940 -6376 8974 -5816
rect 8974 -6376 8985 -5816
rect 9049 -6376 9058 -5816
rect 9058 -6376 9092 -5816
rect 9092 -6376 9101 -5816
rect 9169 -6376 9176 -5816
rect 9176 -6376 9210 -5816
rect 9210 -6376 9221 -5816
rect 9285 -6376 9294 -5816
rect 9294 -6376 9328 -5816
rect 9328 -6376 9337 -5816
rect 9405 -6376 9412 -5816
rect 9412 -6376 9446 -5816
rect 9446 -6376 9457 -5816
rect 9521 -6376 9530 -5816
rect 9530 -6376 9564 -5816
rect 9564 -6376 9573 -5816
rect 9641 -6376 9648 -5816
rect 9648 -6376 9682 -5816
rect 9682 -6376 9693 -5816
rect 9757 -6376 9766 -5816
rect 9766 -6376 9800 -5816
rect 9800 -6376 9809 -5816
rect 9877 -6376 9884 -5816
rect 9884 -6376 9918 -5816
rect 9918 -6376 9929 -5816
rect 9993 -6376 10002 -5816
rect 10002 -6376 10036 -5816
rect 10036 -6376 10045 -5816
rect 10113 -6376 10120 -5816
rect 10120 -6376 10154 -5816
rect 10154 -6376 10165 -5816
rect 10229 -6376 10238 -5816
rect 10238 -6376 10272 -5816
rect 10272 -6376 10281 -5816
rect 10349 -6376 10356 -5816
rect 10356 -6376 10390 -5816
rect 10390 -6376 10401 -5816
rect 10465 -6376 10474 -5816
rect 10474 -6376 10508 -5816
rect 10508 -6376 10517 -5816
rect 10585 -6376 10592 -5816
rect 10592 -6376 10626 -5816
rect 10626 -6376 10637 -5816
rect 10701 -6376 10710 -5816
rect 10710 -6376 10744 -5816
rect 10744 -6376 10753 -5816
rect 4801 -6775 4853 -6525
rect 5037 -6775 5089 -6525
rect 5273 -6775 5325 -6525
rect 5509 -6775 5561 -6525
rect 5745 -6775 5797 -6525
rect 5981 -6775 6033 -6525
rect 6217 -6775 6269 -6525
rect 6453 -6775 6505 -6525
rect 6689 -6775 6741 -6525
rect 6925 -6775 6977 -6525
rect 7161 -6775 7213 -6525
rect 7397 -6775 7449 -6525
rect 7633 -6775 7685 -6525
rect 7869 -6775 7921 -6525
rect 8105 -6775 8157 -6525
rect 8341 -6775 8393 -6525
rect 8577 -6775 8629 -6525
rect 8813 -6775 8865 -6525
rect 9049 -6775 9101 -6525
rect 9285 -6775 9337 -6525
rect 9521 -6775 9573 -6525
rect 9757 -6775 9809 -6525
rect 9993 -6775 10045 -6525
rect 10229 -6775 10281 -6525
rect 10465 -6775 10517 -6525
rect 10701 -6775 10753 -6525
rect 11068 -6752 11120 -6700
rect 11149 -6752 11201 -6700
rect 11230 -6752 11282 -6700
rect 11311 -6752 11363 -6700
rect 11392 -6752 11444 -6700
rect 11473 -6752 11525 -6700
rect 11554 -6752 11606 -6700
rect 11068 -6856 11120 -6804
rect 11149 -6856 11201 -6804
rect 11230 -6856 11282 -6804
rect 11311 -6856 11363 -6804
rect 11392 -6856 11444 -6804
rect 11473 -6856 11525 -6804
rect 11554 -6856 11606 -6804
rect 5759 -6994 5811 -6942
rect 5839 -6994 5891 -6942
rect 5919 -6994 5971 -6942
rect 5999 -6994 6051 -6942
rect 6079 -6994 6131 -6942
rect 6159 -6994 6211 -6942
rect 6239 -6994 6291 -6942
rect 6319 -6994 6371 -6942
rect 6399 -6994 6451 -6942
rect 6479 -6994 6531 -6942
rect 6559 -6994 6611 -6942
rect 6639 -6994 6691 -6942
rect 6719 -6994 6771 -6942
rect 6799 -6994 6851 -6942
rect 6879 -6994 6931 -6942
rect 6959 -6994 7011 -6942
rect 7039 -6994 7091 -6942
rect 7119 -6994 7171 -6942
rect 7199 -6994 7251 -6942
rect 7279 -6994 7331 -6942
rect 7359 -6994 7411 -6942
rect 7439 -6994 7491 -6942
rect 7519 -6994 7571 -6942
rect 7599 -6994 7651 -6942
rect 7679 -6994 7731 -6942
rect 7759 -6994 7811 -6942
rect 7839 -6994 7891 -6942
rect 7919 -6994 7971 -6942
rect 7999 -6994 8051 -6942
rect 8079 -6994 8131 -6942
rect 8159 -6994 8211 -6942
rect 8239 -6994 8291 -6942
rect 8319 -6994 8371 -6942
rect 8399 -6994 8451 -6942
rect 8479 -6994 8531 -6942
rect 8559 -6994 8611 -6942
rect 8639 -6994 8691 -6942
rect 8719 -6994 8771 -6942
rect 8799 -6994 8851 -6942
rect 8879 -6994 8931 -6942
rect 8959 -6994 9011 -6942
rect 9039 -6994 9091 -6942
rect 9119 -6994 9171 -6942
rect 9199 -6994 9251 -6942
rect 9279 -6994 9331 -6942
rect 9359 -6994 9411 -6942
rect 9439 -6994 9491 -6942
rect 9519 -6994 9571 -6942
rect 9599 -6994 9651 -6942
rect 9679 -6994 9731 -6942
rect 9759 -6994 9811 -6942
rect 9839 -6994 9891 -6942
rect 9919 -6994 9971 -6942
rect 9999 -6994 10051 -6942
rect 10079 -6994 10131 -6942
rect 10159 -6994 10211 -6942
rect 10239 -6994 10291 -6942
rect 10319 -6994 10371 -6942
rect 10399 -6994 10451 -6942
rect 10479 -6994 10531 -6942
rect 10559 -6994 10611 -6942
rect 10639 -6994 10691 -6942
rect 10719 -6994 10771 -6942
rect 10799 -6994 10851 -6942
rect 11068 -6960 11120 -6908
rect 11149 -6960 11201 -6908
rect 11230 -6960 11282 -6908
rect 11311 -6960 11363 -6908
rect 11392 -6960 11444 -6908
rect 11473 -6960 11525 -6908
rect 11554 -6960 11606 -6908
rect 4094 -7115 4146 -7063
rect 4175 -7115 4227 -7063
rect 4256 -7115 4308 -7063
rect 4337 -7115 4389 -7063
rect 4418 -7115 4470 -7063
rect 4499 -7115 4551 -7063
rect 4580 -7115 4632 -7063
rect 4662 -7115 4714 -7063
rect 4743 -7115 4795 -7063
rect 4824 -7115 4876 -7063
rect 4905 -7115 4957 -7063
rect 4986 -7115 5038 -7063
rect 5067 -7115 5119 -7063
rect 5148 -7115 5200 -7063
rect 5230 -7115 5282 -7063
rect 5311 -7115 5363 -7063
rect 5392 -7115 5444 -7063
rect 5759 -7074 5811 -7022
rect 5839 -7074 5891 -7022
rect 5919 -7074 5971 -7022
rect 5999 -7074 6051 -7022
rect 6079 -7074 6131 -7022
rect 6159 -7074 6211 -7022
rect 6239 -7074 6291 -7022
rect 6319 -7074 6371 -7022
rect 6399 -7074 6451 -7022
rect 6479 -7074 6531 -7022
rect 6559 -7074 6611 -7022
rect 6639 -7074 6691 -7022
rect 6719 -7074 6771 -7022
rect 6799 -7074 6851 -7022
rect 6879 -7074 6931 -7022
rect 6959 -7074 7011 -7022
rect 7039 -7074 7091 -7022
rect 7119 -7074 7171 -7022
rect 7199 -7074 7251 -7022
rect 7279 -7074 7331 -7022
rect 7359 -7074 7411 -7022
rect 7439 -7074 7491 -7022
rect 7519 -7074 7571 -7022
rect 7599 -7074 7651 -7022
rect 7679 -7074 7731 -7022
rect 7759 -7074 7811 -7022
rect 7839 -7074 7891 -7022
rect 7919 -7074 7971 -7022
rect 7999 -7074 8051 -7022
rect 8079 -7074 8131 -7022
rect 8159 -7074 8211 -7022
rect 8239 -7074 8291 -7022
rect 8319 -7074 8371 -7022
rect 8399 -7074 8451 -7022
rect 8479 -7074 8531 -7022
rect 8559 -7074 8611 -7022
rect 8639 -7074 8691 -7022
rect 8719 -7074 8771 -7022
rect 8799 -7074 8851 -7022
rect 8879 -7074 8931 -7022
rect 8959 -7074 9011 -7022
rect 9039 -7074 9091 -7022
rect 9119 -7074 9171 -7022
rect 9199 -7074 9251 -7022
rect 9279 -7074 9331 -7022
rect 9359 -7074 9411 -7022
rect 9439 -7074 9491 -7022
rect 9519 -7074 9571 -7022
rect 9599 -7074 9651 -7022
rect 9679 -7074 9731 -7022
rect 9759 -7074 9811 -7022
rect 9839 -7074 9891 -7022
rect 9919 -7074 9971 -7022
rect 9999 -7074 10051 -7022
rect 10079 -7074 10131 -7022
rect 10159 -7074 10211 -7022
rect 10239 -7074 10291 -7022
rect 10319 -7074 10371 -7022
rect 10399 -7074 10451 -7022
rect 10479 -7074 10531 -7022
rect 10559 -7074 10611 -7022
rect 10639 -7074 10691 -7022
rect 10719 -7074 10771 -7022
rect 10799 -7074 10851 -7022
rect 4094 -7199 4146 -7167
rect 4175 -7199 4227 -7167
rect 4256 -7199 4308 -7167
rect 4337 -7199 4389 -7167
rect 4418 -7199 4470 -7167
rect 4499 -7199 4551 -7167
rect 4580 -7199 4632 -7167
rect 4662 -7199 4714 -7167
rect 4094 -7219 4098 -7199
rect 4098 -7219 4132 -7199
rect 4132 -7219 4146 -7199
rect 4175 -7219 4204 -7199
rect 4204 -7219 4227 -7199
rect 4256 -7219 4276 -7199
rect 4276 -7219 4308 -7199
rect 4337 -7219 4348 -7199
rect 4348 -7219 4386 -7199
rect 4386 -7219 4389 -7199
rect 4418 -7219 4420 -7199
rect 4420 -7219 4458 -7199
rect 4458 -7219 4470 -7199
rect 4499 -7219 4530 -7199
rect 4530 -7219 4551 -7199
rect 4580 -7219 4602 -7199
rect 4602 -7219 4632 -7199
rect 4662 -7219 4674 -7199
rect 4674 -7219 4708 -7199
rect 4708 -7219 4714 -7199
rect 4743 -7199 4795 -7167
rect 4824 -7199 4876 -7167
rect 4905 -7199 4957 -7167
rect 4986 -7199 5038 -7167
rect 5067 -7199 5119 -7167
rect 5148 -7199 5200 -7167
rect 5230 -7199 5282 -7167
rect 5311 -7199 5363 -7167
rect 4743 -7219 4746 -7199
rect 4746 -7219 4780 -7199
rect 4780 -7219 4795 -7199
rect 4824 -7219 4852 -7199
rect 4852 -7219 4876 -7199
rect 4905 -7219 4924 -7199
rect 4924 -7219 4957 -7199
rect 4986 -7219 4996 -7199
rect 4996 -7219 5034 -7199
rect 5034 -7219 5038 -7199
rect 5067 -7219 5068 -7199
rect 5068 -7219 5106 -7199
rect 5106 -7219 5119 -7199
rect 5148 -7219 5178 -7199
rect 5178 -7219 5200 -7199
rect 5230 -7219 5250 -7199
rect 5250 -7219 5282 -7199
rect 5311 -7219 5322 -7199
rect 5322 -7219 5356 -7199
rect 5356 -7219 5363 -7199
rect 5392 -7199 5444 -7167
rect 5392 -7219 5394 -7199
rect 5394 -7219 5428 -7199
rect 5428 -7219 5444 -7199
rect 9839 -7223 9868 -7206
rect 9868 -7223 9891 -7206
rect 9919 -7223 9940 -7206
rect 9940 -7223 9971 -7206
rect 9999 -7223 10012 -7206
rect 10012 -7223 10050 -7206
rect 10050 -7223 10051 -7206
rect 10079 -7223 10084 -7206
rect 10084 -7223 10122 -7206
rect 10122 -7223 10131 -7206
rect 10159 -7223 10194 -7206
rect 10194 -7223 10211 -7206
rect 10239 -7223 10266 -7206
rect 10266 -7223 10291 -7206
rect 4094 -7273 4146 -7271
rect 4175 -7273 4227 -7271
rect 4256 -7273 4308 -7271
rect 4337 -7273 4389 -7271
rect 4418 -7273 4470 -7271
rect 4499 -7273 4551 -7271
rect 4580 -7273 4632 -7271
rect 4662 -7273 4714 -7271
rect 4094 -7307 4098 -7273
rect 4098 -7307 4132 -7273
rect 4132 -7307 4146 -7273
rect 4175 -7307 4204 -7273
rect 4204 -7307 4227 -7273
rect 4256 -7307 4276 -7273
rect 4276 -7307 4308 -7273
rect 4337 -7307 4348 -7273
rect 4348 -7307 4386 -7273
rect 4386 -7307 4389 -7273
rect 4418 -7307 4420 -7273
rect 4420 -7307 4458 -7273
rect 4458 -7307 4470 -7273
rect 4499 -7307 4530 -7273
rect 4530 -7307 4551 -7273
rect 4580 -7307 4602 -7273
rect 4602 -7307 4632 -7273
rect 4662 -7307 4674 -7273
rect 4674 -7307 4708 -7273
rect 4708 -7307 4714 -7273
rect 4094 -7323 4146 -7307
rect 4175 -7323 4227 -7307
rect 4256 -7323 4308 -7307
rect 4337 -7323 4389 -7307
rect 4418 -7323 4470 -7307
rect 4499 -7323 4551 -7307
rect 4580 -7323 4632 -7307
rect 4662 -7323 4714 -7307
rect 4743 -7273 4795 -7271
rect 4824 -7273 4876 -7271
rect 4905 -7273 4957 -7271
rect 4986 -7273 5038 -7271
rect 5067 -7273 5119 -7271
rect 5148 -7273 5200 -7271
rect 5230 -7273 5282 -7271
rect 5311 -7273 5363 -7271
rect 4743 -7307 4746 -7273
rect 4746 -7307 4780 -7273
rect 4780 -7307 4795 -7273
rect 4824 -7307 4852 -7273
rect 4852 -7307 4876 -7273
rect 4905 -7307 4924 -7273
rect 4924 -7307 4957 -7273
rect 4986 -7307 4996 -7273
rect 4996 -7307 5034 -7273
rect 5034 -7307 5038 -7273
rect 5067 -7307 5068 -7273
rect 5068 -7307 5106 -7273
rect 5106 -7307 5119 -7273
rect 5148 -7307 5178 -7273
rect 5178 -7307 5200 -7273
rect 5230 -7307 5250 -7273
rect 5250 -7307 5282 -7273
rect 5311 -7307 5322 -7273
rect 5322 -7307 5356 -7273
rect 5356 -7307 5363 -7273
rect 4743 -7323 4795 -7307
rect 4824 -7323 4876 -7307
rect 4905 -7323 4957 -7307
rect 4986 -7323 5038 -7307
rect 5067 -7323 5119 -7307
rect 5148 -7323 5200 -7307
rect 5230 -7323 5282 -7307
rect 5311 -7323 5363 -7307
rect 5392 -7273 5444 -7271
rect 5392 -7307 5394 -7273
rect 5394 -7307 5428 -7273
rect 5428 -7307 5444 -7273
rect 5392 -7323 5444 -7307
rect 4094 -7381 4098 -7375
rect 4098 -7381 4132 -7375
rect 4132 -7381 4146 -7375
rect 4175 -7381 4204 -7375
rect 4204 -7381 4227 -7375
rect 4256 -7381 4276 -7375
rect 4276 -7381 4308 -7375
rect 4337 -7381 4348 -7375
rect 4348 -7381 4386 -7375
rect 4386 -7381 4389 -7375
rect 4418 -7381 4420 -7375
rect 4420 -7381 4458 -7375
rect 4458 -7381 4470 -7375
rect 4499 -7381 4530 -7375
rect 4530 -7381 4551 -7375
rect 4580 -7381 4602 -7375
rect 4602 -7381 4632 -7375
rect 4662 -7381 4674 -7375
rect 4674 -7381 4708 -7375
rect 4708 -7381 4714 -7375
rect 4094 -7421 4146 -7381
rect 4175 -7421 4227 -7381
rect 4256 -7421 4308 -7381
rect 4337 -7421 4389 -7381
rect 4418 -7421 4470 -7381
rect 4499 -7421 4551 -7381
rect 4580 -7421 4632 -7381
rect 4662 -7421 4714 -7381
rect 4094 -7427 4098 -7421
rect 4098 -7427 4132 -7421
rect 4132 -7427 4146 -7421
rect 4175 -7427 4204 -7421
rect 4204 -7427 4227 -7421
rect 4256 -7427 4276 -7421
rect 4276 -7427 4308 -7421
rect 4337 -7427 4348 -7421
rect 4348 -7427 4386 -7421
rect 4386 -7427 4389 -7421
rect 4418 -7427 4420 -7421
rect 4420 -7427 4458 -7421
rect 4458 -7427 4470 -7421
rect 4499 -7427 4530 -7421
rect 4530 -7427 4551 -7421
rect 4580 -7427 4602 -7421
rect 4602 -7427 4632 -7421
rect 4662 -7427 4674 -7421
rect 4674 -7427 4708 -7421
rect 4708 -7427 4714 -7421
rect 4743 -7381 4746 -7375
rect 4746 -7381 4780 -7375
rect 4780 -7381 4795 -7375
rect 4824 -7381 4852 -7375
rect 4852 -7381 4876 -7375
rect 4905 -7381 4924 -7375
rect 4924 -7381 4957 -7375
rect 4986 -7381 4996 -7375
rect 4996 -7381 5034 -7375
rect 5034 -7381 5038 -7375
rect 5067 -7381 5068 -7375
rect 5068 -7381 5106 -7375
rect 5106 -7381 5119 -7375
rect 5148 -7381 5178 -7375
rect 5178 -7381 5200 -7375
rect 5230 -7381 5250 -7375
rect 5250 -7381 5282 -7375
rect 5311 -7381 5322 -7375
rect 5322 -7381 5356 -7375
rect 5356 -7381 5363 -7375
rect 4743 -7421 4795 -7381
rect 4824 -7421 4876 -7381
rect 4905 -7421 4957 -7381
rect 4986 -7421 5038 -7381
rect 5067 -7421 5119 -7381
rect 5148 -7421 5200 -7381
rect 5230 -7421 5282 -7381
rect 5311 -7421 5363 -7381
rect 4743 -7427 4746 -7421
rect 4746 -7427 4780 -7421
rect 4780 -7427 4795 -7421
rect 4824 -7427 4852 -7421
rect 4852 -7427 4876 -7421
rect 4905 -7427 4924 -7421
rect 4924 -7427 4957 -7421
rect 4986 -7427 4996 -7421
rect 4996 -7427 5034 -7421
rect 5034 -7427 5038 -7421
rect 5067 -7427 5068 -7421
rect 5068 -7427 5106 -7421
rect 5106 -7427 5119 -7421
rect 5148 -7427 5178 -7421
rect 5178 -7427 5200 -7421
rect 5230 -7427 5250 -7421
rect 5250 -7427 5282 -7421
rect 5311 -7427 5322 -7421
rect 5322 -7427 5356 -7421
rect 5356 -7427 5363 -7421
rect 5392 -7381 5394 -7375
rect 5394 -7381 5428 -7375
rect 5428 -7381 5444 -7375
rect 5392 -7421 5444 -7381
rect 5392 -7427 5394 -7421
rect 5394 -7427 5428 -7421
rect 5428 -7427 5444 -7421
rect 4094 -7495 4146 -7479
rect 4175 -7495 4227 -7479
rect 4256 -7495 4308 -7479
rect 4337 -7495 4389 -7479
rect 4418 -7495 4470 -7479
rect 4499 -7495 4551 -7479
rect 4580 -7495 4632 -7479
rect 4662 -7495 4714 -7479
rect 4094 -7529 4098 -7495
rect 4098 -7529 4132 -7495
rect 4132 -7529 4146 -7495
rect 4175 -7529 4204 -7495
rect 4204 -7529 4227 -7495
rect 4256 -7529 4276 -7495
rect 4276 -7529 4308 -7495
rect 4337 -7529 4348 -7495
rect 4348 -7529 4386 -7495
rect 4386 -7529 4389 -7495
rect 4418 -7529 4420 -7495
rect 4420 -7529 4458 -7495
rect 4458 -7529 4470 -7495
rect 4499 -7529 4530 -7495
rect 4530 -7529 4551 -7495
rect 4580 -7529 4602 -7495
rect 4602 -7529 4632 -7495
rect 4662 -7529 4674 -7495
rect 4674 -7529 4708 -7495
rect 4708 -7529 4714 -7495
rect 4094 -7531 4146 -7529
rect 4175 -7531 4227 -7529
rect 4256 -7531 4308 -7529
rect 4337 -7531 4389 -7529
rect 4418 -7531 4470 -7529
rect 4499 -7531 4551 -7529
rect 4580 -7531 4632 -7529
rect 4662 -7531 4714 -7529
rect 4743 -7495 4795 -7479
rect 4824 -7495 4876 -7479
rect 4905 -7495 4957 -7479
rect 4986 -7495 5038 -7479
rect 5067 -7495 5119 -7479
rect 5148 -7495 5200 -7479
rect 5230 -7495 5282 -7479
rect 5311 -7495 5363 -7479
rect 4743 -7529 4746 -7495
rect 4746 -7529 4780 -7495
rect 4780 -7529 4795 -7495
rect 4824 -7529 4852 -7495
rect 4852 -7529 4876 -7495
rect 4905 -7529 4924 -7495
rect 4924 -7529 4957 -7495
rect 4986 -7529 4996 -7495
rect 4996 -7529 5034 -7495
rect 5034 -7529 5038 -7495
rect 5067 -7529 5068 -7495
rect 5068 -7529 5106 -7495
rect 5106 -7529 5119 -7495
rect 5148 -7529 5178 -7495
rect 5178 -7529 5200 -7495
rect 5230 -7529 5250 -7495
rect 5250 -7529 5282 -7495
rect 5311 -7529 5322 -7495
rect 5322 -7529 5356 -7495
rect 5356 -7529 5363 -7495
rect 4743 -7531 4795 -7529
rect 4824 -7531 4876 -7529
rect 4905 -7531 4957 -7529
rect 4986 -7531 5038 -7529
rect 5067 -7531 5119 -7529
rect 5148 -7531 5200 -7529
rect 5230 -7531 5282 -7529
rect 5311 -7531 5363 -7529
rect 5392 -7495 5444 -7479
rect 5392 -7529 5394 -7495
rect 5394 -7529 5428 -7495
rect 5428 -7529 5444 -7495
rect 5392 -7531 5444 -7529
rect 4094 -7603 4098 -7583
rect 4098 -7603 4132 -7583
rect 4132 -7603 4146 -7583
rect 4175 -7603 4204 -7583
rect 4204 -7603 4227 -7583
rect 4256 -7603 4276 -7583
rect 4276 -7603 4308 -7583
rect 4337 -7603 4348 -7583
rect 4348 -7603 4386 -7583
rect 4386 -7603 4389 -7583
rect 4418 -7603 4420 -7583
rect 4420 -7603 4458 -7583
rect 4458 -7603 4470 -7583
rect 4499 -7603 4530 -7583
rect 4530 -7603 4551 -7583
rect 4580 -7603 4602 -7583
rect 4602 -7603 4632 -7583
rect 4662 -7603 4674 -7583
rect 4674 -7603 4708 -7583
rect 4708 -7603 4714 -7583
rect 4094 -7635 4146 -7603
rect 4175 -7635 4227 -7603
rect 4256 -7635 4308 -7603
rect 4337 -7635 4389 -7603
rect 4418 -7635 4470 -7603
rect 4499 -7635 4551 -7603
rect 4580 -7635 4632 -7603
rect 4662 -7635 4714 -7603
rect 4743 -7603 4746 -7583
rect 4746 -7603 4780 -7583
rect 4780 -7603 4795 -7583
rect 4824 -7603 4852 -7583
rect 4852 -7603 4876 -7583
rect 4905 -7603 4924 -7583
rect 4924 -7603 4957 -7583
rect 4986 -7603 4996 -7583
rect 4996 -7603 5034 -7583
rect 5034 -7603 5038 -7583
rect 5067 -7603 5068 -7583
rect 5068 -7603 5106 -7583
rect 5106 -7603 5119 -7583
rect 5148 -7603 5178 -7583
rect 5178 -7603 5200 -7583
rect 5230 -7603 5250 -7583
rect 5250 -7603 5282 -7583
rect 5311 -7603 5322 -7583
rect 5322 -7603 5356 -7583
rect 5356 -7603 5363 -7583
rect 4743 -7635 4795 -7603
rect 4824 -7635 4876 -7603
rect 4905 -7635 4957 -7603
rect 4986 -7635 5038 -7603
rect 5067 -7635 5119 -7603
rect 5148 -7635 5200 -7603
rect 5230 -7635 5282 -7603
rect 5311 -7635 5363 -7603
rect 5392 -7603 5394 -7583
rect 5394 -7603 5428 -7583
rect 5428 -7603 5444 -7583
rect 5392 -7635 5444 -7603
rect 4094 -7717 4146 -7687
rect 4175 -7717 4227 -7687
rect 4256 -7717 4308 -7687
rect 4337 -7717 4389 -7687
rect 4418 -7717 4470 -7687
rect 4499 -7717 4551 -7687
rect 4580 -7717 4632 -7687
rect 4662 -7717 4714 -7687
rect 4094 -7739 4098 -7717
rect 4098 -7739 4132 -7717
rect 4132 -7739 4146 -7717
rect 4175 -7739 4204 -7717
rect 4204 -7739 4227 -7717
rect 4256 -7739 4276 -7717
rect 4276 -7739 4308 -7717
rect 4337 -7739 4348 -7717
rect 4348 -7739 4386 -7717
rect 4386 -7739 4389 -7717
rect 4418 -7739 4420 -7717
rect 4420 -7739 4458 -7717
rect 4458 -7739 4470 -7717
rect 4499 -7739 4530 -7717
rect 4530 -7739 4551 -7717
rect 4580 -7739 4602 -7717
rect 4602 -7739 4632 -7717
rect 4662 -7739 4674 -7717
rect 4674 -7739 4708 -7717
rect 4708 -7739 4714 -7717
rect 4743 -7717 4795 -7687
rect 4824 -7717 4876 -7687
rect 4905 -7717 4957 -7687
rect 4986 -7717 5038 -7687
rect 5067 -7717 5119 -7687
rect 5148 -7717 5200 -7687
rect 5230 -7717 5282 -7687
rect 5311 -7717 5363 -7687
rect 4743 -7739 4746 -7717
rect 4746 -7739 4780 -7717
rect 4780 -7739 4795 -7717
rect 4824 -7739 4852 -7717
rect 4852 -7739 4876 -7717
rect 4905 -7739 4924 -7717
rect 4924 -7739 4957 -7717
rect 4986 -7739 4996 -7717
rect 4996 -7739 5034 -7717
rect 5034 -7739 5038 -7717
rect 5067 -7739 5068 -7717
rect 5068 -7739 5106 -7717
rect 5106 -7739 5119 -7717
rect 5148 -7739 5178 -7717
rect 5178 -7739 5200 -7717
rect 5230 -7739 5250 -7717
rect 5250 -7739 5282 -7717
rect 5311 -7739 5322 -7717
rect 5322 -7739 5356 -7717
rect 5356 -7739 5363 -7717
rect 5392 -7717 5444 -7687
rect 5392 -7739 5394 -7717
rect 5394 -7739 5428 -7717
rect 5428 -7739 5444 -7717
rect 5867 -7783 5919 -7223
rect 5985 -7783 6037 -7223
rect 6103 -7783 6112 -7223
rect 6112 -7783 6146 -7223
rect 6146 -7783 6155 -7223
rect 6221 -7783 6230 -7223
rect 6230 -7783 6264 -7223
rect 6264 -7783 6273 -7223
rect 6339 -7783 6348 -7223
rect 6348 -7783 6382 -7223
rect 6382 -7783 6391 -7223
rect 6457 -7783 6466 -7223
rect 6466 -7783 6500 -7223
rect 6500 -7783 6509 -7223
rect 6575 -7783 6584 -7223
rect 6584 -7783 6618 -7223
rect 6618 -7783 6627 -7223
rect 6693 -7783 6702 -7223
rect 6702 -7783 6736 -7223
rect 6736 -7783 6745 -7223
rect 6811 -7783 6820 -7223
rect 6820 -7783 6854 -7223
rect 6854 -7783 6863 -7223
rect 6929 -7783 6938 -7223
rect 6938 -7783 6972 -7223
rect 6972 -7783 6981 -7223
rect 7047 -7783 7056 -7223
rect 7056 -7783 7090 -7223
rect 7090 -7783 7099 -7223
rect 7165 -7783 7174 -7223
rect 7174 -7783 7208 -7223
rect 7208 -7783 7217 -7223
rect 7283 -7783 7292 -7223
rect 7292 -7783 7326 -7223
rect 7326 -7783 7335 -7223
rect 7401 -7783 7410 -7223
rect 7410 -7783 7444 -7223
rect 7444 -7783 7453 -7223
rect 7519 -7783 7528 -7223
rect 7528 -7783 7562 -7223
rect 7562 -7783 7571 -7223
rect 7637 -7783 7646 -7223
rect 7646 -7783 7680 -7223
rect 7680 -7783 7689 -7223
rect 7865 -7783 7874 -7223
rect 7874 -7783 7908 -7223
rect 7908 -7783 7917 -7223
rect 7983 -7783 7992 -7223
rect 7992 -7783 8026 -7223
rect 8026 -7783 8035 -7223
rect 8101 -7783 8110 -7223
rect 8110 -7783 8144 -7223
rect 8144 -7783 8153 -7223
rect 8219 -7783 8228 -7223
rect 8228 -7783 8262 -7223
rect 8262 -7783 8271 -7223
rect 8337 -7783 8346 -7223
rect 8346 -7783 8380 -7223
rect 8380 -7783 8389 -7223
rect 8455 -7783 8464 -7223
rect 8464 -7783 8498 -7223
rect 8498 -7783 8507 -7223
rect 8573 -7783 8582 -7223
rect 8582 -7783 8616 -7223
rect 8616 -7783 8625 -7223
rect 8691 -7783 8700 -7223
rect 8700 -7783 8734 -7223
rect 8734 -7783 8743 -7223
rect 8809 -7783 8818 -7223
rect 8818 -7783 8852 -7223
rect 8852 -7783 8861 -7223
rect 8927 -7783 8936 -7223
rect 8936 -7783 8970 -7223
rect 8970 -7783 8979 -7223
rect 9045 -7783 9054 -7223
rect 9054 -7783 9088 -7223
rect 9088 -7783 9097 -7223
rect 9163 -7783 9172 -7223
rect 9172 -7783 9206 -7223
rect 9206 -7783 9215 -7223
rect 9281 -7783 9290 -7223
rect 9290 -7783 9324 -7223
rect 9324 -7783 9333 -7223
rect 9399 -7783 9408 -7223
rect 9408 -7783 9442 -7223
rect 9442 -7783 9451 -7223
rect 9517 -7783 9526 -7223
rect 9526 -7783 9560 -7223
rect 9560 -7783 9569 -7223
rect 9635 -7783 9644 -7223
rect 9644 -7783 9678 -7223
rect 9678 -7783 9687 -7223
rect 9839 -7258 9891 -7223
rect 9919 -7258 9971 -7223
rect 9999 -7258 10051 -7223
rect 10079 -7258 10131 -7223
rect 10159 -7258 10211 -7223
rect 10239 -7258 10291 -7223
rect 10319 -7258 10371 -7206
rect 9839 -7297 9868 -7285
rect 9868 -7297 9891 -7285
rect 9919 -7297 9940 -7285
rect 9940 -7297 9971 -7285
rect 9999 -7297 10012 -7285
rect 10012 -7297 10050 -7285
rect 10050 -7297 10051 -7285
rect 10079 -7297 10084 -7285
rect 10084 -7297 10122 -7285
rect 10122 -7297 10131 -7285
rect 10159 -7297 10194 -7285
rect 10194 -7297 10211 -7285
rect 10239 -7297 10266 -7285
rect 10266 -7297 10291 -7285
rect 9839 -7337 9891 -7297
rect 9919 -7337 9971 -7297
rect 9999 -7337 10051 -7297
rect 10079 -7337 10131 -7297
rect 10159 -7337 10211 -7297
rect 10239 -7337 10291 -7297
rect 10319 -7337 10371 -7285
rect 9839 -7371 9868 -7354
rect 9868 -7371 9891 -7354
rect 9919 -7371 9940 -7354
rect 9940 -7371 9971 -7354
rect 9999 -7371 10012 -7354
rect 10012 -7371 10050 -7354
rect 10050 -7371 10051 -7354
rect 10079 -7371 10084 -7354
rect 10084 -7371 10122 -7354
rect 10122 -7371 10131 -7354
rect 10159 -7371 10194 -7354
rect 10194 -7371 10211 -7354
rect 10239 -7371 10266 -7354
rect 10266 -7371 10291 -7354
rect 9839 -7406 9891 -7371
rect 9919 -7406 9971 -7371
rect 9999 -7406 10051 -7371
rect 10079 -7406 10131 -7371
rect 10159 -7406 10211 -7371
rect 10239 -7406 10291 -7371
rect 10319 -7406 10371 -7354
rect 9839 -7445 9868 -7433
rect 9868 -7445 9891 -7433
rect 9919 -7445 9940 -7433
rect 9940 -7445 9971 -7433
rect 9999 -7445 10012 -7433
rect 10012 -7445 10050 -7433
rect 10050 -7445 10051 -7433
rect 10079 -7445 10084 -7433
rect 10084 -7445 10122 -7433
rect 10122 -7445 10131 -7433
rect 10159 -7445 10194 -7433
rect 10194 -7445 10211 -7433
rect 10239 -7445 10266 -7433
rect 10266 -7445 10291 -7433
rect 9839 -7485 9891 -7445
rect 9919 -7485 9971 -7445
rect 9999 -7485 10051 -7445
rect 10079 -7485 10131 -7445
rect 10159 -7485 10211 -7445
rect 10239 -7485 10291 -7445
rect 10319 -7485 10371 -7433
rect 10513 -7515 10565 -7395
rect 10627 -7515 10679 -7395
rect 10829 -7503 10851 -7395
rect 10851 -7503 10881 -7395
rect 10829 -7515 10881 -7503
rect 10943 -7503 10973 -7395
rect 10973 -7503 10995 -7395
rect 10943 -7515 10995 -7503
rect 11145 -7503 11167 -7395
rect 11167 -7503 11197 -7395
rect 11145 -7515 11197 -7503
rect 11259 -7503 11289 -7395
rect 11289 -7503 11311 -7395
rect 11259 -7515 11311 -7503
rect 11461 -7503 11483 -7395
rect 11483 -7503 11513 -7395
rect 11461 -7515 11513 -7503
rect 11575 -7503 11605 -7395
rect 11605 -7503 11627 -7395
rect 11575 -7515 11627 -7503
rect 11777 -7503 11799 -7395
rect 11799 -7503 11829 -7395
rect 11777 -7515 11829 -7503
rect 11891 -7503 11921 -7395
rect 11921 -7503 11943 -7395
rect 11891 -7515 11943 -7503
rect 12093 -7503 12115 -7395
rect 12115 -7503 12145 -7395
rect 12093 -7515 12145 -7503
rect 12207 -7503 12237 -7395
rect 12237 -7503 12259 -7395
rect 12207 -7515 12259 -7503
rect 4094 -7825 4098 -7791
rect 4098 -7825 4132 -7791
rect 4132 -7825 4146 -7791
rect 4175 -7825 4204 -7791
rect 4204 -7825 4227 -7791
rect 4256 -7825 4276 -7791
rect 4276 -7825 4308 -7791
rect 4337 -7825 4348 -7791
rect 4348 -7825 4386 -7791
rect 4386 -7825 4389 -7791
rect 4418 -7825 4420 -7791
rect 4420 -7825 4458 -7791
rect 4458 -7825 4470 -7791
rect 4499 -7825 4530 -7791
rect 4530 -7825 4551 -7791
rect 4580 -7825 4602 -7791
rect 4602 -7825 4632 -7791
rect 4662 -7825 4674 -7791
rect 4674 -7825 4708 -7791
rect 4708 -7825 4714 -7791
rect 4094 -7843 4146 -7825
rect 4175 -7843 4227 -7825
rect 4256 -7843 4308 -7825
rect 4337 -7843 4389 -7825
rect 4418 -7843 4470 -7825
rect 4499 -7843 4551 -7825
rect 4580 -7843 4632 -7825
rect 4662 -7843 4714 -7825
rect 4743 -7825 4746 -7791
rect 4746 -7825 4780 -7791
rect 4780 -7825 4795 -7791
rect 4824 -7825 4852 -7791
rect 4852 -7825 4876 -7791
rect 4905 -7825 4924 -7791
rect 4924 -7825 4957 -7791
rect 4986 -7825 4996 -7791
rect 4996 -7825 5034 -7791
rect 5034 -7825 5038 -7791
rect 5067 -7825 5068 -7791
rect 5068 -7825 5106 -7791
rect 5106 -7825 5119 -7791
rect 5148 -7825 5178 -7791
rect 5178 -7825 5200 -7791
rect 5230 -7825 5250 -7791
rect 5250 -7825 5282 -7791
rect 5311 -7825 5322 -7791
rect 5322 -7825 5356 -7791
rect 5356 -7825 5363 -7791
rect 4743 -7843 4795 -7825
rect 4824 -7843 4876 -7825
rect 4905 -7843 4957 -7825
rect 4986 -7843 5038 -7825
rect 5067 -7843 5119 -7825
rect 5148 -7843 5200 -7825
rect 5230 -7843 5282 -7825
rect 5311 -7843 5363 -7825
rect 5392 -7825 5394 -7791
rect 5394 -7825 5428 -7791
rect 5428 -7825 5444 -7791
rect 5392 -7843 5444 -7825
rect 4094 -7899 4098 -7895
rect 4098 -7899 4132 -7895
rect 4132 -7899 4146 -7895
rect 4175 -7899 4204 -7895
rect 4204 -7899 4227 -7895
rect 4256 -7899 4276 -7895
rect 4276 -7899 4308 -7895
rect 4337 -7899 4348 -7895
rect 4348 -7899 4386 -7895
rect 4386 -7899 4389 -7895
rect 4418 -7899 4420 -7895
rect 4420 -7899 4458 -7895
rect 4458 -7899 4470 -7895
rect 4499 -7899 4530 -7895
rect 4530 -7899 4551 -7895
rect 4580 -7899 4602 -7895
rect 4602 -7899 4632 -7895
rect 4662 -7899 4674 -7895
rect 4674 -7899 4708 -7895
rect 4708 -7899 4714 -7895
rect 4094 -7939 4146 -7899
rect 4175 -7939 4227 -7899
rect 4256 -7939 4308 -7899
rect 4337 -7939 4389 -7899
rect 4418 -7939 4470 -7899
rect 4499 -7939 4551 -7899
rect 4580 -7939 4632 -7899
rect 4662 -7939 4714 -7899
rect 4094 -7947 4098 -7939
rect 4098 -7947 4132 -7939
rect 4132 -7947 4146 -7939
rect 4175 -7947 4204 -7939
rect 4204 -7947 4227 -7939
rect 4256 -7947 4276 -7939
rect 4276 -7947 4308 -7939
rect 4337 -7947 4348 -7939
rect 4348 -7947 4386 -7939
rect 4386 -7947 4389 -7939
rect 4418 -7947 4420 -7939
rect 4420 -7947 4458 -7939
rect 4458 -7947 4470 -7939
rect 4499 -7947 4530 -7939
rect 4530 -7947 4551 -7939
rect 4580 -7947 4602 -7939
rect 4602 -7947 4632 -7939
rect 4662 -7947 4674 -7939
rect 4674 -7947 4708 -7939
rect 4708 -7947 4714 -7939
rect 4743 -7899 4746 -7895
rect 4746 -7899 4780 -7895
rect 4780 -7899 4795 -7895
rect 4824 -7899 4852 -7895
rect 4852 -7899 4876 -7895
rect 4905 -7899 4924 -7895
rect 4924 -7899 4957 -7895
rect 4986 -7899 4996 -7895
rect 4996 -7899 5034 -7895
rect 5034 -7899 5038 -7895
rect 5067 -7899 5068 -7895
rect 5068 -7899 5106 -7895
rect 5106 -7899 5119 -7895
rect 5148 -7899 5178 -7895
rect 5178 -7899 5200 -7895
rect 5230 -7899 5250 -7895
rect 5250 -7899 5282 -7895
rect 5311 -7899 5322 -7895
rect 5322 -7899 5356 -7895
rect 5356 -7899 5363 -7895
rect 4743 -7939 4795 -7899
rect 4824 -7939 4876 -7899
rect 4905 -7939 4957 -7899
rect 4986 -7939 5038 -7899
rect 5067 -7939 5119 -7899
rect 5148 -7939 5200 -7899
rect 5230 -7939 5282 -7899
rect 5311 -7939 5363 -7899
rect 4743 -7947 4746 -7939
rect 4746 -7947 4780 -7939
rect 4780 -7947 4795 -7939
rect 4824 -7947 4852 -7939
rect 4852 -7947 4876 -7939
rect 4905 -7947 4924 -7939
rect 4924 -7947 4957 -7939
rect 4986 -7947 4996 -7939
rect 4996 -7947 5034 -7939
rect 5034 -7947 5038 -7939
rect 5067 -7947 5068 -7939
rect 5068 -7947 5106 -7939
rect 5106 -7947 5119 -7939
rect 5148 -7947 5178 -7939
rect 5178 -7947 5200 -7939
rect 5230 -7947 5250 -7939
rect 5250 -7947 5282 -7939
rect 5311 -7947 5322 -7939
rect 5322 -7947 5356 -7939
rect 5356 -7947 5363 -7939
rect 5392 -7899 5394 -7895
rect 5394 -7899 5428 -7895
rect 5428 -7899 5444 -7895
rect 5392 -7939 5444 -7899
rect 5392 -7947 5394 -7939
rect 5394 -7947 5428 -7939
rect 5428 -7947 5444 -7939
rect 5923 -7841 5981 -7835
rect 5923 -7875 5935 -7841
rect 5935 -7875 5969 -7841
rect 5969 -7875 5981 -7841
rect 5923 -7949 5981 -7875
rect 5923 -7983 5935 -7949
rect 5935 -7983 5969 -7949
rect 5969 -7983 5981 -7949
rect 5923 -7989 5981 -7983
rect 6041 -7841 6099 -7835
rect 6041 -7875 6053 -7841
rect 6053 -7875 6087 -7841
rect 6087 -7875 6099 -7841
rect 6041 -7949 6099 -7875
rect 6041 -7983 6053 -7949
rect 6053 -7983 6087 -7949
rect 6087 -7983 6099 -7949
rect 6041 -7989 6099 -7983
rect 6159 -7841 6217 -7835
rect 6159 -7875 6171 -7841
rect 6171 -7875 6205 -7841
rect 6205 -7875 6217 -7841
rect 6159 -7949 6217 -7875
rect 6159 -7983 6171 -7949
rect 6171 -7983 6205 -7949
rect 6205 -7983 6217 -7949
rect 6159 -7989 6217 -7983
rect 6277 -7841 6335 -7835
rect 6277 -7875 6289 -7841
rect 6289 -7875 6323 -7841
rect 6323 -7875 6335 -7841
rect 6277 -7949 6335 -7875
rect 6277 -7983 6289 -7949
rect 6289 -7983 6323 -7949
rect 6323 -7983 6335 -7949
rect 6277 -7989 6335 -7983
rect 6395 -7841 6453 -7835
rect 6395 -7875 6407 -7841
rect 6407 -7875 6441 -7841
rect 6441 -7875 6453 -7841
rect 6395 -7949 6453 -7875
rect 6395 -7983 6407 -7949
rect 6407 -7983 6441 -7949
rect 6441 -7983 6453 -7949
rect 6395 -7989 6453 -7983
rect 6513 -7841 6571 -7835
rect 6513 -7875 6525 -7841
rect 6525 -7875 6559 -7841
rect 6559 -7875 6571 -7841
rect 6513 -7949 6571 -7875
rect 6513 -7983 6525 -7949
rect 6525 -7983 6559 -7949
rect 6559 -7983 6571 -7949
rect 6513 -7989 6571 -7983
rect 6631 -7841 6689 -7835
rect 6631 -7875 6643 -7841
rect 6643 -7875 6677 -7841
rect 6677 -7875 6689 -7841
rect 6631 -7949 6689 -7875
rect 6631 -7983 6643 -7949
rect 6643 -7983 6677 -7949
rect 6677 -7983 6689 -7949
rect 6631 -7989 6689 -7983
rect 6749 -7841 6807 -7835
rect 6749 -7875 6761 -7841
rect 6761 -7875 6795 -7841
rect 6795 -7875 6807 -7841
rect 6749 -7949 6807 -7875
rect 6749 -7983 6761 -7949
rect 6761 -7983 6795 -7949
rect 6795 -7983 6807 -7949
rect 6749 -7989 6807 -7983
rect 6867 -7841 6925 -7835
rect 6867 -7875 6879 -7841
rect 6879 -7875 6913 -7841
rect 6913 -7875 6925 -7841
rect 6867 -7949 6925 -7875
rect 6867 -7983 6879 -7949
rect 6879 -7983 6913 -7949
rect 6913 -7983 6925 -7949
rect 6867 -7989 6925 -7983
rect 6985 -7841 7043 -7835
rect 6985 -7875 6997 -7841
rect 6997 -7875 7031 -7841
rect 7031 -7875 7043 -7841
rect 6985 -7949 7043 -7875
rect 6985 -7983 6997 -7949
rect 6997 -7983 7031 -7949
rect 7031 -7983 7043 -7949
rect 6985 -7989 7043 -7983
rect 7103 -7841 7161 -7835
rect 7103 -7875 7115 -7841
rect 7115 -7875 7149 -7841
rect 7149 -7875 7161 -7841
rect 7103 -7949 7161 -7875
rect 7103 -7983 7115 -7949
rect 7115 -7983 7149 -7949
rect 7149 -7983 7161 -7949
rect 7103 -7989 7161 -7983
rect 7221 -7841 7279 -7835
rect 7221 -7875 7233 -7841
rect 7233 -7875 7267 -7841
rect 7267 -7875 7279 -7841
rect 7221 -7949 7279 -7875
rect 7221 -7983 7233 -7949
rect 7233 -7983 7267 -7949
rect 7267 -7983 7279 -7949
rect 7221 -7989 7279 -7983
rect 7339 -7841 7397 -7835
rect 7339 -7875 7351 -7841
rect 7351 -7875 7385 -7841
rect 7385 -7875 7397 -7841
rect 7339 -7949 7397 -7875
rect 7339 -7983 7351 -7949
rect 7351 -7983 7385 -7949
rect 7385 -7983 7397 -7949
rect 7339 -7989 7397 -7983
rect 7457 -7841 7515 -7835
rect 7457 -7875 7469 -7841
rect 7469 -7875 7503 -7841
rect 7503 -7875 7515 -7841
rect 7457 -7949 7515 -7875
rect 7457 -7983 7469 -7949
rect 7469 -7983 7503 -7949
rect 7503 -7983 7515 -7949
rect 7457 -7989 7515 -7983
rect 7575 -7841 7633 -7835
rect 7575 -7875 7587 -7841
rect 7587 -7875 7621 -7841
rect 7621 -7875 7633 -7841
rect 7575 -7949 7633 -7875
rect 7575 -7983 7587 -7949
rect 7587 -7983 7621 -7949
rect 7621 -7983 7633 -7949
rect 7575 -7989 7633 -7983
rect 7921 -7841 7979 -7835
rect 7921 -7875 7933 -7841
rect 7933 -7875 7967 -7841
rect 7967 -7875 7979 -7841
rect 7921 -7949 7979 -7875
rect 7921 -7983 7933 -7949
rect 7933 -7983 7967 -7949
rect 7967 -7983 7979 -7949
rect 7921 -7989 7979 -7983
rect 8039 -7841 8097 -7835
rect 8039 -7875 8051 -7841
rect 8051 -7875 8085 -7841
rect 8085 -7875 8097 -7841
rect 8039 -7949 8097 -7875
rect 8039 -7983 8051 -7949
rect 8051 -7983 8085 -7949
rect 8085 -7983 8097 -7949
rect 8039 -7989 8097 -7983
rect 8157 -7841 8215 -7835
rect 8157 -7875 8169 -7841
rect 8169 -7875 8203 -7841
rect 8203 -7875 8215 -7841
rect 8157 -7949 8215 -7875
rect 8157 -7983 8169 -7949
rect 8169 -7983 8203 -7949
rect 8203 -7983 8215 -7949
rect 8157 -7989 8215 -7983
rect 8275 -7841 8333 -7835
rect 8275 -7875 8287 -7841
rect 8287 -7875 8321 -7841
rect 8321 -7875 8333 -7841
rect 8275 -7949 8333 -7875
rect 8275 -7983 8287 -7949
rect 8287 -7983 8321 -7949
rect 8321 -7983 8333 -7949
rect 8275 -7989 8333 -7983
rect 8393 -7841 8451 -7835
rect 8393 -7875 8405 -7841
rect 8405 -7875 8439 -7841
rect 8439 -7875 8451 -7841
rect 8393 -7949 8451 -7875
rect 8393 -7983 8405 -7949
rect 8405 -7983 8439 -7949
rect 8439 -7983 8451 -7949
rect 8393 -7989 8451 -7983
rect 8511 -7841 8569 -7835
rect 8511 -7875 8523 -7841
rect 8523 -7875 8557 -7841
rect 8557 -7875 8569 -7841
rect 8511 -7949 8569 -7875
rect 8511 -7983 8523 -7949
rect 8523 -7983 8557 -7949
rect 8557 -7983 8569 -7949
rect 8511 -7989 8569 -7983
rect 8629 -7841 8687 -7835
rect 8629 -7875 8641 -7841
rect 8641 -7875 8675 -7841
rect 8675 -7875 8687 -7841
rect 8629 -7949 8687 -7875
rect 8629 -7983 8641 -7949
rect 8641 -7983 8675 -7949
rect 8675 -7983 8687 -7949
rect 8629 -7989 8687 -7983
rect 8747 -7841 8805 -7835
rect 8747 -7875 8759 -7841
rect 8759 -7875 8793 -7841
rect 8793 -7875 8805 -7841
rect 8747 -7949 8805 -7875
rect 8747 -7983 8759 -7949
rect 8759 -7983 8793 -7949
rect 8793 -7983 8805 -7949
rect 8747 -7989 8805 -7983
rect 8865 -7841 8923 -7835
rect 8865 -7875 8877 -7841
rect 8877 -7875 8911 -7841
rect 8911 -7875 8923 -7841
rect 8865 -7949 8923 -7875
rect 8865 -7983 8877 -7949
rect 8877 -7983 8911 -7949
rect 8911 -7983 8923 -7949
rect 8865 -7989 8923 -7983
rect 8983 -7841 9041 -7835
rect 8983 -7875 8995 -7841
rect 8995 -7875 9029 -7841
rect 9029 -7875 9041 -7841
rect 8983 -7949 9041 -7875
rect 8983 -7983 8995 -7949
rect 8995 -7983 9029 -7949
rect 9029 -7983 9041 -7949
rect 8983 -7989 9041 -7983
rect 9101 -7841 9159 -7835
rect 9101 -7875 9113 -7841
rect 9113 -7875 9147 -7841
rect 9147 -7875 9159 -7841
rect 9101 -7949 9159 -7875
rect 9101 -7983 9113 -7949
rect 9113 -7983 9147 -7949
rect 9147 -7983 9159 -7949
rect 9101 -7989 9159 -7983
rect 9219 -7841 9277 -7835
rect 9219 -7875 9231 -7841
rect 9231 -7875 9265 -7841
rect 9265 -7875 9277 -7841
rect 9219 -7949 9277 -7875
rect 9219 -7983 9231 -7949
rect 9231 -7983 9265 -7949
rect 9265 -7983 9277 -7949
rect 9219 -7989 9277 -7983
rect 9337 -7841 9395 -7835
rect 9337 -7875 9349 -7841
rect 9349 -7875 9383 -7841
rect 9383 -7875 9395 -7841
rect 9337 -7949 9395 -7875
rect 9337 -7983 9349 -7949
rect 9349 -7983 9383 -7949
rect 9383 -7983 9395 -7949
rect 9337 -7989 9395 -7983
rect 9455 -7841 9513 -7835
rect 9455 -7875 9467 -7841
rect 9467 -7875 9501 -7841
rect 9501 -7875 9513 -7841
rect 9455 -7949 9513 -7875
rect 9455 -7983 9467 -7949
rect 9467 -7983 9501 -7949
rect 9501 -7983 9513 -7949
rect 9455 -7989 9513 -7983
rect 9573 -7841 9631 -7835
rect 9573 -7875 9585 -7841
rect 9585 -7875 9619 -7841
rect 9619 -7875 9631 -7841
rect 9573 -7949 9631 -7875
rect 9573 -7983 9585 -7949
rect 9585 -7983 9619 -7949
rect 9619 -7983 9631 -7949
rect 9573 -7989 9631 -7983
rect 4094 -8013 4146 -7999
rect 4175 -8013 4227 -7999
rect 4256 -8013 4308 -7999
rect 4337 -8013 4389 -7999
rect 4418 -8013 4470 -7999
rect 4499 -8013 4551 -7999
rect 4580 -8013 4632 -7999
rect 4662 -8013 4714 -7999
rect 4094 -8047 4098 -8013
rect 4098 -8047 4132 -8013
rect 4132 -8047 4146 -8013
rect 4175 -8047 4204 -8013
rect 4204 -8047 4227 -8013
rect 4256 -8047 4276 -8013
rect 4276 -8047 4308 -8013
rect 4337 -8047 4348 -8013
rect 4348 -8047 4386 -8013
rect 4386 -8047 4389 -8013
rect 4418 -8047 4420 -8013
rect 4420 -8047 4458 -8013
rect 4458 -8047 4470 -8013
rect 4499 -8047 4530 -8013
rect 4530 -8047 4551 -8013
rect 4580 -8047 4602 -8013
rect 4602 -8047 4632 -8013
rect 4662 -8047 4674 -8013
rect 4674 -8047 4708 -8013
rect 4708 -8047 4714 -8013
rect 4094 -8051 4146 -8047
rect 4175 -8051 4227 -8047
rect 4256 -8051 4308 -8047
rect 4337 -8051 4389 -8047
rect 4418 -8051 4470 -8047
rect 4499 -8051 4551 -8047
rect 4580 -8051 4632 -8047
rect 4662 -8051 4714 -8047
rect 4743 -8013 4795 -7999
rect 4824 -8013 4876 -7999
rect 4905 -8013 4957 -7999
rect 4986 -8013 5038 -7999
rect 5067 -8013 5119 -7999
rect 5148 -8013 5200 -7999
rect 5230 -8013 5282 -7999
rect 5311 -8013 5363 -7999
rect 4743 -8047 4746 -8013
rect 4746 -8047 4780 -8013
rect 4780 -8047 4795 -8013
rect 4824 -8047 4852 -8013
rect 4852 -8047 4876 -8013
rect 4905 -8047 4924 -8013
rect 4924 -8047 4957 -8013
rect 4986 -8047 4996 -8013
rect 4996 -8047 5034 -8013
rect 5034 -8047 5038 -8013
rect 5067 -8047 5068 -8013
rect 5068 -8047 5106 -8013
rect 5106 -8047 5119 -8013
rect 5148 -8047 5178 -8013
rect 5178 -8047 5200 -8013
rect 5230 -8047 5250 -8013
rect 5250 -8047 5282 -8013
rect 5311 -8047 5322 -8013
rect 5322 -8047 5356 -8013
rect 5356 -8047 5363 -8013
rect 4743 -8051 4795 -8047
rect 4824 -8051 4876 -8047
rect 4905 -8051 4957 -8047
rect 4986 -8051 5038 -8047
rect 5067 -8051 5119 -8047
rect 5148 -8051 5200 -8047
rect 5230 -8051 5282 -8047
rect 5311 -8051 5363 -8047
rect 5392 -8013 5444 -7999
rect 5392 -8047 5394 -8013
rect 5394 -8047 5428 -8013
rect 5428 -8047 5444 -8013
rect 5392 -8051 5444 -8047
rect 4094 -8121 4098 -8103
rect 4098 -8121 4132 -8103
rect 4132 -8121 4146 -8103
rect 4175 -8121 4204 -8103
rect 4204 -8121 4227 -8103
rect 4256 -8121 4276 -8103
rect 4276 -8121 4308 -8103
rect 4337 -8121 4348 -8103
rect 4348 -8121 4386 -8103
rect 4386 -8121 4389 -8103
rect 4418 -8121 4420 -8103
rect 4420 -8121 4458 -8103
rect 4458 -8121 4470 -8103
rect 4499 -8121 4530 -8103
rect 4530 -8121 4551 -8103
rect 4580 -8121 4602 -8103
rect 4602 -8121 4632 -8103
rect 4662 -8121 4674 -8103
rect 4674 -8121 4708 -8103
rect 4708 -8121 4714 -8103
rect 4094 -8155 4146 -8121
rect 4175 -8155 4227 -8121
rect 4256 -8155 4308 -8121
rect 4337 -8155 4389 -8121
rect 4418 -8155 4470 -8121
rect 4499 -8155 4551 -8121
rect 4580 -8155 4632 -8121
rect 4662 -8155 4714 -8121
rect 4743 -8121 4746 -8103
rect 4746 -8121 4780 -8103
rect 4780 -8121 4795 -8103
rect 4824 -8121 4852 -8103
rect 4852 -8121 4876 -8103
rect 4905 -8121 4924 -8103
rect 4924 -8121 4957 -8103
rect 4986 -8121 4996 -8103
rect 4996 -8121 5034 -8103
rect 5034 -8121 5038 -8103
rect 5067 -8121 5068 -8103
rect 5068 -8121 5106 -8103
rect 5106 -8121 5119 -8103
rect 5148 -8121 5178 -8103
rect 5178 -8121 5200 -8103
rect 5230 -8121 5250 -8103
rect 5250 -8121 5282 -8103
rect 5311 -8121 5322 -8103
rect 5322 -8121 5356 -8103
rect 5356 -8121 5363 -8103
rect 4743 -8155 4795 -8121
rect 4824 -8155 4876 -8121
rect 4905 -8155 4957 -8121
rect 4986 -8155 5038 -8121
rect 5067 -8155 5119 -8121
rect 5148 -8155 5200 -8121
rect 5230 -8155 5282 -8121
rect 5311 -8155 5363 -8121
rect 5392 -8121 5394 -8103
rect 5394 -8121 5428 -8103
rect 5428 -8121 5444 -8103
rect 5392 -8155 5444 -8121
rect 4094 -8235 4146 -8207
rect 4175 -8235 4227 -8207
rect 4256 -8235 4308 -8207
rect 4337 -8235 4389 -8207
rect 4418 -8235 4470 -8207
rect 4499 -8235 4551 -8207
rect 4580 -8235 4632 -8207
rect 4662 -8235 4714 -8207
rect 4094 -8259 4098 -8235
rect 4098 -8259 4132 -8235
rect 4132 -8259 4146 -8235
rect 4175 -8259 4204 -8235
rect 4204 -8259 4227 -8235
rect 4256 -8259 4276 -8235
rect 4276 -8259 4308 -8235
rect 4337 -8259 4348 -8235
rect 4348 -8259 4386 -8235
rect 4386 -8259 4389 -8235
rect 4418 -8259 4420 -8235
rect 4420 -8259 4458 -8235
rect 4458 -8259 4470 -8235
rect 4499 -8259 4530 -8235
rect 4530 -8259 4551 -8235
rect 4580 -8259 4602 -8235
rect 4602 -8259 4632 -8235
rect 4662 -8259 4674 -8235
rect 4674 -8259 4708 -8235
rect 4708 -8259 4714 -8235
rect 4743 -8235 4795 -8207
rect 4824 -8235 4876 -8207
rect 4905 -8235 4957 -8207
rect 4986 -8235 5038 -8207
rect 5067 -8235 5119 -8207
rect 5148 -8235 5200 -8207
rect 5230 -8235 5282 -8207
rect 5311 -8235 5363 -8207
rect 4743 -8259 4746 -8235
rect 4746 -8259 4780 -8235
rect 4780 -8259 4795 -8235
rect 4824 -8259 4852 -8235
rect 4852 -8259 4876 -8235
rect 4905 -8259 4924 -8235
rect 4924 -8259 4957 -8235
rect 4986 -8259 4996 -8235
rect 4996 -8259 5034 -8235
rect 5034 -8259 5038 -8235
rect 5067 -8259 5068 -8235
rect 5068 -8259 5106 -8235
rect 5106 -8259 5119 -8235
rect 5148 -8259 5178 -8235
rect 5178 -8259 5200 -8235
rect 5230 -8259 5250 -8235
rect 5250 -8259 5282 -8235
rect 5311 -8259 5322 -8235
rect 5322 -8259 5356 -8235
rect 5356 -8259 5363 -8235
rect 5392 -8235 5444 -8207
rect 5392 -8259 5394 -8235
rect 5394 -8259 5428 -8235
rect 5428 -8259 5444 -8235
rect 4094 -8343 4098 -8311
rect 4098 -8343 4132 -8311
rect 4132 -8343 4146 -8311
rect 4175 -8343 4204 -8311
rect 4204 -8343 4227 -8311
rect 4256 -8343 4276 -8311
rect 4276 -8343 4308 -8311
rect 4337 -8343 4348 -8311
rect 4348 -8343 4386 -8311
rect 4386 -8343 4389 -8311
rect 4418 -8343 4420 -8311
rect 4420 -8343 4458 -8311
rect 4458 -8343 4470 -8311
rect 4499 -8343 4530 -8311
rect 4530 -8343 4551 -8311
rect 4580 -8343 4602 -8311
rect 4602 -8343 4632 -8311
rect 4662 -8343 4674 -8311
rect 4674 -8343 4708 -8311
rect 4708 -8343 4714 -8311
rect 4094 -8363 4146 -8343
rect 4175 -8363 4227 -8343
rect 4256 -8363 4308 -8343
rect 4337 -8363 4389 -8343
rect 4418 -8363 4470 -8343
rect 4499 -8363 4551 -8343
rect 4580 -8363 4632 -8343
rect 4662 -8363 4714 -8343
rect 4743 -8343 4746 -8311
rect 4746 -8343 4780 -8311
rect 4780 -8343 4795 -8311
rect 4824 -8343 4852 -8311
rect 4852 -8343 4876 -8311
rect 4905 -8343 4924 -8311
rect 4924 -8343 4957 -8311
rect 4986 -8343 4996 -8311
rect 4996 -8343 5034 -8311
rect 5034 -8343 5038 -8311
rect 5067 -8343 5068 -8311
rect 5068 -8343 5106 -8311
rect 5106 -8343 5119 -8311
rect 5148 -8343 5178 -8311
rect 5178 -8343 5200 -8311
rect 5230 -8343 5250 -8311
rect 5250 -8343 5282 -8311
rect 5311 -8343 5322 -8311
rect 5322 -8343 5356 -8311
rect 5356 -8343 5363 -8311
rect 4743 -8363 4795 -8343
rect 4824 -8363 4876 -8343
rect 4905 -8363 4957 -8343
rect 4986 -8363 5038 -8343
rect 5067 -8363 5119 -8343
rect 5148 -8363 5200 -8343
rect 5230 -8363 5282 -8343
rect 5311 -8363 5363 -8343
rect 5392 -8343 5394 -8311
rect 5394 -8343 5428 -8311
rect 5428 -8343 5444 -8311
rect 5392 -8363 5444 -8343
rect 4094 -8417 4098 -8415
rect 4098 -8417 4132 -8415
rect 4132 -8417 4146 -8415
rect 4175 -8417 4204 -8415
rect 4204 -8417 4227 -8415
rect 4256 -8417 4276 -8415
rect 4276 -8417 4308 -8415
rect 4337 -8417 4348 -8415
rect 4348 -8417 4386 -8415
rect 4386 -8417 4389 -8415
rect 4418 -8417 4420 -8415
rect 4420 -8417 4458 -8415
rect 4458 -8417 4470 -8415
rect 4499 -8417 4530 -8415
rect 4530 -8417 4551 -8415
rect 4580 -8417 4602 -8415
rect 4602 -8417 4632 -8415
rect 4662 -8417 4674 -8415
rect 4674 -8417 4708 -8415
rect 4708 -8417 4714 -8415
rect 4094 -8457 4146 -8417
rect 4175 -8457 4227 -8417
rect 4256 -8457 4308 -8417
rect 4337 -8457 4389 -8417
rect 4418 -8457 4470 -8417
rect 4499 -8457 4551 -8417
rect 4580 -8457 4632 -8417
rect 4662 -8457 4714 -8417
rect 4094 -8467 4098 -8457
rect 4098 -8467 4132 -8457
rect 4132 -8467 4146 -8457
rect 4175 -8467 4204 -8457
rect 4204 -8467 4227 -8457
rect 4256 -8467 4276 -8457
rect 4276 -8467 4308 -8457
rect 4337 -8467 4348 -8457
rect 4348 -8467 4386 -8457
rect 4386 -8467 4389 -8457
rect 4418 -8467 4420 -8457
rect 4420 -8467 4458 -8457
rect 4458 -8467 4470 -8457
rect 4499 -8467 4530 -8457
rect 4530 -8467 4551 -8457
rect 4580 -8467 4602 -8457
rect 4602 -8467 4632 -8457
rect 4662 -8467 4674 -8457
rect 4674 -8467 4708 -8457
rect 4708 -8467 4714 -8457
rect 4743 -8417 4746 -8415
rect 4746 -8417 4780 -8415
rect 4780 -8417 4795 -8415
rect 4824 -8417 4852 -8415
rect 4852 -8417 4876 -8415
rect 4905 -8417 4924 -8415
rect 4924 -8417 4957 -8415
rect 4986 -8417 4996 -8415
rect 4996 -8417 5034 -8415
rect 5034 -8417 5038 -8415
rect 5067 -8417 5068 -8415
rect 5068 -8417 5106 -8415
rect 5106 -8417 5119 -8415
rect 5148 -8417 5178 -8415
rect 5178 -8417 5200 -8415
rect 5230 -8417 5250 -8415
rect 5250 -8417 5282 -8415
rect 5311 -8417 5322 -8415
rect 5322 -8417 5356 -8415
rect 5356 -8417 5363 -8415
rect 4743 -8457 4795 -8417
rect 4824 -8457 4876 -8417
rect 4905 -8457 4957 -8417
rect 4986 -8457 5038 -8417
rect 5067 -8457 5119 -8417
rect 5148 -8457 5200 -8417
rect 5230 -8457 5282 -8417
rect 5311 -8457 5363 -8417
rect 4743 -8467 4746 -8457
rect 4746 -8467 4780 -8457
rect 4780 -8467 4795 -8457
rect 4824 -8467 4852 -8457
rect 4852 -8467 4876 -8457
rect 4905 -8467 4924 -8457
rect 4924 -8467 4957 -8457
rect 4986 -8467 4996 -8457
rect 4996 -8467 5034 -8457
rect 5034 -8467 5038 -8457
rect 5067 -8467 5068 -8457
rect 5068 -8467 5106 -8457
rect 5106 -8467 5119 -8457
rect 5148 -8467 5178 -8457
rect 5178 -8467 5200 -8457
rect 5230 -8467 5250 -8457
rect 5250 -8467 5282 -8457
rect 5311 -8467 5322 -8457
rect 5322 -8467 5356 -8457
rect 5356 -8467 5363 -8457
rect 5392 -8417 5394 -8415
rect 5394 -8417 5428 -8415
rect 5428 -8417 5444 -8415
rect 5392 -8457 5444 -8417
rect 5392 -8467 5394 -8457
rect 5394 -8467 5428 -8457
rect 5428 -8467 5444 -8457
rect 4094 -8531 4146 -8519
rect 4175 -8531 4227 -8519
rect 4256 -8531 4308 -8519
rect 4337 -8531 4389 -8519
rect 4418 -8531 4470 -8519
rect 4499 -8531 4551 -8519
rect 4580 -8531 4632 -8519
rect 4662 -8531 4714 -8519
rect 4094 -8565 4098 -8531
rect 4098 -8565 4132 -8531
rect 4132 -8565 4146 -8531
rect 4175 -8565 4204 -8531
rect 4204 -8565 4227 -8531
rect 4256 -8565 4276 -8531
rect 4276 -8565 4308 -8531
rect 4337 -8565 4348 -8531
rect 4348 -8565 4386 -8531
rect 4386 -8565 4389 -8531
rect 4418 -8565 4420 -8531
rect 4420 -8565 4458 -8531
rect 4458 -8565 4470 -8531
rect 4499 -8565 4530 -8531
rect 4530 -8565 4551 -8531
rect 4580 -8565 4602 -8531
rect 4602 -8565 4632 -8531
rect 4662 -8565 4674 -8531
rect 4674 -8565 4708 -8531
rect 4708 -8565 4714 -8531
rect 4094 -8571 4146 -8565
rect 4175 -8571 4227 -8565
rect 4256 -8571 4308 -8565
rect 4337 -8571 4389 -8565
rect 4418 -8571 4470 -8565
rect 4499 -8571 4551 -8565
rect 4580 -8571 4632 -8565
rect 4662 -8571 4714 -8565
rect 4743 -8531 4795 -8519
rect 4824 -8531 4876 -8519
rect 4905 -8531 4957 -8519
rect 4986 -8531 5038 -8519
rect 5067 -8531 5119 -8519
rect 5148 -8531 5200 -8519
rect 5230 -8531 5282 -8519
rect 5311 -8531 5363 -8519
rect 4743 -8565 4746 -8531
rect 4746 -8565 4780 -8531
rect 4780 -8565 4795 -8531
rect 4824 -8565 4852 -8531
rect 4852 -8565 4876 -8531
rect 4905 -8565 4924 -8531
rect 4924 -8565 4957 -8531
rect 4986 -8565 4996 -8531
rect 4996 -8565 5034 -8531
rect 5034 -8565 5038 -8531
rect 5067 -8565 5068 -8531
rect 5068 -8565 5106 -8531
rect 5106 -8565 5119 -8531
rect 5148 -8565 5178 -8531
rect 5178 -8565 5200 -8531
rect 5230 -8565 5250 -8531
rect 5250 -8565 5282 -8531
rect 5311 -8565 5322 -8531
rect 5322 -8565 5356 -8531
rect 5356 -8565 5363 -8531
rect 4743 -8571 4795 -8565
rect 4824 -8571 4876 -8565
rect 4905 -8571 4957 -8565
rect 4986 -8571 5038 -8565
rect 5067 -8571 5119 -8565
rect 5148 -8571 5200 -8565
rect 5230 -8571 5282 -8565
rect 5311 -8571 5363 -8565
rect 5392 -8531 5444 -8519
rect 5392 -8565 5394 -8531
rect 5394 -8565 5428 -8531
rect 5428 -8565 5444 -8531
rect 5392 -8571 5444 -8565
rect 5867 -8601 5876 -8041
rect 5876 -8601 5910 -8041
rect 5910 -8601 5919 -8041
rect 5985 -8601 5994 -8041
rect 5994 -8601 6028 -8041
rect 6028 -8601 6037 -8041
rect 6103 -8601 6112 -8041
rect 6112 -8601 6146 -8041
rect 6146 -8601 6155 -8041
rect 6221 -8601 6230 -8041
rect 6230 -8601 6264 -8041
rect 6264 -8601 6273 -8041
rect 6339 -8601 6348 -8041
rect 6348 -8601 6382 -8041
rect 6382 -8601 6391 -8041
rect 6457 -8601 6466 -8041
rect 6466 -8601 6500 -8041
rect 6500 -8601 6509 -8041
rect 6575 -8601 6584 -8041
rect 6584 -8601 6618 -8041
rect 6618 -8601 6627 -8041
rect 6693 -8601 6702 -8041
rect 6702 -8601 6736 -8041
rect 6736 -8601 6745 -8041
rect 6811 -8601 6820 -8041
rect 6820 -8601 6854 -8041
rect 6854 -8601 6863 -8041
rect 6929 -8601 6938 -8041
rect 6938 -8601 6972 -8041
rect 6972 -8601 6981 -8041
rect 7047 -8601 7056 -8041
rect 7056 -8601 7090 -8041
rect 7090 -8601 7099 -8041
rect 7165 -8601 7174 -8041
rect 7174 -8601 7208 -8041
rect 7208 -8601 7217 -8041
rect 7283 -8601 7292 -8041
rect 7292 -8601 7326 -8041
rect 7326 -8601 7335 -8041
rect 7401 -8601 7410 -8041
rect 7410 -8601 7444 -8041
rect 7444 -8601 7453 -8041
rect 7519 -8601 7528 -8041
rect 7528 -8601 7562 -8041
rect 7562 -8601 7571 -8041
rect 7637 -8601 7646 -8041
rect 7646 -8601 7680 -8041
rect 7680 -8601 7689 -8041
rect 7865 -8601 7874 -8041
rect 7874 -8601 7908 -8041
rect 7908 -8601 7917 -8041
rect 7983 -8601 7992 -8041
rect 7992 -8601 8026 -8041
rect 8026 -8601 8035 -8041
rect 8101 -8601 8110 -8041
rect 8110 -8601 8144 -8041
rect 8144 -8601 8153 -8041
rect 8219 -8601 8228 -8041
rect 8228 -8601 8262 -8041
rect 8262 -8601 8271 -8041
rect 8337 -8601 8346 -8041
rect 8346 -8601 8380 -8041
rect 8380 -8601 8389 -8041
rect 8455 -8601 8464 -8041
rect 8464 -8601 8498 -8041
rect 8498 -8601 8507 -8041
rect 8573 -8601 8582 -8041
rect 8582 -8601 8616 -8041
rect 8616 -8601 8625 -8041
rect 8691 -8601 8700 -8041
rect 8700 -8601 8734 -8041
rect 8734 -8601 8743 -8041
rect 8809 -8601 8818 -8041
rect 8818 -8601 8852 -8041
rect 8852 -8601 8861 -8041
rect 8927 -8601 8936 -8041
rect 8936 -8601 8970 -8041
rect 8970 -8601 8979 -8041
rect 9045 -8601 9054 -8041
rect 9054 -8601 9088 -8041
rect 9088 -8601 9097 -8041
rect 9163 -8601 9172 -8041
rect 9172 -8601 9206 -8041
rect 9206 -8601 9215 -8041
rect 9281 -8601 9290 -8041
rect 9290 -8601 9324 -8041
rect 9324 -8601 9333 -8041
rect 9399 -8601 9408 -8041
rect 9408 -8601 9442 -8041
rect 9442 -8601 9451 -8041
rect 9517 -8601 9526 -8041
rect 9526 -8601 9560 -8041
rect 9560 -8601 9569 -8041
rect 9635 -8601 9644 -8041
rect 9644 -8601 9678 -8041
rect 9678 -8601 9687 -8041
rect 12525 -8059 12534 -7219
rect 12534 -8059 12568 -7219
rect 12568 -8059 12577 -7219
rect 12673 -8059 12682 -7219
rect 12682 -8059 12716 -7219
rect 12716 -8059 12725 -7219
rect 12821 -8059 12830 -7219
rect 12830 -8059 12864 -7219
rect 12864 -8059 12873 -7219
rect 12969 -8059 12978 -7219
rect 12978 -8059 13012 -7219
rect 13012 -8059 13021 -7219
rect 13117 -8059 13126 -7219
rect 13126 -8059 13160 -7219
rect 13160 -8059 13169 -7219
rect 13265 -8059 13274 -7219
rect 13274 -8059 13308 -7219
rect 13308 -8059 13317 -7219
rect 13413 -8059 13422 -7219
rect 13422 -8059 13456 -7219
rect 13456 -8059 13465 -7219
rect 13561 -8059 13570 -7219
rect 13570 -8059 13604 -7219
rect 13604 -8059 13613 -7219
rect 13709 -8059 13718 -7219
rect 13718 -8059 13752 -7219
rect 13752 -8059 13761 -7219
rect 13857 -8059 13866 -7219
rect 13866 -8059 13900 -7219
rect 13900 -8059 13909 -7219
rect 14005 -8059 14014 -7219
rect 14014 -8059 14048 -7219
rect 14048 -8059 14057 -7219
rect 14153 -8059 14162 -7219
rect 14162 -8059 14196 -7219
rect 14196 -8059 14205 -7219
rect 14301 -8059 14310 -7219
rect 14310 -8059 14344 -7219
rect 14344 -8059 14353 -7219
rect 14449 -8059 14458 -7219
rect 14458 -8059 14492 -7219
rect 14492 -8059 14501 -7219
rect 14597 -8059 14606 -7219
rect 14606 -8059 14640 -7219
rect 14640 -8059 14649 -7219
rect 14745 -8059 14754 -7219
rect 14754 -8059 14788 -7219
rect 14788 -8059 14797 -7219
rect 14893 -8059 14902 -7219
rect 14902 -8059 14936 -7219
rect 14936 -8059 14945 -7219
rect 15041 -8059 15050 -7219
rect 15050 -8059 15084 -7219
rect 15084 -8059 15093 -7219
rect 15189 -8059 15198 -7219
rect 15198 -8059 15232 -7219
rect 15232 -8059 15241 -7219
rect 15337 -8059 15346 -7219
rect 15346 -8059 15380 -7219
rect 15380 -8059 15389 -7219
rect 15485 -8059 15494 -7219
rect 15494 -8059 15528 -7219
rect 15528 -8059 15537 -7219
rect 15633 -8059 15642 -7219
rect 15642 -8059 15676 -7219
rect 15676 -8059 15685 -7219
rect 15781 -8059 15790 -7219
rect 15790 -8059 15824 -7219
rect 15824 -8059 15833 -7219
rect 15929 -8059 15938 -7219
rect 15938 -8059 15972 -7219
rect 15972 -8059 15981 -7219
rect 16077 -8059 16086 -7219
rect 16086 -8059 16120 -7219
rect 16120 -8059 16129 -7219
rect 16225 -8059 16234 -7219
rect 16234 -8059 16268 -7219
rect 16268 -8059 16277 -7219
rect 16373 -8059 16382 -7219
rect 16382 -8059 16416 -7219
rect 16416 -8059 16425 -7219
rect 16521 -8059 16530 -7219
rect 16530 -8059 16564 -7219
rect 16564 -8059 16573 -7219
rect 16669 -8059 16678 -7219
rect 16678 -8059 16712 -7219
rect 16712 -8059 16721 -7219
rect 16817 -8059 16826 -7219
rect 16826 -8059 16860 -7219
rect 16860 -8059 16869 -7219
rect 16965 -8059 16974 -7219
rect 16974 -8059 17008 -7219
rect 17008 -8059 17017 -7219
rect 17113 -8059 17122 -7219
rect 17122 -8059 17156 -7219
rect 17156 -8059 17165 -7219
rect 17261 -8059 17270 -7219
rect 17270 -8059 17304 -7219
rect 17304 -8059 17313 -7219
rect 17409 -8059 17418 -7219
rect 17418 -8059 17452 -7219
rect 17452 -8059 17461 -7219
rect 17557 -8059 17566 -7219
rect 17566 -8059 17600 -7219
rect 17600 -8059 17609 -7219
rect 17705 -8059 17714 -7219
rect 17714 -8059 17748 -7219
rect 17748 -8059 17757 -7219
rect 17853 -8059 17862 -7219
rect 17862 -8059 17896 -7219
rect 17896 -8059 17905 -7219
rect 18001 -8059 18010 -7219
rect 18010 -8059 18044 -7219
rect 18044 -8059 18053 -7219
rect 18149 -8059 18158 -7219
rect 18158 -8059 18192 -7219
rect 18192 -8059 18201 -7219
rect 18297 -8059 18306 -7219
rect 18306 -8059 18340 -7219
rect 18340 -8059 18349 -7219
rect 18445 -8059 18454 -7219
rect 18454 -8059 18488 -7219
rect 18488 -8059 18497 -7219
rect 18593 -8059 18602 -7219
rect 18602 -8059 18636 -7219
rect 18636 -8059 18645 -7219
rect 18741 -8059 18750 -7219
rect 18750 -8059 18784 -7219
rect 18784 -8059 18793 -7219
rect 18889 -8059 18898 -7219
rect 18898 -8059 18932 -7219
rect 18932 -8059 18941 -7219
rect 19037 -8059 19046 -7219
rect 19046 -8059 19080 -7219
rect 19080 -8059 19089 -7219
rect 19185 -8059 19194 -7219
rect 19194 -8059 19228 -7219
rect 19228 -8059 19237 -7219
rect 19333 -8059 19342 -7219
rect 19342 -8059 19376 -7219
rect 19376 -8059 19385 -7219
rect 19481 -8059 19490 -7219
rect 19490 -8059 19524 -7219
rect 19524 -8059 19533 -7219
rect 19629 -8059 19638 -7219
rect 19638 -8059 19672 -7219
rect 19672 -8059 19681 -7219
rect 19777 -8059 19786 -7219
rect 19786 -8059 19820 -7219
rect 19820 -8059 19829 -7219
rect 19925 -8059 19934 -7219
rect 19934 -8059 19968 -7219
rect 19968 -8059 19977 -7219
rect 20073 -8059 20082 -7219
rect 20082 -8059 20116 -7219
rect 20116 -8059 20125 -7219
rect 20221 -8059 20230 -7219
rect 20230 -8059 20264 -7219
rect 20264 -8059 20273 -7219
rect 20369 -8059 20378 -7219
rect 20378 -8059 20412 -7219
rect 20412 -8059 20421 -7219
rect 20517 -8059 20526 -7219
rect 20526 -8059 20560 -7219
rect 20560 -8059 20569 -7219
rect 20665 -8059 20674 -7219
rect 20674 -8059 20708 -7219
rect 20708 -8059 20717 -7219
rect 20813 -8059 20822 -7219
rect 20822 -8059 20856 -7219
rect 20856 -8059 20865 -7219
rect 20961 -8059 20970 -7219
rect 20970 -8059 21004 -7219
rect 21004 -8059 21013 -7219
rect 21109 -8059 21118 -7219
rect 21118 -8059 21152 -7219
rect 21152 -8059 21161 -7219
rect 21257 -8059 21266 -7219
rect 21266 -8059 21300 -7219
rect 21300 -8059 21309 -7219
rect 21405 -8059 21414 -7219
rect 21414 -8059 21448 -7219
rect 21448 -8059 21457 -7219
rect 21553 -8059 21562 -7219
rect 21562 -8059 21596 -7219
rect 21596 -8059 21605 -7219
rect 21701 -8059 21710 -7219
rect 21710 -8059 21744 -7219
rect 21744 -8059 21753 -7219
rect 21849 -8059 21858 -7219
rect 21858 -8059 21892 -7219
rect 21892 -8059 21901 -7219
rect 21997 -8059 22006 -7219
rect 22006 -8059 22040 -7219
rect 22040 -8059 22049 -7219
rect 22145 -8059 22154 -7219
rect 22154 -8059 22188 -7219
rect 22188 -8059 22197 -7219
rect 22293 -8059 22302 -7219
rect 22302 -8059 22336 -7219
rect 22336 -8059 22345 -7219
rect 22441 -8059 22450 -7219
rect 22450 -8059 22484 -7219
rect 22484 -8059 22493 -7219
rect 22589 -8059 22598 -7219
rect 22598 -8059 22632 -7219
rect 22632 -8059 22641 -7219
rect 22737 -8059 22746 -7219
rect 22746 -8059 22780 -7219
rect 22780 -8059 22789 -7219
rect 22885 -8059 22894 -7219
rect 22894 -8059 22928 -7219
rect 22928 -8059 22937 -7219
rect 23033 -8059 23042 -7219
rect 23042 -8059 23076 -7219
rect 23076 -8059 23085 -7219
rect 23181 -8059 23190 -7219
rect 23190 -8059 23224 -7219
rect 23224 -8059 23233 -7219
rect 23329 -8059 23338 -7219
rect 23338 -8059 23372 -7219
rect 23372 -8059 23381 -7219
rect 23477 -8059 23529 -7219
rect 23625 -8059 23634 -7219
rect 23634 -8059 23668 -7219
rect 23668 -8059 23677 -7219
rect 12580 -8289 12670 -8135
rect 12728 -8141 12818 -8135
rect 12728 -8175 12744 -8141
rect 12744 -8175 12802 -8141
rect 12802 -8175 12818 -8141
rect 12728 -8249 12818 -8175
rect 12728 -8283 12744 -8249
rect 12744 -8283 12802 -8249
rect 12802 -8283 12818 -8249
rect 12728 -8289 12818 -8283
rect 12876 -8141 12966 -8135
rect 12876 -8175 12892 -8141
rect 12892 -8175 12950 -8141
rect 12950 -8175 12966 -8141
rect 12876 -8249 12966 -8175
rect 12876 -8283 12892 -8249
rect 12892 -8283 12950 -8249
rect 12950 -8283 12966 -8249
rect 12876 -8289 12966 -8283
rect 13024 -8141 13114 -8135
rect 13024 -8175 13040 -8141
rect 13040 -8175 13098 -8141
rect 13098 -8175 13114 -8141
rect 13024 -8249 13114 -8175
rect 13024 -8283 13040 -8249
rect 13040 -8283 13098 -8249
rect 13098 -8283 13114 -8249
rect 13024 -8289 13114 -8283
rect 13172 -8141 13262 -8135
rect 13172 -8175 13188 -8141
rect 13188 -8175 13246 -8141
rect 13246 -8175 13262 -8141
rect 13172 -8249 13262 -8175
rect 13172 -8283 13188 -8249
rect 13188 -8283 13246 -8249
rect 13246 -8283 13262 -8249
rect 13172 -8289 13262 -8283
rect 13320 -8141 13410 -8135
rect 13320 -8175 13336 -8141
rect 13336 -8175 13394 -8141
rect 13394 -8175 13410 -8141
rect 13320 -8249 13410 -8175
rect 13320 -8283 13336 -8249
rect 13336 -8283 13394 -8249
rect 13394 -8283 13410 -8249
rect 13320 -8289 13410 -8283
rect 13468 -8141 13558 -8135
rect 13468 -8175 13484 -8141
rect 13484 -8175 13542 -8141
rect 13542 -8175 13558 -8141
rect 13468 -8249 13558 -8175
rect 13468 -8283 13484 -8249
rect 13484 -8283 13542 -8249
rect 13542 -8283 13558 -8249
rect 13468 -8289 13558 -8283
rect 13616 -8141 13706 -8135
rect 13616 -8175 13632 -8141
rect 13632 -8175 13690 -8141
rect 13690 -8175 13706 -8141
rect 13616 -8249 13706 -8175
rect 13616 -8283 13632 -8249
rect 13632 -8283 13690 -8249
rect 13690 -8283 13706 -8249
rect 13616 -8289 13706 -8283
rect 13764 -8141 13854 -8135
rect 13764 -8175 13780 -8141
rect 13780 -8175 13838 -8141
rect 13838 -8175 13854 -8141
rect 13764 -8249 13854 -8175
rect 13764 -8283 13780 -8249
rect 13780 -8283 13838 -8249
rect 13838 -8283 13854 -8249
rect 13764 -8289 13854 -8283
rect 13912 -8141 14002 -8135
rect 13912 -8175 13928 -8141
rect 13928 -8175 13986 -8141
rect 13986 -8175 14002 -8141
rect 13912 -8249 14002 -8175
rect 13912 -8283 13928 -8249
rect 13928 -8283 13986 -8249
rect 13986 -8283 14002 -8249
rect 13912 -8289 14002 -8283
rect 14060 -8141 14150 -8135
rect 14060 -8175 14076 -8141
rect 14076 -8175 14134 -8141
rect 14134 -8175 14150 -8141
rect 14060 -8249 14150 -8175
rect 14060 -8283 14076 -8249
rect 14076 -8283 14134 -8249
rect 14134 -8283 14150 -8249
rect 14060 -8289 14150 -8283
rect 14208 -8141 14298 -8135
rect 14208 -8175 14224 -8141
rect 14224 -8175 14282 -8141
rect 14282 -8175 14298 -8141
rect 14208 -8249 14298 -8175
rect 14208 -8283 14224 -8249
rect 14224 -8283 14282 -8249
rect 14282 -8283 14298 -8249
rect 14208 -8289 14298 -8283
rect 14356 -8141 14446 -8135
rect 14356 -8175 14372 -8141
rect 14372 -8175 14430 -8141
rect 14430 -8175 14446 -8141
rect 14356 -8249 14446 -8175
rect 14356 -8283 14372 -8249
rect 14372 -8283 14430 -8249
rect 14430 -8283 14446 -8249
rect 14356 -8289 14446 -8283
rect 14504 -8141 14594 -8135
rect 14504 -8175 14520 -8141
rect 14520 -8175 14578 -8141
rect 14578 -8175 14594 -8141
rect 14504 -8249 14594 -8175
rect 14504 -8283 14520 -8249
rect 14520 -8283 14578 -8249
rect 14578 -8283 14594 -8249
rect 14504 -8289 14594 -8283
rect 14652 -8141 14742 -8135
rect 14652 -8175 14668 -8141
rect 14668 -8175 14726 -8141
rect 14726 -8175 14742 -8141
rect 14652 -8249 14742 -8175
rect 14652 -8283 14668 -8249
rect 14668 -8283 14726 -8249
rect 14726 -8283 14742 -8249
rect 14652 -8289 14742 -8283
rect 14800 -8141 14890 -8135
rect 14800 -8175 14816 -8141
rect 14816 -8175 14874 -8141
rect 14874 -8175 14890 -8141
rect 14800 -8249 14890 -8175
rect 14800 -8283 14816 -8249
rect 14816 -8283 14874 -8249
rect 14874 -8283 14890 -8249
rect 14800 -8289 14890 -8283
rect 14948 -8141 15038 -8135
rect 14948 -8175 14964 -8141
rect 14964 -8175 15022 -8141
rect 15022 -8175 15038 -8141
rect 14948 -8249 15038 -8175
rect 14948 -8283 14964 -8249
rect 14964 -8283 15022 -8249
rect 15022 -8283 15038 -8249
rect 14948 -8289 15038 -8283
rect 15096 -8141 15186 -8135
rect 15096 -8175 15112 -8141
rect 15112 -8175 15170 -8141
rect 15170 -8175 15186 -8141
rect 15096 -8249 15186 -8175
rect 15096 -8283 15112 -8249
rect 15112 -8283 15170 -8249
rect 15170 -8283 15186 -8249
rect 15096 -8289 15186 -8283
rect 15244 -8141 15334 -8135
rect 15244 -8175 15260 -8141
rect 15260 -8175 15318 -8141
rect 15318 -8175 15334 -8141
rect 15244 -8249 15334 -8175
rect 15244 -8283 15260 -8249
rect 15260 -8283 15318 -8249
rect 15318 -8283 15334 -8249
rect 15244 -8289 15334 -8283
rect 15392 -8141 15482 -8135
rect 15392 -8175 15408 -8141
rect 15408 -8175 15466 -8141
rect 15466 -8175 15482 -8141
rect 15392 -8249 15482 -8175
rect 15392 -8283 15408 -8249
rect 15408 -8283 15466 -8249
rect 15466 -8283 15482 -8249
rect 15392 -8289 15482 -8283
rect 15540 -8141 15630 -8135
rect 15540 -8175 15556 -8141
rect 15556 -8175 15614 -8141
rect 15614 -8175 15630 -8141
rect 15540 -8249 15630 -8175
rect 15540 -8283 15556 -8249
rect 15556 -8283 15614 -8249
rect 15614 -8283 15630 -8249
rect 15540 -8289 15630 -8283
rect 15688 -8141 15778 -8135
rect 15688 -8175 15704 -8141
rect 15704 -8175 15762 -8141
rect 15762 -8175 15778 -8141
rect 15688 -8249 15778 -8175
rect 15688 -8283 15704 -8249
rect 15704 -8283 15762 -8249
rect 15762 -8283 15778 -8249
rect 15688 -8289 15778 -8283
rect 15836 -8141 15926 -8135
rect 15836 -8175 15852 -8141
rect 15852 -8175 15910 -8141
rect 15910 -8175 15926 -8141
rect 15836 -8249 15926 -8175
rect 15836 -8283 15852 -8249
rect 15852 -8283 15910 -8249
rect 15910 -8283 15926 -8249
rect 15836 -8289 15926 -8283
rect 15984 -8141 16074 -8135
rect 15984 -8175 16000 -8141
rect 16000 -8175 16058 -8141
rect 16058 -8175 16074 -8141
rect 15984 -8249 16074 -8175
rect 15984 -8283 16000 -8249
rect 16000 -8283 16058 -8249
rect 16058 -8283 16074 -8249
rect 15984 -8289 16074 -8283
rect 16132 -8141 16222 -8135
rect 16132 -8175 16148 -8141
rect 16148 -8175 16206 -8141
rect 16206 -8175 16222 -8141
rect 16132 -8249 16222 -8175
rect 16132 -8283 16148 -8249
rect 16148 -8283 16206 -8249
rect 16206 -8283 16222 -8249
rect 16132 -8289 16222 -8283
rect 16280 -8141 16370 -8135
rect 16280 -8175 16296 -8141
rect 16296 -8175 16354 -8141
rect 16354 -8175 16370 -8141
rect 16280 -8249 16370 -8175
rect 16280 -8283 16296 -8249
rect 16296 -8283 16354 -8249
rect 16354 -8283 16370 -8249
rect 16280 -8289 16370 -8283
rect 16428 -8141 16518 -8135
rect 16428 -8175 16444 -8141
rect 16444 -8175 16502 -8141
rect 16502 -8175 16518 -8141
rect 16428 -8249 16518 -8175
rect 16428 -8283 16444 -8249
rect 16444 -8283 16502 -8249
rect 16502 -8283 16518 -8249
rect 16428 -8289 16518 -8283
rect 16576 -8141 16666 -8135
rect 16576 -8175 16592 -8141
rect 16592 -8175 16650 -8141
rect 16650 -8175 16666 -8141
rect 16576 -8249 16666 -8175
rect 16576 -8283 16592 -8249
rect 16592 -8283 16650 -8249
rect 16650 -8283 16666 -8249
rect 16576 -8289 16666 -8283
rect 16724 -8141 16814 -8135
rect 16724 -8175 16740 -8141
rect 16740 -8175 16798 -8141
rect 16798 -8175 16814 -8141
rect 16724 -8249 16814 -8175
rect 16724 -8283 16740 -8249
rect 16740 -8283 16798 -8249
rect 16798 -8283 16814 -8249
rect 16724 -8289 16814 -8283
rect 16872 -8141 16962 -8135
rect 16872 -8175 16888 -8141
rect 16888 -8175 16946 -8141
rect 16946 -8175 16962 -8141
rect 16872 -8249 16962 -8175
rect 16872 -8283 16888 -8249
rect 16888 -8283 16946 -8249
rect 16946 -8283 16962 -8249
rect 16872 -8289 16962 -8283
rect 17020 -8141 17110 -8135
rect 17020 -8175 17036 -8141
rect 17036 -8175 17094 -8141
rect 17094 -8175 17110 -8141
rect 17020 -8249 17110 -8175
rect 17020 -8283 17036 -8249
rect 17036 -8283 17094 -8249
rect 17094 -8283 17110 -8249
rect 17020 -8289 17110 -8283
rect 17168 -8141 17258 -8135
rect 17168 -8175 17184 -8141
rect 17184 -8175 17242 -8141
rect 17242 -8175 17258 -8141
rect 17168 -8249 17258 -8175
rect 17168 -8283 17184 -8249
rect 17184 -8283 17242 -8249
rect 17242 -8283 17258 -8249
rect 17168 -8289 17258 -8283
rect 17316 -8141 17406 -8135
rect 17316 -8175 17332 -8141
rect 17332 -8175 17390 -8141
rect 17390 -8175 17406 -8141
rect 17316 -8249 17406 -8175
rect 17316 -8283 17332 -8249
rect 17332 -8283 17390 -8249
rect 17390 -8283 17406 -8249
rect 17316 -8289 17406 -8283
rect 17464 -8141 17554 -8135
rect 17464 -8175 17480 -8141
rect 17480 -8175 17538 -8141
rect 17538 -8175 17554 -8141
rect 17464 -8249 17554 -8175
rect 17464 -8283 17480 -8249
rect 17480 -8283 17538 -8249
rect 17538 -8283 17554 -8249
rect 17464 -8289 17554 -8283
rect 17612 -8141 17702 -8135
rect 17612 -8175 17628 -8141
rect 17628 -8175 17686 -8141
rect 17686 -8175 17702 -8141
rect 17612 -8249 17702 -8175
rect 17612 -8283 17628 -8249
rect 17628 -8283 17686 -8249
rect 17686 -8283 17702 -8249
rect 17612 -8289 17702 -8283
rect 17760 -8141 17850 -8135
rect 17760 -8175 17776 -8141
rect 17776 -8175 17834 -8141
rect 17834 -8175 17850 -8141
rect 17760 -8249 17850 -8175
rect 17760 -8283 17776 -8249
rect 17776 -8283 17834 -8249
rect 17834 -8283 17850 -8249
rect 17760 -8289 17850 -8283
rect 17908 -8141 17998 -8135
rect 17908 -8175 17924 -8141
rect 17924 -8175 17982 -8141
rect 17982 -8175 17998 -8141
rect 17908 -8249 17998 -8175
rect 17908 -8283 17924 -8249
rect 17924 -8283 17982 -8249
rect 17982 -8283 17998 -8249
rect 17908 -8289 17998 -8283
rect 18056 -8141 18146 -8135
rect 18056 -8175 18072 -8141
rect 18072 -8175 18130 -8141
rect 18130 -8175 18146 -8141
rect 18056 -8249 18146 -8175
rect 18056 -8283 18072 -8249
rect 18072 -8283 18130 -8249
rect 18130 -8283 18146 -8249
rect 18056 -8289 18146 -8283
rect 18204 -8141 18294 -8135
rect 18204 -8175 18220 -8141
rect 18220 -8175 18278 -8141
rect 18278 -8175 18294 -8141
rect 18204 -8249 18294 -8175
rect 18204 -8283 18220 -8249
rect 18220 -8283 18278 -8249
rect 18278 -8283 18294 -8249
rect 18204 -8289 18294 -8283
rect 18352 -8141 18442 -8135
rect 18352 -8175 18368 -8141
rect 18368 -8175 18426 -8141
rect 18426 -8175 18442 -8141
rect 18352 -8249 18442 -8175
rect 18352 -8283 18368 -8249
rect 18368 -8283 18426 -8249
rect 18426 -8283 18442 -8249
rect 18352 -8289 18442 -8283
rect 18500 -8141 18590 -8135
rect 18500 -8175 18516 -8141
rect 18516 -8175 18574 -8141
rect 18574 -8175 18590 -8141
rect 18500 -8249 18590 -8175
rect 18500 -8283 18516 -8249
rect 18516 -8283 18574 -8249
rect 18574 -8283 18590 -8249
rect 18500 -8289 18590 -8283
rect 18648 -8141 18738 -8135
rect 18648 -8175 18664 -8141
rect 18664 -8175 18722 -8141
rect 18722 -8175 18738 -8141
rect 18648 -8249 18738 -8175
rect 18648 -8283 18664 -8249
rect 18664 -8283 18722 -8249
rect 18722 -8283 18738 -8249
rect 18648 -8289 18738 -8283
rect 18796 -8141 18886 -8135
rect 18796 -8175 18812 -8141
rect 18812 -8175 18870 -8141
rect 18870 -8175 18886 -8141
rect 18796 -8249 18886 -8175
rect 18796 -8283 18812 -8249
rect 18812 -8283 18870 -8249
rect 18870 -8283 18886 -8249
rect 18796 -8289 18886 -8283
rect 18944 -8141 19034 -8135
rect 18944 -8175 18960 -8141
rect 18960 -8175 19018 -8141
rect 19018 -8175 19034 -8141
rect 18944 -8249 19034 -8175
rect 18944 -8283 18960 -8249
rect 18960 -8283 19018 -8249
rect 19018 -8283 19034 -8249
rect 18944 -8289 19034 -8283
rect 19092 -8141 19182 -8135
rect 19092 -8175 19108 -8141
rect 19108 -8175 19166 -8141
rect 19166 -8175 19182 -8141
rect 19092 -8249 19182 -8175
rect 19092 -8283 19108 -8249
rect 19108 -8283 19166 -8249
rect 19166 -8283 19182 -8249
rect 19092 -8289 19182 -8283
rect 19240 -8141 19330 -8135
rect 19240 -8175 19256 -8141
rect 19256 -8175 19314 -8141
rect 19314 -8175 19330 -8141
rect 19240 -8249 19330 -8175
rect 19240 -8283 19256 -8249
rect 19256 -8283 19314 -8249
rect 19314 -8283 19330 -8249
rect 19240 -8289 19330 -8283
rect 19388 -8141 19478 -8135
rect 19388 -8175 19404 -8141
rect 19404 -8175 19462 -8141
rect 19462 -8175 19478 -8141
rect 19388 -8249 19478 -8175
rect 19388 -8283 19404 -8249
rect 19404 -8283 19462 -8249
rect 19462 -8283 19478 -8249
rect 19388 -8289 19478 -8283
rect 19536 -8141 19626 -8135
rect 19536 -8175 19552 -8141
rect 19552 -8175 19610 -8141
rect 19610 -8175 19626 -8141
rect 19536 -8249 19626 -8175
rect 19536 -8283 19552 -8249
rect 19552 -8283 19610 -8249
rect 19610 -8283 19626 -8249
rect 19536 -8289 19626 -8283
rect 19684 -8141 19774 -8135
rect 19684 -8175 19700 -8141
rect 19700 -8175 19758 -8141
rect 19758 -8175 19774 -8141
rect 19684 -8249 19774 -8175
rect 19684 -8283 19700 -8249
rect 19700 -8283 19758 -8249
rect 19758 -8283 19774 -8249
rect 19684 -8289 19774 -8283
rect 19832 -8141 19922 -8135
rect 19832 -8175 19848 -8141
rect 19848 -8175 19906 -8141
rect 19906 -8175 19922 -8141
rect 19832 -8249 19922 -8175
rect 19832 -8283 19848 -8249
rect 19848 -8283 19906 -8249
rect 19906 -8283 19922 -8249
rect 19832 -8289 19922 -8283
rect 19980 -8141 20070 -8135
rect 19980 -8175 19996 -8141
rect 19996 -8175 20054 -8141
rect 20054 -8175 20070 -8141
rect 19980 -8249 20070 -8175
rect 19980 -8283 19996 -8249
rect 19996 -8283 20054 -8249
rect 20054 -8283 20070 -8249
rect 19980 -8289 20070 -8283
rect 20128 -8141 20218 -8135
rect 20128 -8175 20144 -8141
rect 20144 -8175 20202 -8141
rect 20202 -8175 20218 -8141
rect 20128 -8249 20218 -8175
rect 20128 -8283 20144 -8249
rect 20144 -8283 20202 -8249
rect 20202 -8283 20218 -8249
rect 20128 -8289 20218 -8283
rect 20276 -8141 20366 -8135
rect 20276 -8175 20292 -8141
rect 20292 -8175 20350 -8141
rect 20350 -8175 20366 -8141
rect 20276 -8249 20366 -8175
rect 20276 -8283 20292 -8249
rect 20292 -8283 20350 -8249
rect 20350 -8283 20366 -8249
rect 20276 -8289 20366 -8283
rect 20424 -8141 20514 -8135
rect 20424 -8175 20440 -8141
rect 20440 -8175 20498 -8141
rect 20498 -8175 20514 -8141
rect 20424 -8249 20514 -8175
rect 20424 -8283 20440 -8249
rect 20440 -8283 20498 -8249
rect 20498 -8283 20514 -8249
rect 20424 -8289 20514 -8283
rect 20572 -8141 20662 -8135
rect 20572 -8175 20588 -8141
rect 20588 -8175 20646 -8141
rect 20646 -8175 20662 -8141
rect 20572 -8249 20662 -8175
rect 20572 -8283 20588 -8249
rect 20588 -8283 20646 -8249
rect 20646 -8283 20662 -8249
rect 20572 -8289 20662 -8283
rect 20720 -8141 20810 -8135
rect 20720 -8175 20736 -8141
rect 20736 -8175 20794 -8141
rect 20794 -8175 20810 -8141
rect 20720 -8249 20810 -8175
rect 20720 -8283 20736 -8249
rect 20736 -8283 20794 -8249
rect 20794 -8283 20810 -8249
rect 20720 -8289 20810 -8283
rect 20868 -8141 20958 -8135
rect 20868 -8175 20884 -8141
rect 20884 -8175 20942 -8141
rect 20942 -8175 20958 -8141
rect 20868 -8249 20958 -8175
rect 20868 -8283 20884 -8249
rect 20884 -8283 20942 -8249
rect 20942 -8283 20958 -8249
rect 20868 -8289 20958 -8283
rect 21016 -8141 21106 -8135
rect 21016 -8175 21032 -8141
rect 21032 -8175 21090 -8141
rect 21090 -8175 21106 -8141
rect 21016 -8249 21106 -8175
rect 21016 -8283 21032 -8249
rect 21032 -8283 21090 -8249
rect 21090 -8283 21106 -8249
rect 21016 -8289 21106 -8283
rect 21164 -8141 21254 -8135
rect 21164 -8175 21180 -8141
rect 21180 -8175 21238 -8141
rect 21238 -8175 21254 -8141
rect 21164 -8249 21254 -8175
rect 21164 -8283 21180 -8249
rect 21180 -8283 21238 -8249
rect 21238 -8283 21254 -8249
rect 21164 -8289 21254 -8283
rect 21312 -8141 21402 -8135
rect 21312 -8175 21328 -8141
rect 21328 -8175 21386 -8141
rect 21386 -8175 21402 -8141
rect 21312 -8249 21402 -8175
rect 21312 -8283 21328 -8249
rect 21328 -8283 21386 -8249
rect 21386 -8283 21402 -8249
rect 21312 -8289 21402 -8283
rect 21460 -8141 21550 -8135
rect 21460 -8175 21476 -8141
rect 21476 -8175 21534 -8141
rect 21534 -8175 21550 -8141
rect 21460 -8249 21550 -8175
rect 21460 -8283 21476 -8249
rect 21476 -8283 21534 -8249
rect 21534 -8283 21550 -8249
rect 21460 -8289 21550 -8283
rect 21608 -8141 21698 -8135
rect 21608 -8175 21624 -8141
rect 21624 -8175 21682 -8141
rect 21682 -8175 21698 -8141
rect 21608 -8249 21698 -8175
rect 21608 -8283 21624 -8249
rect 21624 -8283 21682 -8249
rect 21682 -8283 21698 -8249
rect 21608 -8289 21698 -8283
rect 21756 -8141 21846 -8135
rect 21756 -8175 21772 -8141
rect 21772 -8175 21830 -8141
rect 21830 -8175 21846 -8141
rect 21756 -8249 21846 -8175
rect 21756 -8283 21772 -8249
rect 21772 -8283 21830 -8249
rect 21830 -8283 21846 -8249
rect 21756 -8289 21846 -8283
rect 21904 -8141 21994 -8135
rect 21904 -8175 21920 -8141
rect 21920 -8175 21978 -8141
rect 21978 -8175 21994 -8141
rect 21904 -8249 21994 -8175
rect 21904 -8283 21920 -8249
rect 21920 -8283 21978 -8249
rect 21978 -8283 21994 -8249
rect 21904 -8289 21994 -8283
rect 22052 -8141 22142 -8135
rect 22052 -8175 22068 -8141
rect 22068 -8175 22126 -8141
rect 22126 -8175 22142 -8141
rect 22052 -8249 22142 -8175
rect 22052 -8283 22068 -8249
rect 22068 -8283 22126 -8249
rect 22126 -8283 22142 -8249
rect 22052 -8289 22142 -8283
rect 22200 -8141 22290 -8135
rect 22200 -8175 22216 -8141
rect 22216 -8175 22274 -8141
rect 22274 -8175 22290 -8141
rect 22200 -8249 22290 -8175
rect 22200 -8283 22216 -8249
rect 22216 -8283 22274 -8249
rect 22274 -8283 22290 -8249
rect 22200 -8289 22290 -8283
rect 22348 -8141 22438 -8135
rect 22348 -8175 22364 -8141
rect 22364 -8175 22422 -8141
rect 22422 -8175 22438 -8141
rect 22348 -8249 22438 -8175
rect 22348 -8283 22364 -8249
rect 22364 -8283 22422 -8249
rect 22422 -8283 22438 -8249
rect 22348 -8289 22438 -8283
rect 22496 -8141 22586 -8135
rect 22496 -8175 22512 -8141
rect 22512 -8175 22570 -8141
rect 22570 -8175 22586 -8141
rect 22496 -8249 22586 -8175
rect 22496 -8283 22512 -8249
rect 22512 -8283 22570 -8249
rect 22570 -8283 22586 -8249
rect 22496 -8289 22586 -8283
rect 22644 -8141 22734 -8135
rect 22644 -8175 22660 -8141
rect 22660 -8175 22718 -8141
rect 22718 -8175 22734 -8141
rect 22644 -8249 22734 -8175
rect 22644 -8283 22660 -8249
rect 22660 -8283 22718 -8249
rect 22718 -8283 22734 -8249
rect 22644 -8289 22734 -8283
rect 22792 -8141 22882 -8135
rect 22792 -8175 22808 -8141
rect 22808 -8175 22866 -8141
rect 22866 -8175 22882 -8141
rect 22792 -8249 22882 -8175
rect 22792 -8283 22808 -8249
rect 22808 -8283 22866 -8249
rect 22866 -8283 22882 -8249
rect 22792 -8289 22882 -8283
rect 22940 -8141 23030 -8135
rect 22940 -8175 22956 -8141
rect 22956 -8175 23014 -8141
rect 23014 -8175 23030 -8141
rect 22940 -8249 23030 -8175
rect 22940 -8283 22956 -8249
rect 22956 -8283 23014 -8249
rect 23014 -8283 23030 -8249
rect 22940 -8289 23030 -8283
rect 23088 -8141 23178 -8135
rect 23088 -8175 23104 -8141
rect 23104 -8175 23162 -8141
rect 23162 -8175 23178 -8141
rect 23088 -8249 23178 -8175
rect 23088 -8283 23104 -8249
rect 23104 -8283 23162 -8249
rect 23162 -8283 23178 -8249
rect 23088 -8289 23178 -8283
rect 23236 -8141 23326 -8135
rect 23236 -8175 23252 -8141
rect 23252 -8175 23310 -8141
rect 23310 -8175 23326 -8141
rect 23236 -8249 23326 -8175
rect 23236 -8283 23252 -8249
rect 23252 -8283 23310 -8249
rect 23310 -8283 23326 -8249
rect 23236 -8289 23326 -8283
rect 23384 -8141 23474 -8135
rect 23384 -8175 23400 -8141
rect 23400 -8175 23458 -8141
rect 23458 -8175 23474 -8141
rect 23384 -8249 23474 -8175
rect 23384 -8283 23400 -8249
rect 23400 -8283 23458 -8249
rect 23458 -8283 23474 -8249
rect 23384 -8289 23474 -8283
rect 23532 -8141 23622 -8135
rect 23532 -8175 23548 -8141
rect 23548 -8175 23606 -8141
rect 23606 -8175 23622 -8141
rect 23532 -8249 23622 -8175
rect 23532 -8283 23548 -8249
rect 23548 -8283 23606 -8249
rect 23606 -8283 23622 -8249
rect 23532 -8289 23622 -8283
rect 9839 -8555 9868 -8538
rect 9868 -8555 9891 -8538
rect 9919 -8555 9940 -8538
rect 9940 -8555 9971 -8538
rect 9999 -8555 10012 -8538
rect 10012 -8555 10050 -8538
rect 10050 -8555 10051 -8538
rect 10079 -8555 10084 -8538
rect 10084 -8555 10122 -8538
rect 10122 -8555 10131 -8538
rect 10159 -8555 10194 -8538
rect 10194 -8555 10211 -8538
rect 10239 -8555 10266 -8538
rect 10266 -8555 10291 -8538
rect 10319 -8555 10338 -8538
rect 10338 -8555 10371 -8538
rect 10399 -8555 10410 -8538
rect 10410 -8555 10444 -8538
rect 10444 -8555 10451 -8538
rect 9839 -8590 9891 -8555
rect 9919 -8590 9971 -8555
rect 9999 -8590 10051 -8555
rect 10079 -8590 10131 -8555
rect 10159 -8590 10211 -8555
rect 10239 -8590 10291 -8555
rect 10319 -8590 10371 -8555
rect 10399 -8590 10451 -8555
rect 10479 -8555 10482 -8538
rect 10482 -8555 10516 -8538
rect 10516 -8555 10531 -8538
rect 10559 -8555 10588 -8538
rect 10588 -8555 10611 -8538
rect 10479 -8590 10531 -8555
rect 10559 -8590 10611 -8555
rect 9839 -8629 9868 -8617
rect 9868 -8629 9891 -8617
rect 9919 -8629 9940 -8617
rect 9940 -8629 9971 -8617
rect 9999 -8629 10012 -8617
rect 10012 -8629 10050 -8617
rect 10050 -8629 10051 -8617
rect 10079 -8629 10084 -8617
rect 10084 -8629 10122 -8617
rect 10122 -8629 10131 -8617
rect 10159 -8629 10194 -8617
rect 10194 -8629 10211 -8617
rect 10239 -8629 10266 -8617
rect 10266 -8629 10291 -8617
rect 10319 -8629 10338 -8617
rect 10338 -8629 10371 -8617
rect 10399 -8629 10410 -8617
rect 10410 -8629 10444 -8617
rect 10444 -8629 10451 -8617
rect 9839 -8669 9891 -8629
rect 9919 -8669 9971 -8629
rect 9999 -8669 10051 -8629
rect 10079 -8669 10131 -8629
rect 10159 -8669 10211 -8629
rect 10239 -8669 10291 -8629
rect 10319 -8669 10371 -8629
rect 10399 -8669 10451 -8629
rect 10479 -8629 10482 -8617
rect 10482 -8629 10516 -8617
rect 10516 -8629 10531 -8617
rect 10559 -8629 10588 -8617
rect 10588 -8629 10611 -8617
rect 10479 -8669 10531 -8629
rect 10559 -8669 10611 -8629
rect 5759 -8881 5811 -8829
rect 5839 -8881 5891 -8829
rect 5919 -8881 5971 -8829
rect 5999 -8881 6051 -8829
rect 6079 -8881 6131 -8829
rect 6159 -8881 6211 -8829
rect 6239 -8881 6291 -8829
rect 6319 -8881 6371 -8829
rect 6399 -8881 6451 -8829
rect 6479 -8881 6531 -8829
rect 6559 -8881 6611 -8829
rect 6639 -8881 6691 -8829
rect 6719 -8881 6771 -8829
rect 6799 -8881 6851 -8829
rect 6879 -8881 6931 -8829
rect 6959 -8881 7011 -8829
rect 7039 -8881 7091 -8829
rect 7119 -8881 7171 -8829
rect 7199 -8881 7251 -8829
rect 7279 -8881 7331 -8829
rect 7359 -8881 7411 -8829
rect 7439 -8881 7491 -8829
rect 7519 -8881 7571 -8829
rect 7599 -8881 7651 -8829
rect 7679 -8881 7731 -8829
rect 7759 -8881 7811 -8829
rect 7839 -8881 7891 -8829
rect 7919 -8881 7971 -8829
rect 7999 -8881 8051 -8829
rect 8079 -8881 8131 -8829
rect 8159 -8881 8211 -8829
rect 8239 -8881 8291 -8829
rect 8319 -8881 8371 -8829
rect 8399 -8881 8451 -8829
rect 8479 -8881 8531 -8829
rect 8559 -8881 8611 -8829
rect 8639 -8881 8691 -8829
rect 8719 -8881 8771 -8829
rect 8799 -8881 8851 -8829
rect 8879 -8881 8931 -8829
rect 8959 -8881 9011 -8829
rect 9039 -8881 9091 -8829
rect 9119 -8881 9171 -8829
rect 9199 -8881 9251 -8829
rect 9279 -8881 9331 -8829
rect 9359 -8881 9411 -8829
rect 9439 -8881 9491 -8829
rect 9519 -8881 9571 -8829
rect 9599 -8881 9651 -8829
rect 9679 -8881 9731 -8829
rect 9759 -8881 9811 -8829
rect 9839 -8881 9891 -8829
rect 9919 -8881 9971 -8829
rect 9999 -8881 10051 -8829
rect 10079 -8881 10131 -8829
rect 10159 -8881 10211 -8829
rect 10239 -8881 10291 -8829
rect 10319 -8881 10371 -8829
rect 10399 -8881 10451 -8829
rect 10479 -8881 10531 -8829
rect 10559 -8881 10611 -8829
rect 10639 -8881 10691 -8829
rect 10719 -8881 10771 -8829
rect 10799 -8881 10851 -8829
rect 5759 -8945 5811 -8909
rect 5759 -8961 5774 -8945
rect 5774 -8961 5808 -8945
rect 5808 -8961 5811 -8945
rect 5839 -8945 5891 -8909
rect 5839 -8961 5846 -8945
rect 5846 -8961 5880 -8945
rect 5880 -8961 5891 -8945
rect 5919 -8945 5971 -8909
rect 5919 -8961 5928 -8945
rect 5928 -8961 5962 -8945
rect 5962 -8961 5971 -8945
rect 5999 -8945 6051 -8909
rect 5999 -8961 6000 -8945
rect 6000 -8961 6034 -8945
rect 6034 -8961 6051 -8945
rect 6079 -8945 6131 -8909
rect 6159 -8945 6211 -8909
rect 6239 -8945 6291 -8909
rect 6319 -8945 6371 -8909
rect 6399 -8945 6451 -8909
rect 6479 -8945 6531 -8909
rect 6559 -8945 6611 -8909
rect 6639 -8945 6691 -8909
rect 6719 -8945 6771 -8909
rect 6799 -8945 6851 -8909
rect 6879 -8945 6931 -8909
rect 6959 -8945 7011 -8909
rect 7039 -8945 7091 -8909
rect 7119 -8945 7171 -8909
rect 7199 -8945 7251 -8909
rect 7279 -8945 7331 -8909
rect 7359 -8945 7411 -8909
rect 7439 -8945 7491 -8909
rect 7519 -8945 7571 -8909
rect 7599 -8945 7651 -8909
rect 7679 -8945 7731 -8909
rect 6079 -8961 6082 -8945
rect 6082 -8961 6116 -8945
rect 6116 -8961 6131 -8945
rect 6159 -8961 6188 -8945
rect 6188 -8961 6211 -8945
rect 6239 -8961 6270 -8945
rect 6270 -8961 6291 -8945
rect 6319 -8961 6342 -8945
rect 6342 -8961 6371 -8945
rect 6399 -8961 6424 -8945
rect 6424 -8961 6451 -8945
rect 6479 -8961 6496 -8945
rect 6496 -8961 6531 -8945
rect 6559 -8961 6578 -8945
rect 6578 -8961 6611 -8945
rect 6639 -8961 6650 -8945
rect 6650 -8961 6691 -8945
rect 6719 -8961 6732 -8945
rect 6732 -8961 6770 -8945
rect 6770 -8961 6771 -8945
rect 6799 -8961 6804 -8945
rect 6804 -8961 6851 -8945
rect 6879 -8961 6886 -8945
rect 6886 -8961 6924 -8945
rect 6924 -8961 6931 -8945
rect 6959 -8961 7006 -8945
rect 7006 -8961 7011 -8945
rect 7039 -8961 7040 -8945
rect 7040 -8961 7078 -8945
rect 7078 -8961 7091 -8945
rect 7119 -8961 7160 -8945
rect 7160 -8961 7171 -8945
rect 7199 -8961 7232 -8945
rect 7232 -8961 7251 -8945
rect 7279 -8961 7314 -8945
rect 7314 -8961 7331 -8945
rect 7359 -8961 7386 -8945
rect 7386 -8961 7411 -8945
rect 7439 -8961 7468 -8945
rect 7468 -8961 7491 -8945
rect 7519 -8961 7540 -8945
rect 7540 -8961 7571 -8945
rect 7599 -8961 7622 -8945
rect 7622 -8961 7651 -8945
rect 7679 -8961 7694 -8945
rect 7694 -8961 7728 -8945
rect 7728 -8961 7731 -8945
rect 7759 -8945 7811 -8909
rect 7759 -8961 7776 -8945
rect 7776 -8961 7810 -8945
rect 7810 -8961 7811 -8945
rect 7839 -8945 7891 -8909
rect 7839 -8961 7848 -8945
rect 7848 -8961 7882 -8945
rect 7882 -8961 7891 -8945
rect 7919 -8945 7971 -8909
rect 7919 -8961 7930 -8945
rect 7930 -8961 7964 -8945
rect 7964 -8961 7971 -8945
rect 7999 -8945 8051 -8909
rect 7999 -8961 8002 -8945
rect 8002 -8961 8036 -8945
rect 8036 -8961 8051 -8945
rect 8079 -8945 8131 -8909
rect 8159 -8945 8211 -8909
rect 8239 -8945 8291 -8909
rect 8319 -8945 8371 -8909
rect 8399 -8945 8451 -8909
rect 8479 -8945 8531 -8909
rect 8559 -8945 8611 -8909
rect 8639 -8945 8691 -8909
rect 8719 -8945 8771 -8909
rect 8799 -8945 8851 -8909
rect 8879 -8945 8931 -8909
rect 8959 -8945 9011 -8909
rect 9039 -8945 9091 -8909
rect 9119 -8945 9171 -8909
rect 9199 -8945 9251 -8909
rect 9279 -8945 9331 -8909
rect 9359 -8945 9411 -8909
rect 9439 -8945 9491 -8909
rect 9519 -8945 9571 -8909
rect 9599 -8945 9651 -8909
rect 9679 -8945 9731 -8909
rect 8079 -8961 8084 -8945
rect 8084 -8961 8118 -8945
rect 8118 -8961 8131 -8945
rect 8159 -8961 8190 -8945
rect 8190 -8961 8211 -8945
rect 8239 -8961 8272 -8945
rect 8272 -8961 8291 -8945
rect 8319 -8961 8344 -8945
rect 8344 -8961 8371 -8945
rect 8399 -8961 8426 -8945
rect 8426 -8961 8451 -8945
rect 8479 -8961 8498 -8945
rect 8498 -8961 8531 -8945
rect 8559 -8961 8580 -8945
rect 8580 -8961 8611 -8945
rect 8639 -8961 8652 -8945
rect 8652 -8961 8691 -8945
rect 8719 -8961 8734 -8945
rect 8734 -8961 8771 -8945
rect 8799 -8961 8806 -8945
rect 8806 -8961 8851 -8945
rect 8879 -8961 8888 -8945
rect 8888 -8961 8926 -8945
rect 8926 -8961 8931 -8945
rect 8959 -8961 8960 -8945
rect 8960 -8961 9008 -8945
rect 9008 -8961 9011 -8945
rect 9039 -8961 9042 -8945
rect 9042 -8961 9080 -8945
rect 9080 -8961 9091 -8945
rect 9119 -8961 9162 -8945
rect 9162 -8961 9171 -8945
rect 9199 -8961 9234 -8945
rect 9234 -8961 9251 -8945
rect 9279 -8961 9316 -8945
rect 9316 -8961 9331 -8945
rect 9359 -8961 9388 -8945
rect 9388 -8961 9411 -8945
rect 9439 -8961 9470 -8945
rect 9470 -8961 9491 -8945
rect 9519 -8961 9542 -8945
rect 9542 -8961 9571 -8945
rect 9599 -8961 9624 -8945
rect 9624 -8961 9651 -8945
rect 9679 -8961 9696 -8945
rect 9696 -8961 9730 -8945
rect 9730 -8961 9731 -8945
rect 9759 -8945 9811 -8909
rect 9839 -8945 9891 -8909
rect 9759 -8961 9778 -8945
rect 9778 -8961 9811 -8945
rect 9839 -8961 9850 -8945
rect 9850 -8961 9884 -8945
rect 9884 -8961 9891 -8945
rect 9919 -8945 9971 -8909
rect 9919 -8961 9932 -8945
rect 9932 -8961 9966 -8945
rect 9966 -8961 9971 -8945
rect 9999 -8945 10051 -8909
rect 9999 -8961 10004 -8945
rect 10004 -8961 10038 -8945
rect 10038 -8961 10051 -8945
rect 10079 -8945 10131 -8909
rect 10159 -8945 10211 -8909
rect 10079 -8961 10086 -8945
rect 10086 -8961 10120 -8945
rect 10120 -8961 10131 -8945
rect 10159 -8961 10192 -8945
rect 10192 -8961 10211 -8945
rect 10239 -8945 10291 -8909
rect 10319 -8945 10371 -8909
rect 10399 -8945 10451 -8909
rect 10479 -8945 10531 -8909
rect 10559 -8945 10611 -8909
rect 10639 -8945 10691 -8909
rect 10719 -8945 10771 -8909
rect 10799 -8945 10851 -8909
rect 10239 -8961 10240 -8945
rect 10240 -8961 10274 -8945
rect 10274 -8961 10291 -8945
rect 10319 -8961 10346 -8945
rect 10346 -8961 10371 -8945
rect 10399 -8961 10428 -8945
rect 10428 -8961 10451 -8945
rect 10479 -8961 10500 -8945
rect 10500 -8961 10531 -8945
rect 10559 -8961 10582 -8945
rect 10582 -8961 10611 -8945
rect 10639 -8961 10654 -8945
rect 10654 -8961 10691 -8945
rect 10719 -8961 10736 -8945
rect 10736 -8961 10771 -8945
rect 10799 -8961 10808 -8945
rect 10808 -8961 10851 -8945
rect 12525 -9205 12534 -8365
rect 12534 -9205 12568 -8365
rect 12568 -9205 12577 -8365
rect 12673 -9205 12682 -8365
rect 12682 -9205 12716 -8365
rect 12716 -9205 12725 -8365
rect 12821 -9205 12830 -8365
rect 12830 -9205 12864 -8365
rect 12864 -9205 12873 -8365
rect 12969 -9205 12978 -8365
rect 12978 -9205 13012 -8365
rect 13012 -9205 13021 -8365
rect 13117 -9205 13126 -8365
rect 13126 -9205 13160 -8365
rect 13160 -9205 13169 -8365
rect 13265 -9205 13274 -8365
rect 13274 -9205 13308 -8365
rect 13308 -9205 13317 -8365
rect 13413 -9205 13422 -8365
rect 13422 -9205 13456 -8365
rect 13456 -9205 13465 -8365
rect 13561 -9205 13570 -8365
rect 13570 -9205 13604 -8365
rect 13604 -9205 13613 -8365
rect 13709 -9205 13718 -8365
rect 13718 -9205 13752 -8365
rect 13752 -9205 13761 -8365
rect 13857 -9205 13866 -8365
rect 13866 -9205 13900 -8365
rect 13900 -9205 13909 -8365
rect 14005 -9205 14014 -8365
rect 14014 -9205 14048 -8365
rect 14048 -9205 14057 -8365
rect 14153 -9205 14162 -8365
rect 14162 -9205 14196 -8365
rect 14196 -9205 14205 -8365
rect 14301 -9205 14310 -8365
rect 14310 -9205 14344 -8365
rect 14344 -9205 14353 -8365
rect 14449 -9205 14458 -8365
rect 14458 -9205 14492 -8365
rect 14492 -9205 14501 -8365
rect 14597 -9205 14606 -8365
rect 14606 -9205 14640 -8365
rect 14640 -9205 14649 -8365
rect 14745 -9205 14754 -8365
rect 14754 -9205 14788 -8365
rect 14788 -9205 14797 -8365
rect 14893 -9205 14902 -8365
rect 14902 -9205 14936 -8365
rect 14936 -9205 14945 -8365
rect 15041 -9205 15050 -8365
rect 15050 -9205 15084 -8365
rect 15084 -9205 15093 -8365
rect 15189 -9205 15198 -8365
rect 15198 -9205 15232 -8365
rect 15232 -9205 15241 -8365
rect 15337 -9205 15346 -8365
rect 15346 -9205 15380 -8365
rect 15380 -9205 15389 -8365
rect 15485 -9205 15494 -8365
rect 15494 -9205 15528 -8365
rect 15528 -9205 15537 -8365
rect 15633 -9205 15642 -8365
rect 15642 -9205 15676 -8365
rect 15676 -9205 15685 -8365
rect 15781 -9205 15790 -8365
rect 15790 -9205 15824 -8365
rect 15824 -9205 15833 -8365
rect 15929 -9205 15938 -8365
rect 15938 -9205 15972 -8365
rect 15972 -9205 15981 -8365
rect 16077 -9205 16086 -8365
rect 16086 -9205 16120 -8365
rect 16120 -9205 16129 -8365
rect 16225 -9205 16234 -8365
rect 16234 -9205 16268 -8365
rect 16268 -9205 16277 -8365
rect 16373 -9205 16382 -8365
rect 16382 -9205 16416 -8365
rect 16416 -9205 16425 -8365
rect 16521 -9205 16530 -8365
rect 16530 -9205 16564 -8365
rect 16564 -9205 16573 -8365
rect 16669 -9205 16678 -8365
rect 16678 -9205 16712 -8365
rect 16712 -9205 16721 -8365
rect 16817 -9205 16826 -8365
rect 16826 -9205 16860 -8365
rect 16860 -9205 16869 -8365
rect 16965 -9205 16974 -8365
rect 16974 -9205 17008 -8365
rect 17008 -9205 17017 -8365
rect 17113 -9205 17122 -8365
rect 17122 -9205 17156 -8365
rect 17156 -9205 17165 -8365
rect 17261 -9205 17270 -8365
rect 17270 -9205 17304 -8365
rect 17304 -9205 17313 -8365
rect 17409 -9205 17418 -8365
rect 17418 -9205 17452 -8365
rect 17452 -9205 17461 -8365
rect 17557 -9205 17566 -8365
rect 17566 -9205 17600 -8365
rect 17600 -9205 17609 -8365
rect 17705 -9205 17714 -8365
rect 17714 -9205 17748 -8365
rect 17748 -9205 17757 -8365
rect 17853 -9205 17862 -8365
rect 17862 -9205 17896 -8365
rect 17896 -9205 17905 -8365
rect 18001 -9205 18010 -8365
rect 18010 -9205 18044 -8365
rect 18044 -9205 18053 -8365
rect 18149 -9205 18158 -8365
rect 18158 -9205 18192 -8365
rect 18192 -9205 18201 -8365
rect 18297 -9205 18306 -8365
rect 18306 -9205 18340 -8365
rect 18340 -9205 18349 -8365
rect 18445 -9205 18454 -8365
rect 18454 -9205 18488 -8365
rect 18488 -9205 18497 -8365
rect 18593 -9205 18602 -8365
rect 18602 -9205 18636 -8365
rect 18636 -9205 18645 -8365
rect 18741 -9205 18750 -8365
rect 18750 -9205 18784 -8365
rect 18784 -9205 18793 -8365
rect 18889 -9205 18898 -8365
rect 18898 -9205 18932 -8365
rect 18932 -9205 18941 -8365
rect 19037 -9205 19046 -8365
rect 19046 -9205 19080 -8365
rect 19080 -9205 19089 -8365
rect 19185 -9205 19194 -8365
rect 19194 -9205 19228 -8365
rect 19228 -9205 19237 -8365
rect 19333 -9205 19342 -8365
rect 19342 -9205 19376 -8365
rect 19376 -9205 19385 -8365
rect 19481 -9205 19490 -8365
rect 19490 -9205 19524 -8365
rect 19524 -9205 19533 -8365
rect 19629 -9205 19638 -8365
rect 19638 -9205 19672 -8365
rect 19672 -9205 19681 -8365
rect 19777 -9205 19786 -8365
rect 19786 -9205 19820 -8365
rect 19820 -9205 19829 -8365
rect 19925 -9205 19934 -8365
rect 19934 -9205 19968 -8365
rect 19968 -9205 19977 -8365
rect 20073 -9205 20082 -8365
rect 20082 -9205 20116 -8365
rect 20116 -9205 20125 -8365
rect 20221 -9205 20230 -8365
rect 20230 -9205 20264 -8365
rect 20264 -9205 20273 -8365
rect 20369 -9205 20378 -8365
rect 20378 -9205 20412 -8365
rect 20412 -9205 20421 -8365
rect 20517 -9205 20526 -8365
rect 20526 -9205 20560 -8365
rect 20560 -9205 20569 -8365
rect 20665 -9205 20674 -8365
rect 20674 -9205 20708 -8365
rect 20708 -9205 20717 -8365
rect 20813 -9205 20822 -8365
rect 20822 -9205 20856 -8365
rect 20856 -9205 20865 -8365
rect 20961 -9205 20970 -8365
rect 20970 -9205 21004 -8365
rect 21004 -9205 21013 -8365
rect 21109 -9205 21118 -8365
rect 21118 -9205 21152 -8365
rect 21152 -9205 21161 -8365
rect 21257 -9205 21266 -8365
rect 21266 -9205 21300 -8365
rect 21300 -9205 21309 -8365
rect 21405 -9205 21414 -8365
rect 21414 -9205 21448 -8365
rect 21448 -9205 21457 -8365
rect 21553 -9205 21562 -8365
rect 21562 -9205 21596 -8365
rect 21596 -9205 21605 -8365
rect 21701 -9205 21710 -8365
rect 21710 -9205 21744 -8365
rect 21744 -9205 21753 -8365
rect 21849 -9205 21858 -8365
rect 21858 -9205 21892 -8365
rect 21892 -9205 21901 -8365
rect 21997 -9205 22006 -8365
rect 22006 -9205 22040 -8365
rect 22040 -9205 22049 -8365
rect 22145 -9205 22154 -8365
rect 22154 -9205 22188 -8365
rect 22188 -9205 22197 -8365
rect 22293 -9205 22302 -8365
rect 22302 -9205 22336 -8365
rect 22336 -9205 22345 -8365
rect 22441 -9205 22450 -8365
rect 22450 -9205 22484 -8365
rect 22484 -9205 22493 -8365
rect 22589 -9205 22598 -8365
rect 22598 -9205 22632 -8365
rect 22632 -9205 22641 -8365
rect 22737 -9205 22746 -8365
rect 22746 -9205 22780 -8365
rect 22780 -9205 22789 -8365
rect 22885 -9205 22894 -8365
rect 22894 -9205 22928 -8365
rect 22928 -9205 22937 -8365
rect 23033 -9205 23042 -8365
rect 23042 -9205 23076 -8365
rect 23076 -9205 23085 -8365
rect 23181 -9205 23190 -8365
rect 23190 -9205 23224 -8365
rect 23224 -9205 23233 -8365
rect 23329 -9205 23338 -8365
rect 23338 -9205 23372 -8365
rect 23372 -9205 23381 -8365
rect 23477 -9205 23529 -8365
rect 23625 -9205 23677 -8365
rect 4055 -9735 4107 -9683
rect 4055 -9839 4107 -9787
rect 4055 -9943 4107 -9891
rect 4136 -9735 4188 -9683
rect 4136 -9839 4188 -9787
rect 4136 -9943 4188 -9891
rect 4217 -9735 4269 -9683
rect 4217 -9839 4269 -9787
rect 4217 -9943 4269 -9891
rect 4298 -9735 4350 -9683
rect 4379 -9735 4431 -9683
rect 4460 -9735 4512 -9683
rect 4541 -9735 4593 -9683
rect 4623 -9735 4675 -9683
rect 4704 -9735 4756 -9683
rect 4785 -9735 4837 -9683
rect 4298 -9839 4350 -9787
rect 4379 -9839 4431 -9787
rect 4460 -9839 4512 -9787
rect 4541 -9839 4593 -9787
rect 4623 -9839 4675 -9787
rect 4704 -9839 4756 -9787
rect 4785 -9839 4837 -9787
rect 4298 -9943 4350 -9891
rect 4379 -9943 4431 -9891
rect 4460 -9943 4512 -9891
rect 4541 -9943 4593 -9891
rect 4623 -9943 4675 -9891
rect 4704 -9943 4756 -9891
rect 4785 -9943 4837 -9891
rect 4866 -9735 4918 -9683
rect 4866 -9839 4918 -9787
rect 4866 -9943 4918 -9891
rect 4947 -9735 4999 -9683
rect 4947 -9839 4999 -9787
rect 4947 -9943 4999 -9891
rect 5028 -9735 5080 -9683
rect 5028 -9839 5080 -9787
rect 5028 -9943 5080 -9891
rect 5109 -9735 5161 -9683
rect 5191 -9735 5243 -9683
rect 5272 -9735 5324 -9683
rect 5353 -9735 5405 -9683
rect 5434 -9735 5486 -9683
rect 5515 -9735 5567 -9683
rect 5596 -9735 5648 -9683
rect 5677 -9735 5729 -9683
rect 5109 -9839 5161 -9787
rect 5191 -9839 5243 -9787
rect 5272 -9839 5324 -9787
rect 5353 -9839 5405 -9787
rect 5434 -9839 5486 -9787
rect 5515 -9839 5567 -9787
rect 5596 -9839 5648 -9787
rect 5677 -9839 5729 -9787
rect 5109 -9943 5161 -9891
rect 5191 -9943 5243 -9891
rect 5272 -9943 5324 -9891
rect 5353 -9943 5405 -9891
rect 5434 -9943 5486 -9891
rect 5515 -9943 5567 -9891
rect 5596 -9943 5648 -9891
rect 5677 -9943 5729 -9891
rect 5759 -9735 5811 -9683
rect 5759 -9839 5811 -9787
rect 5759 -9943 5811 -9891
rect 5840 -9735 5892 -9683
rect 5840 -9839 5892 -9787
rect 5840 -9943 5892 -9891
rect 5921 -9735 5973 -9683
rect 5921 -9839 5973 -9787
rect 5921 -9943 5973 -9891
rect 6002 -9735 6054 -9683
rect 6083 -9735 6135 -9683
rect 6164 -9735 6216 -9683
rect 6245 -9735 6297 -9683
rect 6327 -9735 6379 -9683
rect 6408 -9735 6460 -9683
rect 6489 -9735 6541 -9683
rect 6002 -9839 6054 -9787
rect 6083 -9839 6135 -9787
rect 6164 -9839 6216 -9787
rect 6245 -9839 6297 -9787
rect 6327 -9839 6379 -9787
rect 6408 -9839 6460 -9787
rect 6489 -9839 6541 -9787
rect 6002 -9943 6054 -9891
rect 6083 -9943 6135 -9891
rect 6164 -9943 6216 -9891
rect 6245 -9943 6297 -9891
rect 6327 -9943 6379 -9891
rect 6408 -9943 6460 -9891
rect 6489 -9943 6541 -9891
rect 6570 -9735 6622 -9683
rect 6570 -9839 6622 -9787
rect 6570 -9943 6622 -9891
rect 6651 -9735 6703 -9683
rect 6651 -9839 6703 -9787
rect 6651 -9943 6703 -9891
rect 6732 -9735 6784 -9683
rect 6732 -9839 6784 -9787
rect 6732 -9943 6784 -9891
rect 6813 -9735 6865 -9683
rect 6895 -9735 6947 -9683
rect 6976 -9735 7028 -9683
rect 7057 -9735 7109 -9683
rect 7138 -9735 7190 -9683
rect 7219 -9735 7271 -9683
rect 7300 -9735 7352 -9683
rect 7381 -9735 7433 -9683
rect 6813 -9839 6865 -9787
rect 6895 -9839 6947 -9787
rect 6976 -9839 7028 -9787
rect 7057 -9839 7109 -9787
rect 7138 -9839 7190 -9787
rect 7219 -9839 7271 -9787
rect 7300 -9839 7352 -9787
rect 7381 -9839 7433 -9787
rect 6813 -9943 6865 -9891
rect 6895 -9943 6947 -9891
rect 6976 -9943 7028 -9891
rect 7057 -9943 7109 -9891
rect 7138 -9943 7190 -9891
rect 7219 -9943 7271 -9891
rect 7300 -9943 7352 -9891
rect 7381 -9943 7433 -9891
rect 7463 -9735 7515 -9683
rect 7463 -9839 7515 -9787
rect 7463 -9943 7515 -9891
rect 7544 -9735 7596 -9683
rect 7544 -9839 7596 -9787
rect 7544 -9943 7596 -9891
rect 7625 -9735 7677 -9683
rect 7706 -9735 7758 -9683
rect 7787 -9735 7839 -9683
rect 7868 -9735 7920 -9683
rect 7949 -9735 8001 -9683
rect 8031 -9735 8083 -9683
rect 8112 -9735 8164 -9683
rect 8193 -9735 8245 -9683
rect 7625 -9839 7677 -9787
rect 7706 -9839 7758 -9787
rect 7787 -9839 7839 -9787
rect 7868 -9839 7920 -9787
rect 7949 -9839 8001 -9787
rect 8031 -9839 8083 -9787
rect 8112 -9839 8164 -9787
rect 8193 -9839 8245 -9787
rect 7625 -9943 7677 -9891
rect 7706 -9943 7758 -9891
rect 7787 -9943 7839 -9891
rect 7868 -9943 7920 -9891
rect 7949 -9943 8001 -9891
rect 8031 -9943 8083 -9891
rect 8112 -9943 8164 -9891
rect 8193 -9943 8245 -9891
rect 8274 -9735 8326 -9683
rect 8274 -9839 8326 -9787
rect 8274 -9943 8326 -9891
rect 8355 -9735 8407 -9683
rect 8355 -9839 8407 -9787
rect 8355 -9943 8407 -9891
rect 8436 -9735 8488 -9683
rect 8436 -9839 8488 -9787
rect 8436 -9943 8488 -9891
rect 8517 -9735 8569 -9683
rect 8599 -9735 8651 -9683
rect 8680 -9735 8732 -9683
rect 8761 -9735 8813 -9683
rect 8842 -9735 8894 -9683
rect 8923 -9735 8975 -9683
rect 9004 -9735 9056 -9683
rect 8517 -9839 8569 -9787
rect 8599 -9839 8651 -9787
rect 8680 -9839 8732 -9787
rect 8761 -9839 8813 -9787
rect 8842 -9839 8894 -9787
rect 8923 -9839 8975 -9787
rect 9004 -9839 9056 -9787
rect 8517 -9943 8569 -9891
rect 8599 -9943 8651 -9891
rect 8680 -9943 8732 -9891
rect 8761 -9943 8813 -9891
rect 8842 -9943 8894 -9891
rect 8923 -9943 8975 -9891
rect 9004 -9943 9056 -9891
rect 9085 -9735 9137 -9683
rect 9085 -9839 9137 -9787
rect 9085 -9943 9137 -9891
rect 9167 -9735 9219 -9683
rect 9167 -9839 9219 -9787
rect 9167 -9943 9219 -9891
rect 9248 -9735 9300 -9683
rect 9248 -9839 9300 -9787
rect 9248 -9943 9300 -9891
rect 9329 -9735 9381 -9683
rect 9410 -9735 9462 -9683
rect 9491 -9735 9543 -9683
rect 9572 -9735 9624 -9683
rect 9653 -9735 9705 -9683
rect 9735 -9735 9787 -9683
rect 9816 -9735 9868 -9683
rect 9897 -9735 9949 -9683
rect 9329 -9839 9381 -9787
rect 9410 -9839 9462 -9787
rect 9491 -9839 9543 -9787
rect 9572 -9839 9624 -9787
rect 9653 -9839 9705 -9787
rect 9735 -9839 9787 -9787
rect 9816 -9839 9868 -9787
rect 9897 -9839 9949 -9787
rect 9329 -9943 9381 -9891
rect 9410 -9943 9462 -9891
rect 9491 -9943 9543 -9891
rect 9572 -9943 9624 -9891
rect 9653 -9943 9705 -9891
rect 9735 -9943 9787 -9891
rect 9816 -9943 9868 -9891
rect 9897 -9943 9949 -9891
rect 9978 -9735 10030 -9683
rect 9978 -9839 10030 -9787
rect 9978 -9943 10030 -9891
rect 10059 -9735 10111 -9683
rect 10059 -9839 10111 -9787
rect 10059 -9943 10111 -9891
rect 10140 -9735 10192 -9683
rect 10221 -9735 10273 -9683
rect 10303 -9735 10355 -9683
rect 10384 -9735 10436 -9683
rect 10465 -9735 10517 -9683
rect 10546 -9735 10598 -9683
rect 10627 -9735 10679 -9683
rect 10708 -9735 10760 -9683
rect 10140 -9839 10192 -9787
rect 10221 -9839 10273 -9787
rect 10303 -9839 10355 -9787
rect 10384 -9839 10436 -9787
rect 10465 -9839 10517 -9787
rect 10546 -9839 10598 -9787
rect 10627 -9839 10679 -9787
rect 10708 -9839 10760 -9787
rect 10140 -9943 10192 -9891
rect 10221 -9943 10273 -9891
rect 10303 -9943 10355 -9891
rect 10384 -9943 10436 -9891
rect 10465 -9943 10517 -9891
rect 10546 -9943 10598 -9891
rect 10627 -9943 10679 -9891
rect 10708 -9943 10760 -9891
rect 10789 -9735 10841 -9683
rect 10789 -9839 10841 -9787
rect 10789 -9943 10841 -9891
rect 10871 -9735 10923 -9683
rect 10871 -9839 10923 -9787
rect 10871 -9943 10923 -9891
rect 10952 -9735 11004 -9683
rect 10952 -9839 11004 -9787
rect 10952 -9943 11004 -9891
rect 11033 -9735 11085 -9683
rect 11114 -9735 11166 -9683
rect 11195 -9735 11247 -9683
rect 11276 -9735 11328 -9683
rect 11357 -9735 11409 -9683
rect 11439 -9735 11491 -9683
rect 11520 -9735 11572 -9683
rect 11033 -9839 11085 -9787
rect 11114 -9839 11166 -9787
rect 11195 -9839 11247 -9787
rect 11276 -9839 11328 -9787
rect 11357 -9839 11409 -9787
rect 11439 -9839 11491 -9787
rect 11520 -9839 11572 -9787
rect 11033 -9943 11085 -9891
rect 11114 -9943 11166 -9891
rect 11195 -9943 11247 -9891
rect 11276 -9943 11328 -9891
rect 11357 -9943 11409 -9891
rect 11439 -9943 11491 -9891
rect 11520 -9943 11572 -9891
rect 11601 -9735 11653 -9683
rect 11601 -9839 11653 -9787
rect 11601 -9943 11653 -9891
rect 11682 -9735 11734 -9683
rect 11682 -9839 11734 -9787
rect 11682 -9943 11734 -9891
rect 11763 -9735 11815 -9683
rect 11763 -9839 11815 -9787
rect 11763 -9943 11815 -9891
rect 11844 -9735 11896 -9683
rect 11925 -9735 11977 -9683
rect 12007 -9735 12059 -9683
rect 12088 -9735 12140 -9683
rect 12169 -9735 12221 -9683
rect 12250 -9735 12302 -9683
rect 12331 -9735 12383 -9683
rect 12412 -9735 12464 -9683
rect 11844 -9839 11896 -9787
rect 11925 -9839 11977 -9787
rect 12007 -9839 12059 -9787
rect 12088 -9839 12140 -9787
rect 12169 -9839 12221 -9787
rect 12250 -9839 12302 -9787
rect 12331 -9839 12383 -9787
rect 12412 -9839 12464 -9787
rect 11844 -9943 11896 -9891
rect 11925 -9943 11977 -9891
rect 12007 -9943 12059 -9891
rect 12088 -9943 12140 -9891
rect 12169 -9943 12221 -9891
rect 12250 -9943 12302 -9891
rect 12331 -9943 12383 -9891
rect 12412 -9943 12464 -9891
rect 12493 -9735 12545 -9683
rect 12493 -9839 12545 -9787
rect 12493 -9943 12545 -9891
rect 12575 -9735 12627 -9683
rect 12575 -9839 12627 -9787
rect 12575 -9943 12627 -9891
rect 12656 -9735 12708 -9683
rect 12737 -9735 12789 -9683
rect 12818 -9735 12870 -9683
rect 12899 -9735 12951 -9683
rect 12980 -9735 13032 -9683
rect 13061 -9735 13113 -9683
rect 13143 -9735 13195 -9683
rect 13224 -9735 13276 -9683
rect 12656 -9839 12708 -9787
rect 12737 -9839 12789 -9787
rect 12818 -9839 12870 -9787
rect 12899 -9839 12951 -9787
rect 12980 -9839 13032 -9787
rect 13061 -9839 13113 -9787
rect 13143 -9839 13195 -9787
rect 13224 -9839 13276 -9787
rect 12656 -9943 12708 -9891
rect 12737 -9943 12789 -9891
rect 12818 -9943 12870 -9891
rect 12899 -9943 12951 -9891
rect 12980 -9943 13032 -9891
rect 13061 -9943 13113 -9891
rect 13143 -9943 13195 -9891
rect 13224 -9943 13276 -9891
rect 13305 -9735 13357 -9683
rect 13305 -9839 13357 -9787
rect 13305 -9943 13357 -9891
rect 13386 -9735 13438 -9683
rect 13386 -9839 13438 -9787
rect 13386 -9943 13438 -9891
rect 13467 -9735 13519 -9683
rect 13467 -9839 13519 -9787
rect 13467 -9943 13519 -9891
rect 13548 -9735 13600 -9683
rect 13629 -9735 13681 -9683
rect 13711 -9735 13763 -9683
rect 13792 -9735 13844 -9683
rect 13873 -9735 13925 -9683
rect 13954 -9735 14006 -9683
rect 14035 -9735 14087 -9683
rect 13548 -9839 13600 -9787
rect 13629 -9839 13681 -9787
rect 13711 -9839 13763 -9787
rect 13792 -9839 13844 -9787
rect 13873 -9839 13925 -9787
rect 13954 -9839 14006 -9787
rect 14035 -9839 14087 -9787
rect 13548 -9943 13600 -9891
rect 13629 -9943 13681 -9891
rect 13711 -9943 13763 -9891
rect 13792 -9943 13844 -9891
rect 13873 -9943 13925 -9891
rect 13954 -9943 14006 -9891
rect 14035 -9943 14087 -9891
rect 14116 -9735 14168 -9683
rect 14116 -9839 14168 -9787
rect 14116 -9943 14168 -9891
rect 14197 -9735 14249 -9683
rect 14197 -9839 14249 -9787
rect 14197 -9943 14249 -9891
rect 14279 -9735 14331 -9683
rect 14279 -9839 14331 -9787
rect 14279 -9943 14331 -9891
rect 14360 -9735 14412 -9683
rect 14441 -9735 14493 -9683
rect 14522 -9735 14574 -9683
rect 14603 -9735 14655 -9683
rect 14684 -9735 14736 -9683
rect 14765 -9735 14817 -9683
rect 14847 -9735 14899 -9683
rect 14928 -9735 14980 -9683
rect 14360 -9839 14412 -9787
rect 14441 -9839 14493 -9787
rect 14522 -9839 14574 -9787
rect 14603 -9839 14655 -9787
rect 14684 -9839 14736 -9787
rect 14765 -9839 14817 -9787
rect 14847 -9839 14899 -9787
rect 14928 -9839 14980 -9787
rect 14360 -9943 14412 -9891
rect 14441 -9943 14493 -9891
rect 14522 -9943 14574 -9891
rect 14603 -9943 14655 -9891
rect 14684 -9943 14736 -9891
rect 14765 -9943 14817 -9891
rect 14847 -9943 14899 -9891
rect 14928 -9943 14980 -9891
rect 15009 -9735 15061 -9683
rect 15009 -9839 15061 -9787
rect 15009 -9943 15061 -9891
rect 15090 -9735 15142 -9683
rect 15090 -9839 15142 -9787
rect 15090 -9943 15142 -9891
rect 15171 -9735 15223 -9683
rect 15171 -9839 15223 -9787
rect 15171 -9943 15223 -9891
rect 15252 -9735 15304 -9683
rect 15333 -9735 15385 -9683
rect 15415 -9735 15467 -9683
rect 15496 -9735 15548 -9683
rect 15577 -9735 15629 -9683
rect 15658 -9735 15710 -9683
rect 15739 -9735 15791 -9683
rect 15252 -9839 15304 -9787
rect 15333 -9839 15385 -9787
rect 15415 -9839 15467 -9787
rect 15496 -9839 15548 -9787
rect 15577 -9839 15629 -9787
rect 15658 -9839 15710 -9787
rect 15739 -9839 15791 -9787
rect 15252 -9943 15304 -9891
rect 15333 -9943 15385 -9891
rect 15415 -9943 15467 -9891
rect 15496 -9943 15548 -9891
rect 15577 -9943 15629 -9891
rect 15658 -9943 15710 -9891
rect 15739 -9943 15791 -9891
rect 15820 -9735 15872 -9683
rect 15820 -9839 15872 -9787
rect 15820 -9943 15872 -9891
rect 15901 -9735 15953 -9683
rect 15901 -9839 15953 -9787
rect 15901 -9943 15953 -9891
rect 15983 -9735 16035 -9683
rect 15983 -9839 16035 -9787
rect 15983 -9943 16035 -9891
rect 16064 -9735 16116 -9683
rect 16145 -9735 16197 -9683
rect 16226 -9735 16278 -9683
rect 16307 -9735 16359 -9683
rect 16388 -9735 16440 -9683
rect 16469 -9735 16521 -9683
rect 16551 -9735 16603 -9683
rect 16064 -9839 16116 -9787
rect 16145 -9839 16197 -9787
rect 16226 -9839 16278 -9787
rect 16307 -9839 16359 -9787
rect 16388 -9839 16440 -9787
rect 16469 -9839 16521 -9787
rect 16551 -9839 16603 -9787
rect 16064 -9943 16116 -9891
rect 16145 -9943 16197 -9891
rect 16226 -9943 16278 -9891
rect 16307 -9943 16359 -9891
rect 16388 -9943 16440 -9891
rect 16469 -9943 16521 -9891
rect 16551 -9943 16603 -9891
rect 16632 -9735 16684 -9683
rect 16632 -9839 16684 -9787
rect 16632 -9943 16684 -9891
rect 16713 -9735 16765 -9683
rect 16713 -9839 16765 -9787
rect 16713 -9943 16765 -9891
rect 16794 -9735 16846 -9683
rect 16794 -9839 16846 -9787
rect 16794 -9943 16846 -9891
rect 16875 -9735 16927 -9683
rect 16956 -9735 17008 -9683
rect 17037 -9735 17089 -9683
rect 17119 -9735 17171 -9683
rect 17200 -9735 17252 -9683
rect 17281 -9735 17333 -9683
rect 17362 -9735 17414 -9683
rect 17443 -9735 17495 -9683
rect 16875 -9839 16927 -9787
rect 16956 -9839 17008 -9787
rect 17037 -9839 17089 -9787
rect 17119 -9839 17171 -9787
rect 17200 -9839 17252 -9787
rect 17281 -9839 17333 -9787
rect 17362 -9839 17414 -9787
rect 17443 -9839 17495 -9787
rect 16875 -9943 16927 -9891
rect 16956 -9943 17008 -9891
rect 17037 -9943 17089 -9891
rect 17119 -9943 17171 -9891
rect 17200 -9943 17252 -9891
rect 17281 -9943 17333 -9891
rect 17362 -9943 17414 -9891
rect 17443 -9943 17495 -9891
rect 17524 -9735 17576 -9683
rect 17524 -9839 17576 -9787
rect 17524 -9943 17576 -9891
rect 17605 -9735 17657 -9683
rect 17605 -9839 17657 -9787
rect 17605 -9943 17657 -9891
rect 17686 -9735 17738 -9683
rect 17686 -9839 17738 -9787
rect 17686 -9943 17738 -9891
rect 17767 -9735 17819 -9683
rect 17848 -9735 17900 -9683
rect 17929 -9735 17981 -9683
rect 18010 -9735 18062 -9683
rect 18091 -9735 18143 -9683
rect 18173 -9735 18225 -9683
rect 18254 -9735 18306 -9683
rect 17767 -9839 17819 -9787
rect 17848 -9839 17900 -9787
rect 17929 -9839 17981 -9787
rect 18010 -9839 18062 -9787
rect 18091 -9839 18143 -9787
rect 18173 -9839 18225 -9787
rect 18254 -9839 18306 -9787
rect 17767 -9943 17819 -9891
rect 17848 -9943 17900 -9891
rect 17929 -9943 17981 -9891
rect 18010 -9943 18062 -9891
rect 18091 -9943 18143 -9891
rect 18173 -9943 18225 -9891
rect 18254 -9943 18306 -9891
rect 18335 -9735 18387 -9683
rect 18335 -9839 18387 -9787
rect 18335 -9943 18387 -9891
rect 18416 -9735 18468 -9683
rect 18416 -9839 18468 -9787
rect 18416 -9943 18468 -9891
rect 18497 -9735 18549 -9683
rect 18497 -9839 18549 -9787
rect 18497 -9943 18549 -9891
rect 18578 -9735 18630 -9683
rect 18659 -9735 18711 -9683
rect 18741 -9735 18793 -9683
rect 18822 -9735 18874 -9683
rect 18903 -9735 18955 -9683
rect 18984 -9735 19036 -9683
rect 19065 -9735 19117 -9683
rect 19146 -9735 19198 -9683
rect 18578 -9839 18630 -9787
rect 18659 -9839 18711 -9787
rect 18741 -9839 18793 -9787
rect 18822 -9839 18874 -9787
rect 18903 -9839 18955 -9787
rect 18984 -9839 19036 -9787
rect 19065 -9839 19117 -9787
rect 19146 -9839 19198 -9787
rect 18578 -9943 18630 -9891
rect 18659 -9943 18711 -9891
rect 18741 -9943 18793 -9891
rect 18822 -9943 18874 -9891
rect 18903 -9943 18955 -9891
rect 18984 -9943 19036 -9891
rect 19065 -9943 19117 -9891
rect 19146 -9943 19198 -9891
rect 19227 -9735 19279 -9683
rect 19227 -9839 19279 -9787
rect 19227 -9943 19279 -9891
rect 19309 -9735 19361 -9683
rect 19309 -9839 19361 -9787
rect 19309 -9943 19361 -9891
rect 19390 -9735 19442 -9683
rect 19471 -9735 19523 -9683
rect 19552 -9735 19604 -9683
rect 19633 -9735 19685 -9683
rect 19714 -9735 19766 -9683
rect 19795 -9735 19847 -9683
rect 19877 -9735 19929 -9683
rect 19958 -9735 20010 -9683
rect 19390 -9839 19442 -9787
rect 19471 -9839 19523 -9787
rect 19552 -9839 19604 -9787
rect 19633 -9839 19685 -9787
rect 19714 -9839 19766 -9787
rect 19795 -9839 19847 -9787
rect 19877 -9839 19929 -9787
rect 19958 -9839 20010 -9787
rect 19390 -9943 19442 -9891
rect 19471 -9943 19523 -9891
rect 19552 -9943 19604 -9891
rect 19633 -9943 19685 -9891
rect 19714 -9943 19766 -9891
rect 19795 -9943 19847 -9891
rect 19877 -9943 19929 -9891
rect 19958 -9943 20010 -9891
rect 20039 -9735 20091 -9683
rect 20039 -9839 20091 -9787
rect 20039 -9943 20091 -9891
rect 20120 -9735 20172 -9683
rect 20120 -9839 20172 -9787
rect 20120 -9943 20172 -9891
rect 20201 -9735 20253 -9683
rect 20201 -9839 20253 -9787
rect 20201 -9943 20253 -9891
rect 20282 -9735 20334 -9683
rect 20363 -9735 20415 -9683
rect 20445 -9735 20497 -9683
rect 20526 -9735 20578 -9683
rect 20607 -9735 20659 -9683
rect 20688 -9735 20740 -9683
rect 20769 -9735 20821 -9683
rect 20282 -9839 20334 -9787
rect 20363 -9839 20415 -9787
rect 20445 -9839 20497 -9787
rect 20526 -9839 20578 -9787
rect 20607 -9839 20659 -9787
rect 20688 -9839 20740 -9787
rect 20769 -9839 20821 -9787
rect 20282 -9943 20334 -9891
rect 20363 -9943 20415 -9891
rect 20445 -9943 20497 -9891
rect 20526 -9943 20578 -9891
rect 20607 -9943 20659 -9891
rect 20688 -9943 20740 -9891
rect 20769 -9943 20821 -9891
rect 20850 -9735 20902 -9683
rect 20850 -9839 20902 -9787
rect 20850 -9943 20902 -9891
rect 20931 -9735 20983 -9683
rect 20931 -9839 20983 -9787
rect 20931 -9943 20983 -9891
rect 21013 -9735 21065 -9683
rect 21013 -9839 21065 -9787
rect 21013 -9943 21065 -9891
rect 21094 -9735 21146 -9683
rect 21175 -9735 21227 -9683
rect 21256 -9735 21308 -9683
rect 21337 -9735 21389 -9683
rect 21418 -9735 21470 -9683
rect 21499 -9735 21551 -9683
rect 21581 -9735 21633 -9683
rect 21662 -9735 21714 -9683
rect 21094 -9839 21146 -9787
rect 21175 -9839 21227 -9787
rect 21256 -9839 21308 -9787
rect 21337 -9839 21389 -9787
rect 21418 -9839 21470 -9787
rect 21499 -9839 21551 -9787
rect 21581 -9839 21633 -9787
rect 21662 -9839 21714 -9787
rect 21094 -9943 21146 -9891
rect 21175 -9943 21227 -9891
rect 21256 -9943 21308 -9891
rect 21337 -9943 21389 -9891
rect 21418 -9943 21470 -9891
rect 21499 -9943 21551 -9891
rect 21581 -9943 21633 -9891
rect 21662 -9943 21714 -9891
rect 21743 -9735 21795 -9683
rect 21743 -9839 21795 -9787
rect 21743 -9943 21795 -9891
rect 21824 -9735 21876 -9683
rect 21824 -9839 21876 -9787
rect 21824 -9943 21876 -9891
rect 21905 -9735 21957 -9683
rect 21905 -9839 21957 -9787
rect 21905 -9943 21957 -9891
rect 21986 -9735 22038 -9683
rect 22067 -9735 22119 -9683
rect 22149 -9735 22201 -9683
rect 22230 -9735 22282 -9683
rect 22311 -9735 22363 -9683
rect 22392 -9735 22444 -9683
rect 22473 -9735 22525 -9683
rect 21986 -9839 22038 -9787
rect 22067 -9839 22119 -9787
rect 22149 -9839 22201 -9787
rect 22230 -9839 22282 -9787
rect 22311 -9839 22363 -9787
rect 22392 -9839 22444 -9787
rect 22473 -9839 22525 -9787
rect 21986 -9943 22038 -9891
rect 22067 -9943 22119 -9891
rect 22149 -9943 22201 -9891
rect 22230 -9943 22282 -9891
rect 22311 -9943 22363 -9891
rect 22392 -9943 22444 -9891
rect 22473 -9943 22525 -9891
rect 22554 -9735 22606 -9683
rect 22554 -9839 22606 -9787
rect 22554 -9943 22606 -9891
rect 22635 -9735 22687 -9683
rect 22635 -9839 22687 -9787
rect 22635 -9943 22687 -9891
rect 22717 -9735 22769 -9683
rect 22717 -9839 22769 -9787
rect 22717 -9943 22769 -9891
rect 22798 -9735 22850 -9683
rect 22879 -9735 22931 -9683
rect 22960 -9735 23012 -9683
rect 23041 -9735 23093 -9683
rect 23122 -9735 23174 -9683
rect 23203 -9735 23255 -9683
rect 23285 -9735 23337 -9683
rect 22798 -9839 22850 -9787
rect 22879 -9839 22931 -9787
rect 22960 -9839 23012 -9787
rect 23041 -9839 23093 -9787
rect 23122 -9839 23174 -9787
rect 23203 -9839 23255 -9787
rect 23285 -9839 23337 -9787
rect 22798 -9943 22850 -9891
rect 22879 -9943 22931 -9891
rect 22960 -9943 23012 -9891
rect 23041 -9943 23093 -9891
rect 23122 -9943 23174 -9891
rect 23203 -9943 23255 -9891
rect 23285 -9943 23337 -9891
rect 23366 -9735 23418 -9683
rect 23366 -9839 23418 -9787
rect 23366 -9943 23418 -9891
rect 23447 -9735 23499 -9683
rect 23447 -9839 23499 -9787
rect 23447 -9943 23499 -9891
rect 23528 -9735 23580 -9683
rect 23528 -9839 23580 -9787
rect 23528 -9943 23580 -9891
rect 23609 -9735 23661 -9683
rect 23690 -9735 23742 -9683
rect 23771 -9735 23823 -9683
rect 23853 -9735 23905 -9683
rect 23934 -9735 23986 -9683
rect 24015 -9735 24067 -9683
rect 24096 -9735 24148 -9683
rect 24177 -9735 24229 -9683
rect 23609 -9839 23661 -9787
rect 23690 -9839 23742 -9787
rect 23771 -9839 23823 -9787
rect 23853 -9839 23905 -9787
rect 23934 -9839 23986 -9787
rect 24015 -9839 24067 -9787
rect 24096 -9839 24148 -9787
rect 24177 -9839 24229 -9787
rect 23609 -9943 23661 -9891
rect 23690 -9943 23742 -9891
rect 23771 -9943 23823 -9891
rect 23853 -9943 23905 -9891
rect 23934 -9943 23986 -9891
rect 24015 -9943 24067 -9891
rect 24096 -9943 24148 -9891
rect 24177 -9943 24229 -9891
rect 24258 -9735 24310 -9683
rect 24258 -9839 24310 -9787
rect 24258 -9943 24310 -9891
rect 24339 -9735 24391 -9683
rect 24339 -9839 24391 -9787
rect 24339 -9943 24391 -9891
rect 24421 -9735 24473 -9683
rect 24421 -9839 24473 -9787
rect 24421 -9943 24473 -9891
rect 24502 -9735 24554 -9683
rect 24583 -9735 24635 -9683
rect 24664 -9735 24716 -9683
rect 24745 -9735 24797 -9683
rect 24826 -9735 24878 -9683
rect 24907 -9735 24959 -9683
rect 24989 -9735 25041 -9683
rect 24502 -9839 24554 -9787
rect 24583 -9839 24635 -9787
rect 24664 -9839 24716 -9787
rect 24745 -9839 24797 -9787
rect 24826 -9839 24878 -9787
rect 24907 -9839 24959 -9787
rect 24989 -9839 25041 -9787
rect 24502 -9943 24554 -9891
rect 24583 -9943 24635 -9891
rect 24664 -9943 24716 -9891
rect 24745 -9943 24797 -9891
rect 24826 -9943 24878 -9891
rect 24907 -9943 24959 -9891
rect 24989 -9943 25041 -9891
rect 25070 -9735 25122 -9683
rect 25070 -9839 25122 -9787
rect 25070 -9943 25122 -9891
rect 25151 -9735 25203 -9683
rect 25151 -9839 25203 -9787
rect 25151 -9943 25203 -9891
rect 25232 -9735 25284 -9683
rect 25232 -9839 25284 -9787
rect 25232 -9943 25284 -9891
rect 25313 -9735 25365 -9683
rect 25394 -9735 25446 -9683
rect 25475 -9735 25527 -9683
rect 25557 -9735 25609 -9683
rect 25638 -9735 25690 -9683
rect 25719 -9735 25771 -9683
rect 25800 -9735 25852 -9683
rect 25881 -9735 25933 -9683
rect 25313 -9839 25365 -9787
rect 25394 -9839 25446 -9787
rect 25475 -9839 25527 -9787
rect 25557 -9839 25609 -9787
rect 25638 -9839 25690 -9787
rect 25719 -9839 25771 -9787
rect 25800 -9839 25852 -9787
rect 25881 -9839 25933 -9787
rect 25313 -9943 25365 -9891
rect 25394 -9943 25446 -9891
rect 25475 -9943 25527 -9891
rect 25557 -9943 25609 -9891
rect 25638 -9943 25690 -9891
rect 25719 -9943 25771 -9891
rect 25800 -9943 25852 -9891
rect 25881 -9943 25933 -9891
rect 25962 -9735 26014 -9683
rect 25962 -9839 26014 -9787
rect 25962 -9943 26014 -9891
rect 26043 -9735 26095 -9683
rect 26043 -9839 26095 -9787
rect 26043 -9943 26095 -9891
rect 26125 -9735 26177 -9683
rect 26206 -9735 26258 -9683
rect 26125 -9839 26177 -9787
rect 26206 -9839 26258 -9787
rect 26125 -9943 26177 -9891
rect 26206 -9943 26258 -9891
<< metal2 >>
rect 23903 3182 25067 3183
rect 3012 3174 25067 3182
rect 3012 3118 3036 3174
rect 3092 3118 3118 3174
rect 3174 3118 3199 3174
rect 3255 3118 3280 3174
rect 3336 3118 3361 3174
rect 3417 3118 3442 3174
rect 3498 3118 3523 3174
rect 3579 3118 3604 3174
rect 3660 3118 3686 3174
rect 3742 3118 3767 3174
rect 3823 3118 3848 3174
rect 3904 3118 3929 3174
rect 3985 3118 4010 3174
rect 4066 3118 4091 3174
rect 4147 3118 4172 3174
rect 4228 3118 4254 3174
rect 4310 3118 4335 3174
rect 4391 3118 4416 3174
rect 4472 3118 4497 3174
rect 4553 3118 4578 3174
rect 4634 3118 4659 3174
rect 4715 3118 4740 3174
rect 4796 3118 4822 3174
rect 4878 3118 4903 3174
rect 4959 3118 4984 3174
rect 5040 3118 5065 3174
rect 5121 3118 5146 3174
rect 5202 3118 5227 3174
rect 5283 3118 5308 3174
rect 5364 3118 5390 3174
rect 5446 3118 5471 3174
rect 5527 3118 5552 3174
rect 5608 3118 5633 3174
rect 5689 3118 5714 3174
rect 5770 3118 5795 3174
rect 5851 3118 5876 3174
rect 5932 3118 5958 3174
rect 6014 3118 6039 3174
rect 6095 3118 6120 3174
rect 6176 3118 6201 3174
rect 6257 3118 6282 3174
rect 6338 3118 6363 3174
rect 6419 3118 6444 3174
rect 6500 3118 6526 3174
rect 6582 3118 6607 3174
rect 6663 3118 6688 3174
rect 6744 3118 6769 3174
rect 6825 3118 6850 3174
rect 6906 3118 6931 3174
rect 6987 3118 7012 3174
rect 7068 3118 7094 3174
rect 7150 3118 7175 3174
rect 7231 3118 7256 3174
rect 7312 3118 7337 3174
rect 7393 3118 7418 3174
rect 7474 3118 7499 3174
rect 7555 3118 7580 3174
rect 7636 3118 7662 3174
rect 7718 3118 7743 3174
rect 7799 3118 7824 3174
rect 7880 3118 7905 3174
rect 7961 3118 7986 3174
rect 8042 3118 8067 3174
rect 8123 3118 8148 3174
rect 8204 3118 8230 3174
rect 8286 3118 8311 3174
rect 8367 3118 8392 3174
rect 8448 3118 8473 3174
rect 8529 3118 8554 3174
rect 8610 3118 8635 3174
rect 8691 3118 8716 3174
rect 8772 3118 8798 3174
rect 8854 3118 8879 3174
rect 8935 3118 8960 3174
rect 9016 3118 9041 3174
rect 9097 3118 9122 3174
rect 9178 3118 9203 3174
rect 9259 3118 9284 3174
rect 9340 3118 9366 3174
rect 9422 3118 9447 3174
rect 9503 3118 9528 3174
rect 9584 3118 9609 3174
rect 9665 3118 9690 3174
rect 9746 3118 9771 3174
rect 9827 3118 9852 3174
rect 9908 3118 9934 3174
rect 9990 3118 10015 3174
rect 10071 3118 10096 3174
rect 10152 3118 10177 3174
rect 10233 3118 10258 3174
rect 10314 3118 10339 3174
rect 10395 3118 10420 3174
rect 10476 3118 10502 3174
rect 10558 3118 10583 3174
rect 10639 3118 10664 3174
rect 10720 3118 10745 3174
rect 10801 3118 10826 3174
rect 10882 3118 10907 3174
rect 10963 3118 10988 3174
rect 11044 3118 11116 3174
rect 11172 3118 11197 3174
rect 11253 3118 11278 3174
rect 11334 3118 11359 3174
rect 11415 3118 11440 3174
rect 11496 3118 11521 3174
rect 11577 3118 11602 3174
rect 11658 3118 11684 3174
rect 11740 3118 11765 3174
rect 11821 3118 11846 3174
rect 11902 3118 11927 3174
rect 11983 3118 12008 3174
rect 12064 3118 12089 3174
rect 12145 3118 12170 3174
rect 12226 3118 12252 3174
rect 12308 3118 12333 3174
rect 12389 3118 12414 3174
rect 12470 3118 12495 3174
rect 12551 3118 12576 3174
rect 12632 3118 12657 3174
rect 12713 3118 12738 3174
rect 12794 3118 12820 3174
rect 12876 3118 12901 3174
rect 12957 3118 12982 3174
rect 13038 3118 13063 3174
rect 13119 3118 13144 3174
rect 13200 3118 13225 3174
rect 13281 3118 13306 3174
rect 13362 3118 13388 3174
rect 13444 3118 13469 3174
rect 13525 3118 13550 3174
rect 13606 3118 13631 3174
rect 13687 3118 13712 3174
rect 13768 3118 13793 3174
rect 13849 3118 13874 3174
rect 13930 3118 13956 3174
rect 14012 3118 14037 3174
rect 14093 3118 14118 3174
rect 14174 3118 14199 3174
rect 14255 3118 14280 3174
rect 14336 3118 14361 3174
rect 14417 3118 14442 3174
rect 14498 3118 14524 3174
rect 14580 3118 14605 3174
rect 14661 3118 14686 3174
rect 14742 3118 14767 3174
rect 14823 3118 14848 3174
rect 14904 3118 14929 3174
rect 14985 3118 15010 3174
rect 15066 3118 15092 3174
rect 15148 3118 15173 3174
rect 15229 3118 15254 3174
rect 15310 3118 15335 3174
rect 15391 3118 15416 3174
rect 15472 3118 15497 3174
rect 15553 3118 15578 3174
rect 15634 3118 15660 3174
rect 15716 3118 15741 3174
rect 15797 3118 15822 3174
rect 15878 3118 15903 3174
rect 15959 3118 15984 3174
rect 16040 3118 16065 3174
rect 16121 3118 16146 3174
rect 16202 3118 16228 3174
rect 16284 3118 16309 3174
rect 16365 3118 16390 3174
rect 16446 3118 16471 3174
rect 16527 3118 16552 3174
rect 16608 3118 16633 3174
rect 16689 3118 16714 3174
rect 16770 3118 16796 3174
rect 16852 3118 16877 3174
rect 16933 3118 16958 3174
rect 17014 3118 17039 3174
rect 17095 3118 17120 3174
rect 17176 3118 17201 3174
rect 17257 3118 17282 3174
rect 17338 3118 17364 3174
rect 17420 3118 17445 3174
rect 17501 3118 17526 3174
rect 17582 3118 17607 3174
rect 17663 3118 17688 3174
rect 17744 3118 17769 3174
rect 17825 3118 17850 3174
rect 17906 3118 17932 3174
rect 17988 3118 18013 3174
rect 18069 3118 18094 3174
rect 18150 3118 18175 3174
rect 18231 3118 18256 3174
rect 18312 3118 18337 3174
rect 18393 3118 18418 3174
rect 18474 3118 18500 3174
rect 18556 3118 18581 3174
rect 18637 3118 18662 3174
rect 18718 3118 18743 3174
rect 18799 3118 18824 3174
rect 18880 3118 18905 3174
rect 18961 3118 18986 3174
rect 19042 3118 19068 3174
rect 19124 3118 19149 3174
rect 19205 3118 19230 3174
rect 19286 3118 19311 3174
rect 19367 3118 19392 3174
rect 19448 3118 19473 3174
rect 19529 3118 19554 3174
rect 19610 3118 19636 3174
rect 19692 3118 19717 3174
rect 19773 3118 19798 3174
rect 19854 3118 19879 3174
rect 19935 3118 19960 3174
rect 20016 3118 20041 3174
rect 20097 3118 20122 3174
rect 20178 3118 20204 3174
rect 20260 3118 20285 3174
rect 20341 3118 20366 3174
rect 20422 3118 20447 3174
rect 20503 3118 20528 3174
rect 20584 3118 20609 3174
rect 20665 3118 20690 3174
rect 20746 3118 20772 3174
rect 20828 3118 20853 3174
rect 20909 3118 20934 3174
rect 20990 3118 21015 3174
rect 21071 3118 21096 3174
rect 21152 3118 21177 3174
rect 21233 3118 21258 3174
rect 21314 3118 21340 3174
rect 21396 3118 21421 3174
rect 21477 3118 21502 3174
rect 21558 3118 21583 3174
rect 21639 3118 21664 3174
rect 21720 3118 21745 3174
rect 21801 3118 21826 3174
rect 21882 3118 21908 3174
rect 21964 3118 21989 3174
rect 22045 3118 22070 3174
rect 22126 3118 22151 3174
rect 22207 3118 22232 3174
rect 22288 3118 22313 3174
rect 22369 3118 22394 3174
rect 22450 3118 22476 3174
rect 22532 3118 22557 3174
rect 22613 3118 22638 3174
rect 22694 3118 22719 3174
rect 22775 3118 22800 3174
rect 22856 3118 22881 3174
rect 22937 3118 22962 3174
rect 23018 3118 23044 3174
rect 23100 3118 23125 3174
rect 23181 3118 23206 3174
rect 23262 3118 23287 3174
rect 23343 3118 23368 3174
rect 23424 3118 23449 3174
rect 23505 3118 23530 3174
rect 23586 3118 23612 3174
rect 23668 3118 23693 3174
rect 23749 3118 23774 3174
rect 23830 3118 23855 3174
rect 23911 3118 23936 3174
rect 23992 3118 24017 3174
rect 24073 3118 24098 3174
rect 24154 3118 24180 3174
rect 24236 3118 24261 3174
rect 24317 3118 24342 3174
rect 24398 3118 24423 3174
rect 24479 3118 24504 3174
rect 24560 3118 24585 3174
rect 24641 3118 24666 3174
rect 24722 3118 25067 3174
rect 3012 3070 25067 3118
rect 3012 3014 3036 3070
rect 3092 3014 3118 3070
rect 3174 3014 3199 3070
rect 3255 3014 3280 3070
rect 3336 3014 3361 3070
rect 3417 3014 3442 3070
rect 3498 3014 3523 3070
rect 3579 3014 3604 3070
rect 3660 3014 3686 3070
rect 3742 3014 3767 3070
rect 3823 3014 3848 3070
rect 3904 3014 3929 3070
rect 3985 3014 4010 3070
rect 4066 3014 4091 3070
rect 4147 3014 4172 3070
rect 4228 3014 4254 3070
rect 4310 3014 4335 3070
rect 4391 3014 4416 3070
rect 4472 3014 4497 3070
rect 4553 3014 4578 3070
rect 4634 3014 4659 3070
rect 4715 3014 4740 3070
rect 4796 3014 4822 3070
rect 4878 3014 4903 3070
rect 4959 3014 4984 3070
rect 5040 3014 5065 3070
rect 5121 3014 5146 3070
rect 5202 3014 5227 3070
rect 5283 3014 5308 3070
rect 5364 3014 5390 3070
rect 5446 3014 5471 3070
rect 5527 3014 5552 3070
rect 5608 3014 5633 3070
rect 5689 3014 5714 3070
rect 5770 3014 5795 3070
rect 5851 3014 5876 3070
rect 5932 3014 5958 3070
rect 6014 3014 6039 3070
rect 6095 3014 6120 3070
rect 6176 3014 6201 3070
rect 6257 3014 6282 3070
rect 6338 3014 6363 3070
rect 6419 3014 6444 3070
rect 6500 3014 6526 3070
rect 6582 3014 6607 3070
rect 6663 3014 6688 3070
rect 6744 3014 6769 3070
rect 6825 3014 6850 3070
rect 6906 3014 6931 3070
rect 6987 3014 7012 3070
rect 7068 3014 7094 3070
rect 7150 3014 7175 3070
rect 7231 3014 7256 3070
rect 7312 3014 7337 3070
rect 7393 3014 7418 3070
rect 7474 3014 7499 3070
rect 7555 3014 7580 3070
rect 7636 3014 7662 3070
rect 7718 3014 7743 3070
rect 7799 3014 7824 3070
rect 7880 3014 7905 3070
rect 7961 3014 7986 3070
rect 8042 3014 8067 3070
rect 8123 3014 8148 3070
rect 8204 3014 8230 3070
rect 8286 3014 8311 3070
rect 8367 3014 8392 3070
rect 8448 3014 8473 3070
rect 8529 3014 8554 3070
rect 8610 3014 8635 3070
rect 8691 3014 8716 3070
rect 8772 3014 8798 3070
rect 8854 3014 8879 3070
rect 8935 3014 8960 3070
rect 9016 3014 9041 3070
rect 9097 3014 9122 3070
rect 9178 3014 9203 3070
rect 9259 3014 9284 3070
rect 9340 3014 9366 3070
rect 9422 3014 9447 3070
rect 9503 3014 9528 3070
rect 9584 3014 9609 3070
rect 9665 3014 9690 3070
rect 9746 3014 9771 3070
rect 9827 3014 9852 3070
rect 9908 3014 9934 3070
rect 9990 3014 10015 3070
rect 10071 3014 10096 3070
rect 10152 3014 10177 3070
rect 10233 3014 10258 3070
rect 10314 3014 10339 3070
rect 10395 3014 10420 3070
rect 10476 3014 10502 3070
rect 10558 3014 10583 3070
rect 10639 3014 10664 3070
rect 10720 3014 10745 3070
rect 10801 3014 10826 3070
rect 10882 3014 10907 3070
rect 10963 3014 10988 3070
rect 11044 3014 11116 3070
rect 11172 3014 11197 3070
rect 11253 3014 11278 3070
rect 11334 3014 11359 3070
rect 11415 3014 11440 3070
rect 11496 3014 11521 3070
rect 11577 3014 11602 3070
rect 11658 3014 11684 3070
rect 11740 3014 11765 3070
rect 11821 3014 11846 3070
rect 11902 3014 11927 3070
rect 11983 3014 12008 3070
rect 12064 3014 12089 3070
rect 12145 3014 12170 3070
rect 12226 3014 12252 3070
rect 12308 3014 12333 3070
rect 12389 3014 12414 3070
rect 12470 3014 12495 3070
rect 12551 3014 12576 3070
rect 12632 3014 12657 3070
rect 12713 3014 12738 3070
rect 12794 3014 12820 3070
rect 12876 3014 12901 3070
rect 12957 3014 12982 3070
rect 13038 3014 13063 3070
rect 13119 3014 13144 3070
rect 13200 3014 13225 3070
rect 13281 3014 13306 3070
rect 13362 3014 13388 3070
rect 13444 3014 13469 3070
rect 13525 3014 13550 3070
rect 13606 3014 13631 3070
rect 13687 3014 13712 3070
rect 13768 3014 13793 3070
rect 13849 3014 13874 3070
rect 13930 3014 13956 3070
rect 14012 3014 14037 3070
rect 14093 3014 14118 3070
rect 14174 3014 14199 3070
rect 14255 3014 14280 3070
rect 14336 3014 14361 3070
rect 14417 3014 14442 3070
rect 14498 3014 14524 3070
rect 14580 3014 14605 3070
rect 14661 3014 14686 3070
rect 14742 3014 14767 3070
rect 14823 3014 14848 3070
rect 14904 3014 14929 3070
rect 14985 3014 15010 3070
rect 15066 3014 15092 3070
rect 15148 3014 15173 3070
rect 15229 3014 15254 3070
rect 15310 3014 15335 3070
rect 15391 3014 15416 3070
rect 15472 3014 15497 3070
rect 15553 3014 15578 3070
rect 15634 3014 15660 3070
rect 15716 3014 15741 3070
rect 15797 3014 15822 3070
rect 15878 3014 15903 3070
rect 15959 3014 15984 3070
rect 16040 3014 16065 3070
rect 16121 3014 16146 3070
rect 16202 3014 16228 3070
rect 16284 3014 16309 3070
rect 16365 3014 16390 3070
rect 16446 3014 16471 3070
rect 16527 3014 16552 3070
rect 16608 3014 16633 3070
rect 16689 3014 16714 3070
rect 16770 3014 16796 3070
rect 16852 3014 16877 3070
rect 16933 3014 16958 3070
rect 17014 3014 17039 3070
rect 17095 3014 17120 3070
rect 17176 3014 17201 3070
rect 17257 3014 17282 3070
rect 17338 3014 17364 3070
rect 17420 3014 17445 3070
rect 17501 3014 17526 3070
rect 17582 3014 17607 3070
rect 17663 3014 17688 3070
rect 17744 3014 17769 3070
rect 17825 3014 17850 3070
rect 17906 3014 17932 3070
rect 17988 3014 18013 3070
rect 18069 3014 18094 3070
rect 18150 3014 18175 3070
rect 18231 3014 18256 3070
rect 18312 3014 18337 3070
rect 18393 3014 18418 3070
rect 18474 3014 18500 3070
rect 18556 3014 18581 3070
rect 18637 3014 18662 3070
rect 18718 3014 18743 3070
rect 18799 3014 18824 3070
rect 18880 3014 18905 3070
rect 18961 3014 18986 3070
rect 19042 3014 19068 3070
rect 19124 3014 19149 3070
rect 19205 3014 19230 3070
rect 19286 3014 19311 3070
rect 19367 3014 19392 3070
rect 19448 3014 19473 3070
rect 19529 3014 19554 3070
rect 19610 3014 19636 3070
rect 19692 3014 19717 3070
rect 19773 3014 19798 3070
rect 19854 3014 19879 3070
rect 19935 3014 19960 3070
rect 20016 3014 20041 3070
rect 20097 3014 20122 3070
rect 20178 3014 20204 3070
rect 20260 3014 20285 3070
rect 20341 3014 20366 3070
rect 20422 3014 20447 3070
rect 20503 3014 20528 3070
rect 20584 3014 20609 3070
rect 20665 3014 20690 3070
rect 20746 3014 20772 3070
rect 20828 3014 20853 3070
rect 20909 3014 20934 3070
rect 20990 3014 21015 3070
rect 21071 3014 21096 3070
rect 21152 3014 21177 3070
rect 21233 3014 21258 3070
rect 21314 3014 21340 3070
rect 21396 3014 21421 3070
rect 21477 3014 21502 3070
rect 21558 3014 21583 3070
rect 21639 3014 21664 3070
rect 21720 3014 21745 3070
rect 21801 3014 21826 3070
rect 21882 3014 21908 3070
rect 21964 3014 21989 3070
rect 22045 3014 22070 3070
rect 22126 3014 22151 3070
rect 22207 3014 22232 3070
rect 22288 3014 22313 3070
rect 22369 3014 22394 3070
rect 22450 3014 22476 3070
rect 22532 3014 22557 3070
rect 22613 3014 22638 3070
rect 22694 3014 22719 3070
rect 22775 3014 22800 3070
rect 22856 3014 22881 3070
rect 22937 3014 22962 3070
rect 23018 3014 23044 3070
rect 23100 3014 23125 3070
rect 23181 3014 23206 3070
rect 23262 3014 23287 3070
rect 23343 3014 23368 3070
rect 23424 3014 23449 3070
rect 23505 3014 23530 3070
rect 23586 3014 23612 3070
rect 23668 3014 23693 3070
rect 23749 3014 23774 3070
rect 23830 3014 23855 3070
rect 23911 3014 23936 3070
rect 23992 3014 24017 3070
rect 24073 3014 24098 3070
rect 24154 3014 24180 3070
rect 24236 3014 24261 3070
rect 24317 3014 24342 3070
rect 24398 3014 24423 3070
rect 24479 3014 24504 3070
rect 24560 3014 24585 3070
rect 24641 3014 24666 3070
rect 24722 3014 25067 3070
rect 3012 2966 25067 3014
rect 3012 2910 3036 2966
rect 3092 2910 3118 2966
rect 3174 2910 3199 2966
rect 3255 2910 3280 2966
rect 3336 2910 3361 2966
rect 3417 2910 3442 2966
rect 3498 2910 3523 2966
rect 3579 2910 3604 2966
rect 3660 2910 3686 2966
rect 3742 2910 3767 2966
rect 3823 2910 3848 2966
rect 3904 2910 3929 2966
rect 3985 2910 4010 2966
rect 4066 2910 4091 2966
rect 4147 2910 4172 2966
rect 4228 2910 4254 2966
rect 4310 2910 4335 2966
rect 4391 2910 4416 2966
rect 4472 2910 4497 2966
rect 4553 2910 4578 2966
rect 4634 2910 4659 2966
rect 4715 2910 4740 2966
rect 4796 2910 4822 2966
rect 4878 2910 4903 2966
rect 4959 2910 4984 2966
rect 5040 2910 5065 2966
rect 5121 2910 5146 2966
rect 5202 2910 5227 2966
rect 5283 2910 5308 2966
rect 5364 2910 5390 2966
rect 5446 2910 5471 2966
rect 5527 2910 5552 2966
rect 5608 2910 5633 2966
rect 5689 2910 5714 2966
rect 5770 2910 5795 2966
rect 5851 2910 5876 2966
rect 5932 2910 5958 2966
rect 6014 2910 6039 2966
rect 6095 2910 6120 2966
rect 6176 2910 6201 2966
rect 6257 2910 6282 2966
rect 6338 2910 6363 2966
rect 6419 2910 6444 2966
rect 6500 2910 6526 2966
rect 6582 2910 6607 2966
rect 6663 2910 6688 2966
rect 6744 2910 6769 2966
rect 6825 2910 6850 2966
rect 6906 2910 6931 2966
rect 6987 2910 7012 2966
rect 7068 2910 7094 2966
rect 7150 2910 7175 2966
rect 7231 2910 7256 2966
rect 7312 2910 7337 2966
rect 7393 2910 7418 2966
rect 7474 2910 7499 2966
rect 7555 2910 7580 2966
rect 7636 2910 7662 2966
rect 7718 2910 7743 2966
rect 7799 2910 7824 2966
rect 7880 2910 7905 2966
rect 7961 2910 7986 2966
rect 8042 2910 8067 2966
rect 8123 2910 8148 2966
rect 8204 2910 8230 2966
rect 8286 2910 8311 2966
rect 8367 2910 8392 2966
rect 8448 2910 8473 2966
rect 8529 2910 8554 2966
rect 8610 2910 8635 2966
rect 8691 2910 8716 2966
rect 8772 2910 8798 2966
rect 8854 2910 8879 2966
rect 8935 2910 8960 2966
rect 9016 2910 9041 2966
rect 9097 2910 9122 2966
rect 9178 2910 9203 2966
rect 9259 2910 9284 2966
rect 9340 2910 9366 2966
rect 9422 2910 9447 2966
rect 9503 2910 9528 2966
rect 9584 2910 9609 2966
rect 9665 2910 9690 2966
rect 9746 2910 9771 2966
rect 9827 2910 9852 2966
rect 9908 2910 9934 2966
rect 9990 2910 10015 2966
rect 10071 2910 10096 2966
rect 10152 2910 10177 2966
rect 10233 2910 10258 2966
rect 10314 2910 10339 2966
rect 10395 2910 10420 2966
rect 10476 2910 10502 2966
rect 10558 2910 10583 2966
rect 10639 2910 10664 2966
rect 10720 2910 10745 2966
rect 10801 2910 10826 2966
rect 10882 2910 10907 2966
rect 10963 2910 10988 2966
rect 11044 2910 11116 2966
rect 11172 2910 11197 2966
rect 11253 2910 11278 2966
rect 11334 2910 11359 2966
rect 11415 2910 11440 2966
rect 11496 2910 11521 2966
rect 11577 2910 11602 2966
rect 11658 2910 11684 2966
rect 11740 2910 11765 2966
rect 11821 2910 11846 2966
rect 11902 2910 11927 2966
rect 11983 2910 12008 2966
rect 12064 2910 12089 2966
rect 12145 2910 12170 2966
rect 12226 2910 12252 2966
rect 12308 2910 12333 2966
rect 12389 2910 12414 2966
rect 12470 2910 12495 2966
rect 12551 2910 12576 2966
rect 12632 2910 12657 2966
rect 12713 2910 12738 2966
rect 12794 2910 12820 2966
rect 12876 2910 12901 2966
rect 12957 2910 12982 2966
rect 13038 2910 13063 2966
rect 13119 2910 13144 2966
rect 13200 2910 13225 2966
rect 13281 2910 13306 2966
rect 13362 2910 13388 2966
rect 13444 2910 13469 2966
rect 13525 2910 13550 2966
rect 13606 2910 13631 2966
rect 13687 2910 13712 2966
rect 13768 2910 13793 2966
rect 13849 2910 13874 2966
rect 13930 2910 13956 2966
rect 14012 2910 14037 2966
rect 14093 2910 14118 2966
rect 14174 2910 14199 2966
rect 14255 2910 14280 2966
rect 14336 2910 14361 2966
rect 14417 2910 14442 2966
rect 14498 2910 14524 2966
rect 14580 2910 14605 2966
rect 14661 2910 14686 2966
rect 14742 2910 14767 2966
rect 14823 2910 14848 2966
rect 14904 2910 14929 2966
rect 14985 2910 15010 2966
rect 15066 2910 15092 2966
rect 15148 2910 15173 2966
rect 15229 2910 15254 2966
rect 15310 2910 15335 2966
rect 15391 2910 15416 2966
rect 15472 2910 15497 2966
rect 15553 2910 15578 2966
rect 15634 2910 15660 2966
rect 15716 2910 15741 2966
rect 15797 2910 15822 2966
rect 15878 2910 15903 2966
rect 15959 2910 15984 2966
rect 16040 2910 16065 2966
rect 16121 2910 16146 2966
rect 16202 2910 16228 2966
rect 16284 2910 16309 2966
rect 16365 2910 16390 2966
rect 16446 2910 16471 2966
rect 16527 2910 16552 2966
rect 16608 2910 16633 2966
rect 16689 2910 16714 2966
rect 16770 2910 16796 2966
rect 16852 2910 16877 2966
rect 16933 2910 16958 2966
rect 17014 2910 17039 2966
rect 17095 2910 17120 2966
rect 17176 2910 17201 2966
rect 17257 2910 17282 2966
rect 17338 2910 17364 2966
rect 17420 2910 17445 2966
rect 17501 2910 17526 2966
rect 17582 2910 17607 2966
rect 17663 2910 17688 2966
rect 17744 2910 17769 2966
rect 17825 2910 17850 2966
rect 17906 2910 17932 2966
rect 17988 2910 18013 2966
rect 18069 2910 18094 2966
rect 18150 2910 18175 2966
rect 18231 2910 18256 2966
rect 18312 2910 18337 2966
rect 18393 2910 18418 2966
rect 18474 2910 18500 2966
rect 18556 2910 18581 2966
rect 18637 2910 18662 2966
rect 18718 2910 18743 2966
rect 18799 2910 18824 2966
rect 18880 2910 18905 2966
rect 18961 2910 18986 2966
rect 19042 2910 19068 2966
rect 19124 2910 19149 2966
rect 19205 2910 19230 2966
rect 19286 2910 19311 2966
rect 19367 2910 19392 2966
rect 19448 2910 19473 2966
rect 19529 2910 19554 2966
rect 19610 2910 19636 2966
rect 19692 2910 19717 2966
rect 19773 2910 19798 2966
rect 19854 2910 19879 2966
rect 19935 2910 19960 2966
rect 20016 2910 20041 2966
rect 20097 2910 20122 2966
rect 20178 2910 20204 2966
rect 20260 2910 20285 2966
rect 20341 2910 20366 2966
rect 20422 2910 20447 2966
rect 20503 2910 20528 2966
rect 20584 2910 20609 2966
rect 20665 2910 20690 2966
rect 20746 2910 20772 2966
rect 20828 2910 20853 2966
rect 20909 2910 20934 2966
rect 20990 2910 21015 2966
rect 21071 2910 21096 2966
rect 21152 2910 21177 2966
rect 21233 2910 21258 2966
rect 21314 2910 21340 2966
rect 21396 2910 21421 2966
rect 21477 2910 21502 2966
rect 21558 2910 21583 2966
rect 21639 2910 21664 2966
rect 21720 2910 21745 2966
rect 21801 2910 21826 2966
rect 21882 2910 21908 2966
rect 21964 2910 21989 2966
rect 22045 2910 22070 2966
rect 22126 2910 22151 2966
rect 22207 2910 22232 2966
rect 22288 2910 22313 2966
rect 22369 2910 22394 2966
rect 22450 2910 22476 2966
rect 22532 2910 22557 2966
rect 22613 2910 22638 2966
rect 22694 2910 22719 2966
rect 22775 2910 22800 2966
rect 22856 2910 22881 2966
rect 22937 2910 22962 2966
rect 23018 2910 23044 2966
rect 23100 2910 23125 2966
rect 23181 2910 23206 2966
rect 23262 2910 23287 2966
rect 23343 2910 23368 2966
rect 23424 2910 23449 2966
rect 23505 2910 23530 2966
rect 23586 2910 23612 2966
rect 23668 2910 23693 2966
rect 23749 2910 23774 2966
rect 23830 2910 23855 2966
rect 23911 2910 23936 2966
rect 23992 2910 24017 2966
rect 24073 2910 24098 2966
rect 24154 2910 24180 2966
rect 24236 2910 24261 2966
rect 24317 2910 24342 2966
rect 24398 2910 24423 2966
rect 24479 2910 24504 2966
rect 24560 2910 24585 2966
rect 24641 2910 24666 2966
rect 24722 2910 25067 2966
rect 3012 2905 25067 2910
rect 4919 2667 4971 2677
rect 4919 2054 4971 2107
rect 5155 2667 5207 2677
rect 5155 2054 5207 2107
rect 5391 2667 5443 2677
rect 5391 2054 5443 2107
rect 5627 2667 5679 2677
rect 5627 2054 5679 2107
rect 5863 2667 5915 2677
rect 5863 2054 5915 2107
rect 6099 2667 6151 2677
rect 6099 2054 6151 2107
rect 6335 2667 6387 2677
rect 6335 2054 6387 2107
rect 6571 2667 6623 2677
rect 6571 2054 6623 2107
rect 6915 2667 6971 2677
rect 6915 2097 6971 2107
rect 7151 2667 7207 2677
rect 7151 2097 7207 2107
rect 7387 2667 7443 2677
rect 7387 2097 7443 2107
rect 7623 2667 7679 2677
rect 7623 2097 7679 2107
rect 7859 2667 7915 2677
rect 7859 2097 7915 2107
rect 8095 2667 8151 2677
rect 8095 2097 8151 2107
rect 8331 2667 8387 2677
rect 8331 2097 8387 2107
rect 8567 2667 8623 2677
rect 8567 2097 8623 2107
rect 8913 2667 8969 2677
rect 8913 2097 8969 2107
rect 9149 2667 9205 2677
rect 9149 2097 9205 2107
rect 9385 2667 9441 2677
rect 9385 2097 9441 2107
rect 9621 2667 9677 2677
rect 9621 2097 9677 2107
rect 9857 2667 9913 2677
rect 9857 2097 9913 2107
rect 10093 2667 10149 2677
rect 10093 2097 10149 2107
rect 10329 2667 10385 2677
rect 10329 2097 10385 2107
rect 10565 2667 10621 2677
rect 10565 2097 10621 2107
rect 12491 2666 12543 2905
rect 12491 2096 12543 2106
rect 12607 2666 12663 2676
rect 12607 2096 12663 2106
rect 12727 2666 12779 2905
rect 12727 2096 12779 2106
rect 12843 2666 12899 2676
rect 12843 2096 12899 2106
rect 12963 2666 13015 2905
rect 12963 2096 13015 2106
rect 13079 2666 13135 2676
rect 13079 2096 13135 2106
rect 13199 2666 13251 2905
rect 13199 2096 13251 2106
rect 13315 2666 13371 2676
rect 13315 2096 13371 2106
rect 13435 2666 13487 2905
rect 13435 2096 13487 2106
rect 13551 2666 13607 2676
rect 13551 2096 13607 2106
rect 13671 2666 13723 2905
rect 13671 2096 13723 2106
rect 13787 2666 13843 2676
rect 13787 2096 13843 2106
rect 13907 2666 13959 2905
rect 13907 2096 13959 2106
rect 14023 2666 14079 2676
rect 14023 2096 14079 2106
rect 14143 2666 14195 2905
rect 14143 2096 14195 2106
rect 14259 2666 14315 2676
rect 14259 2096 14315 2106
rect 14379 2666 14431 2905
rect 14379 2096 14431 2106
rect 14495 2666 14551 2676
rect 14495 2096 14551 2106
rect 14615 2666 14667 2905
rect 14615 2096 14667 2106
rect 14731 2666 14787 2676
rect 14731 2096 14787 2106
rect 14851 2666 14903 2905
rect 14851 2096 14903 2106
rect 14967 2666 15023 2676
rect 14967 2096 15023 2106
rect 15087 2666 15139 2905
rect 15087 2096 15139 2106
rect 15203 2666 15259 2676
rect 15203 2096 15259 2106
rect 15323 2666 15375 2905
rect 15323 2096 15375 2106
rect 15439 2666 15495 2676
rect 15439 2096 15495 2106
rect 16614 2666 16666 2905
rect 16614 2096 16666 2106
rect 16730 2666 16786 2676
rect 16730 2096 16786 2106
rect 16850 2666 16902 2905
rect 16850 2096 16902 2106
rect 16966 2666 17022 2676
rect 16966 2096 17022 2106
rect 17086 2666 17138 2905
rect 17086 2096 17138 2106
rect 17202 2666 17258 2676
rect 17202 2096 17258 2106
rect 17322 2666 17374 2905
rect 17322 2096 17374 2106
rect 17438 2666 17494 2676
rect 17438 2096 17494 2106
rect 17558 2666 17610 2905
rect 17558 2096 17610 2106
rect 17674 2666 17730 2676
rect 17674 2096 17730 2106
rect 17794 2666 17846 2905
rect 17794 2096 17846 2106
rect 17910 2666 17966 2676
rect 17910 2096 17966 2106
rect 18030 2666 18082 2905
rect 18030 2096 18082 2106
rect 18146 2666 18202 2676
rect 18146 2096 18202 2106
rect 18266 2666 18318 2905
rect 18266 2096 18318 2106
rect 18382 2666 18438 2676
rect 18382 2096 18438 2106
rect 18502 2666 18554 2905
rect 18502 2096 18554 2106
rect 18618 2666 18674 2676
rect 18618 2096 18674 2106
rect 18738 2666 18790 2905
rect 18738 2096 18790 2106
rect 18854 2666 18910 2676
rect 18854 2096 18910 2106
rect 18974 2666 19026 2905
rect 18974 2096 19026 2106
rect 19090 2666 19146 2676
rect 19090 2096 19146 2106
rect 19210 2666 19262 2905
rect 19210 2096 19262 2106
rect 19326 2666 19382 2676
rect 19326 2096 19382 2106
rect 19446 2666 19498 2905
rect 19446 2096 19498 2106
rect 19562 2666 19618 2676
rect 19562 2096 19618 2106
rect 20737 2666 20789 2905
rect 20737 2096 20789 2106
rect 20853 2666 20909 2676
rect 20853 2096 20909 2106
rect 20973 2666 21025 2905
rect 20973 2096 21025 2106
rect 21089 2666 21145 2676
rect 21089 2096 21145 2106
rect 21209 2666 21261 2905
rect 21209 2096 21261 2106
rect 21325 2666 21381 2676
rect 21325 2096 21381 2106
rect 21445 2666 21497 2905
rect 21445 2096 21497 2106
rect 21561 2666 21617 2676
rect 21561 2096 21617 2106
rect 21681 2666 21733 2905
rect 21681 2096 21733 2106
rect 21797 2666 21853 2676
rect 21797 2096 21853 2106
rect 21917 2666 21969 2905
rect 21917 2096 21969 2106
rect 22033 2666 22089 2676
rect 22033 2096 22089 2106
rect 22153 2666 22205 2905
rect 22153 2096 22205 2106
rect 22269 2666 22325 2676
rect 22269 2096 22325 2106
rect 22389 2666 22441 2905
rect 22389 2096 22441 2106
rect 22505 2666 22561 2676
rect 22505 2096 22561 2106
rect 22625 2666 22677 2905
rect 22625 2096 22677 2106
rect 22741 2666 22797 2676
rect 22741 2096 22797 2106
rect 22861 2666 22913 2905
rect 22861 2096 22913 2106
rect 22977 2666 23033 2676
rect 22977 2096 23033 2106
rect 23097 2666 23149 2905
rect 23097 2096 23149 2106
rect 23213 2666 23269 2676
rect 23213 2096 23269 2106
rect 23333 2666 23385 2905
rect 23333 2096 23385 2106
rect 23449 2666 23505 2676
rect 23449 2096 23505 2106
rect 23569 2666 23621 2905
rect 23569 2096 23621 2106
rect 23685 2666 23741 2676
rect 23903 2667 25067 2905
rect 23685 2096 23741 2106
rect 23895 2653 25067 2667
rect 23947 2601 23975 2653
rect 24027 2601 24055 2653
rect 24107 2601 24135 2653
rect 24187 2601 24215 2653
rect 24267 2601 24295 2653
rect 24347 2601 24375 2653
rect 24427 2601 24455 2653
rect 24507 2601 24535 2653
rect 24587 2601 24615 2653
rect 24667 2601 24695 2653
rect 24747 2601 24775 2653
rect 24827 2601 24855 2653
rect 24907 2601 24935 2653
rect 24987 2601 25015 2653
rect 23895 2573 25067 2601
rect 23947 2521 23975 2573
rect 24027 2521 24055 2573
rect 24107 2521 24135 2573
rect 24187 2521 24215 2573
rect 24267 2521 24295 2573
rect 24347 2521 24375 2573
rect 24427 2521 24455 2573
rect 24507 2521 24535 2573
rect 24587 2521 24615 2573
rect 24667 2521 24695 2573
rect 24747 2521 24775 2573
rect 24827 2521 24855 2573
rect 24907 2521 24935 2573
rect 24987 2521 25015 2573
rect 23895 2493 25067 2521
rect 23947 2441 23975 2493
rect 24027 2441 24055 2493
rect 24107 2441 24135 2493
rect 24187 2441 24215 2493
rect 24267 2441 24295 2493
rect 24347 2441 24375 2493
rect 24427 2441 24455 2493
rect 24507 2441 24535 2493
rect 24587 2441 24615 2493
rect 24667 2441 24695 2493
rect 24747 2441 24775 2493
rect 24827 2441 24855 2493
rect 24907 2441 24935 2493
rect 24987 2441 25015 2493
rect 23895 2413 25067 2441
rect 23947 2361 23975 2413
rect 24027 2361 24055 2413
rect 24107 2361 24135 2413
rect 24187 2361 24215 2413
rect 24267 2361 24295 2413
rect 24347 2361 24375 2413
rect 24427 2361 24455 2413
rect 24507 2361 24535 2413
rect 24587 2361 24615 2413
rect 24667 2361 24695 2413
rect 24747 2361 24775 2413
rect 24827 2361 24855 2413
rect 24907 2361 24935 2413
rect 24987 2361 25015 2413
rect 23895 2333 25067 2361
rect 23947 2281 23975 2333
rect 24027 2281 24055 2333
rect 24107 2281 24135 2333
rect 24187 2281 24215 2333
rect 24267 2281 24295 2333
rect 24347 2281 24375 2333
rect 24427 2281 24455 2333
rect 24507 2281 24535 2333
rect 24587 2281 24615 2333
rect 24667 2281 24695 2333
rect 24747 2281 24775 2333
rect 24827 2281 24855 2333
rect 24907 2281 24935 2333
rect 24987 2281 25015 2333
rect 23895 2253 25067 2281
rect 23947 2201 23975 2253
rect 24027 2201 24055 2253
rect 24107 2201 24135 2253
rect 24187 2201 24215 2253
rect 24267 2201 24295 2253
rect 24347 2201 24375 2253
rect 24427 2201 24455 2253
rect 24507 2201 24535 2253
rect 24587 2201 24615 2253
rect 24667 2201 24695 2253
rect 24747 2201 24775 2253
rect 24827 2201 24855 2253
rect 24907 2201 24935 2253
rect 24987 2201 25015 2253
rect 23895 2173 25067 2201
rect 23947 2121 23975 2173
rect 24027 2121 24055 2173
rect 24107 2121 24135 2173
rect 24187 2121 24215 2173
rect 24267 2121 24295 2173
rect 24347 2121 24375 2173
rect 24427 2121 24455 2173
rect 24507 2121 24535 2173
rect 24587 2121 24615 2173
rect 24667 2121 24695 2173
rect 24747 2121 24775 2173
rect 24827 2121 24855 2173
rect 24907 2121 24935 2173
rect 24987 2121 25015 2173
rect 23895 2093 25067 2121
rect 2069 2045 23720 2054
rect 2069 2044 12547 2045
rect 2069 1952 4857 2044
rect 4915 1952 4975 2044
rect 5033 1952 5093 2044
rect 5151 1952 5211 2044
rect 5269 1952 5329 2044
rect 5387 1952 5447 2044
rect 5505 1952 5565 2044
rect 5623 1952 5683 2044
rect 5741 1952 5801 2044
rect 5859 1952 5919 2044
rect 5977 1952 6037 2044
rect 6095 1952 6155 2044
rect 6213 1952 6273 2044
rect 6331 1952 6391 2044
rect 6449 1952 6509 2044
rect 6567 1952 6855 2044
rect 6913 1952 6973 2044
rect 7031 1952 7091 2044
rect 7149 1952 7209 2044
rect 7267 1952 7327 2044
rect 7385 1952 7445 2044
rect 7503 1952 7563 2044
rect 7621 1952 7681 2044
rect 7739 1952 7799 2044
rect 7857 1952 7917 2044
rect 7975 1952 8035 2044
rect 8093 1952 8153 2044
rect 8211 1952 8271 2044
rect 8329 1952 8389 2044
rect 8447 1952 8507 2044
rect 8565 1952 8853 2044
rect 8911 1952 8971 2044
rect 9029 1952 9089 2044
rect 9147 1952 9207 2044
rect 9265 1952 9325 2044
rect 9383 1952 9443 2044
rect 9501 1952 9561 2044
rect 9619 1952 9679 2044
rect 9737 1952 9797 2044
rect 9855 1952 9915 2044
rect 9973 1952 10033 2044
rect 10091 1952 10151 2044
rect 10209 1952 10269 2044
rect 10327 1952 10387 2044
rect 10445 1952 10505 2044
rect 10563 1952 12547 2044
rect 2069 1891 12547 1952
rect 12605 1891 12665 2045
rect 12723 1891 12783 2045
rect 12841 1891 12901 2045
rect 12959 1891 13019 2045
rect 13077 1891 13137 2045
rect 13195 1891 13255 2045
rect 13313 1891 13373 2045
rect 13431 1891 13491 2045
rect 13549 1891 13609 2045
rect 13667 1891 13727 2045
rect 13785 1891 13845 2045
rect 13903 1891 13963 2045
rect 14021 1891 14081 2045
rect 14139 1891 14199 2045
rect 14257 1891 14317 2045
rect 14375 1891 14435 2045
rect 14493 1891 14553 2045
rect 14611 1891 14671 2045
rect 14729 1891 14789 2045
rect 14847 1891 14907 2045
rect 14965 1891 15025 2045
rect 15083 1891 15143 2045
rect 15201 1891 15261 2045
rect 15319 1891 15379 2045
rect 15437 1891 16670 2045
rect 16728 1891 16788 2045
rect 16846 1891 16906 2045
rect 16964 1891 17024 2045
rect 17082 1891 17142 2045
rect 17200 1891 17260 2045
rect 17318 1891 17378 2045
rect 17436 1891 17496 2045
rect 17554 1891 17614 2045
rect 17672 1891 17732 2045
rect 17790 1891 17850 2045
rect 17908 1891 17968 2045
rect 18026 1891 18086 2045
rect 18144 1891 18204 2045
rect 18262 1891 18322 2045
rect 18380 1891 18440 2045
rect 18498 1891 18558 2045
rect 18616 1891 18676 2045
rect 18734 1891 18794 2045
rect 18852 1891 18912 2045
rect 18970 1891 19030 2045
rect 19088 1891 19148 2045
rect 19206 1891 19266 2045
rect 19324 1891 19384 2045
rect 19442 1891 19502 2045
rect 19560 1891 20793 2045
rect 20851 1891 20911 2045
rect 20969 1891 21029 2045
rect 21087 1891 21147 2045
rect 21205 1891 21265 2045
rect 21323 1891 21383 2045
rect 21441 1891 21501 2045
rect 21559 1891 21619 2045
rect 21677 1891 21737 2045
rect 21795 1891 21855 2045
rect 21913 1891 21973 2045
rect 22031 1891 22091 2045
rect 22149 1891 22209 2045
rect 22267 1891 22327 2045
rect 22385 1891 22445 2045
rect 22503 1891 22563 2045
rect 22621 1891 22681 2045
rect 22739 1891 22799 2045
rect 22857 1891 22917 2045
rect 22975 1891 23035 2045
rect 23093 1891 23153 2045
rect 23211 1891 23271 2045
rect 23329 1891 23389 2045
rect 23447 1891 23507 2045
rect 23565 1891 23625 2045
rect 23683 1891 23720 2045
rect 2069 1881 23720 1891
rect 23947 2041 23975 2093
rect 24027 2041 24055 2093
rect 24107 2041 24135 2093
rect 24187 2041 24215 2093
rect 24267 2041 24295 2093
rect 24347 2041 24375 2093
rect 24427 2041 24455 2093
rect 24507 2041 24535 2093
rect 24587 2041 24615 2093
rect 24667 2041 24695 2093
rect 24747 2041 24775 2093
rect 24827 2041 24855 2093
rect 24907 2041 24935 2093
rect 24987 2041 25015 2093
rect 23895 2013 25067 2041
rect 23947 1961 23975 2013
rect 24027 1961 24055 2013
rect 24107 1961 24135 2013
rect 24187 1961 24215 2013
rect 24267 1961 24295 2013
rect 24347 1961 24375 2013
rect 24427 1961 24455 2013
rect 24507 1961 24535 2013
rect 24587 1961 24615 2013
rect 24667 1961 24695 2013
rect 24747 1961 24775 2013
rect 24827 1961 24855 2013
rect 24907 1961 24935 2013
rect 24987 1961 25015 2013
rect 23895 1933 25067 1961
rect 23947 1881 23975 1933
rect 24027 1881 24055 1933
rect 24107 1881 24135 1933
rect 24187 1881 24215 1933
rect 24267 1881 24295 1933
rect 24347 1881 24375 1933
rect 24427 1881 24455 1933
rect 24507 1881 24535 1933
rect 24587 1881 24615 1933
rect 24667 1881 24695 1933
rect 24747 1881 24775 1933
rect 24827 1881 24855 1933
rect 24907 1881 24935 1933
rect 24987 1881 25015 1933
rect 23895 1853 25067 1881
rect 12491 1830 12543 1840
rect 4760 1593 11628 1601
rect 4760 1537 4775 1593
rect 4831 1569 4856 1593
rect 4853 1537 4856 1569
rect 4912 1537 4937 1593
rect 4993 1537 5018 1593
rect 5074 1569 5099 1593
rect 5089 1537 5099 1569
rect 5155 1537 5180 1593
rect 5236 1537 5261 1593
rect 5317 1569 5363 1593
rect 5325 1537 5363 1569
rect 5419 1537 5444 1593
rect 5500 1569 5525 1593
rect 5500 1537 5509 1569
rect 5581 1537 5606 1593
rect 5662 1537 5687 1593
rect 5743 1569 5768 1593
rect 5743 1537 5745 1569
rect 5824 1537 5849 1593
rect 5905 1537 5951 1593
rect 6007 1569 6032 1593
rect 6088 1537 6113 1593
rect 6169 1537 6194 1593
rect 6250 1569 6275 1593
rect 6269 1537 6275 1569
rect 6331 1537 6356 1593
rect 6412 1537 6437 1593
rect 6493 1569 6517 1593
rect 6505 1537 6517 1569
rect 6573 1537 6598 1593
rect 6654 1537 6679 1593
rect 6735 1569 6760 1593
rect 6741 1537 6760 1569
rect 6816 1537 6841 1593
rect 6897 1537 6922 1593
rect 6978 1537 7003 1593
rect 7059 1537 7090 1593
rect 7146 1569 7171 1593
rect 7146 1537 7161 1569
rect 7227 1537 7252 1593
rect 7308 1537 7333 1593
rect 7389 1569 7414 1593
rect 7389 1537 7397 1569
rect 7470 1537 7495 1593
rect 7551 1537 7576 1593
rect 7632 1569 7656 1593
rect 7632 1537 7633 1569
rect 7712 1537 7737 1593
rect 7793 1537 7818 1593
rect 7874 1569 7899 1593
rect 7955 1537 7980 1593
rect 8036 1537 8061 1593
rect 8117 1569 8142 1593
rect 8198 1537 8222 1593
rect 8278 1537 8303 1593
rect 8359 1569 8384 1593
rect 8440 1537 8465 1593
rect 8521 1537 8546 1593
rect 8602 1569 8627 1593
rect 8683 1537 8708 1593
rect 8764 1537 8788 1593
rect 8844 1569 8869 1593
rect 8865 1537 8869 1569
rect 8925 1537 8950 1593
rect 9006 1537 9031 1593
rect 9087 1569 9112 1593
rect 9101 1537 9112 1569
rect 9168 1537 9193 1593
rect 9249 1537 9274 1593
rect 9330 1569 9357 1593
rect 9337 1537 9357 1569
rect 9413 1537 9438 1593
rect 9494 1537 9519 1593
rect 9575 1537 9600 1593
rect 9656 1537 9681 1593
rect 9737 1569 9762 1593
rect 9737 1537 9757 1569
rect 9818 1537 9843 1593
rect 9899 1537 9923 1593
rect 9979 1569 10004 1593
rect 9979 1537 9993 1569
rect 10060 1537 10085 1593
rect 10141 1537 10166 1593
rect 10222 1569 10247 1593
rect 10222 1537 10229 1569
rect 10303 1537 10328 1593
rect 10384 1537 10409 1593
rect 10465 1569 10489 1593
rect 10545 1537 10570 1593
rect 10626 1537 10651 1593
rect 10707 1569 10732 1593
rect 10788 1537 10813 1593
rect 10869 1537 10894 1593
rect 10950 1537 10975 1593
rect 11031 1537 11055 1593
rect 11111 1537 11136 1593
rect 11192 1537 11217 1593
rect 11273 1537 11298 1593
rect 11354 1537 11379 1593
rect 11435 1537 11460 1593
rect 11516 1537 11541 1593
rect 11597 1537 11628 1593
rect 4760 1489 4801 1537
rect 4853 1489 5037 1537
rect 5089 1489 5273 1537
rect 5325 1489 5509 1537
rect 5561 1489 5745 1537
rect 5797 1489 5981 1537
rect 6033 1489 6217 1537
rect 6269 1489 6453 1537
rect 6505 1489 6689 1537
rect 6741 1489 6925 1537
rect 6977 1489 7161 1537
rect 7213 1489 7397 1537
rect 7449 1489 7633 1537
rect 7685 1489 7869 1537
rect 7921 1489 8105 1537
rect 8157 1489 8341 1537
rect 8393 1489 8577 1537
rect 8629 1489 8813 1537
rect 8865 1489 9049 1537
rect 9101 1489 9285 1537
rect 9337 1489 9521 1537
rect 9573 1489 9757 1537
rect 9809 1489 9993 1537
rect 10045 1489 10229 1537
rect 10281 1489 10465 1537
rect 10517 1489 10701 1537
rect 10753 1489 11628 1537
rect 4760 1433 4775 1489
rect 4853 1433 4856 1489
rect 4912 1433 4937 1489
rect 4993 1433 5018 1489
rect 5089 1433 5099 1489
rect 5155 1433 5180 1489
rect 5236 1433 5261 1489
rect 5325 1433 5363 1489
rect 5419 1433 5444 1489
rect 5500 1433 5509 1489
rect 5581 1433 5606 1489
rect 5662 1433 5687 1489
rect 5743 1433 5745 1489
rect 5824 1433 5849 1489
rect 5905 1433 5951 1489
rect 6088 1433 6113 1489
rect 6169 1433 6194 1489
rect 6269 1433 6275 1489
rect 6331 1433 6356 1489
rect 6412 1433 6437 1489
rect 6505 1433 6517 1489
rect 6573 1433 6598 1489
rect 6654 1433 6679 1489
rect 6741 1433 6760 1489
rect 6816 1433 6841 1489
rect 6897 1433 6922 1489
rect 6978 1433 7003 1489
rect 7059 1433 7090 1489
rect 7146 1433 7161 1489
rect 7227 1433 7252 1489
rect 7308 1433 7333 1489
rect 7389 1433 7397 1489
rect 7470 1433 7495 1489
rect 7551 1433 7576 1489
rect 7632 1433 7633 1489
rect 7712 1433 7737 1489
rect 7793 1433 7818 1489
rect 7955 1433 7980 1489
rect 8036 1433 8061 1489
rect 8198 1433 8222 1489
rect 8278 1433 8303 1489
rect 8440 1433 8465 1489
rect 8521 1433 8546 1489
rect 8683 1433 8708 1489
rect 8764 1433 8788 1489
rect 8865 1433 8869 1489
rect 8925 1433 8950 1489
rect 9006 1433 9031 1489
rect 9101 1433 9112 1489
rect 9168 1433 9193 1489
rect 9249 1433 9274 1489
rect 9337 1433 9357 1489
rect 9413 1433 9438 1489
rect 9494 1433 9519 1489
rect 9575 1433 9600 1489
rect 9656 1433 9681 1489
rect 9737 1433 9757 1489
rect 9818 1433 9843 1489
rect 9899 1433 9923 1489
rect 9979 1433 9993 1489
rect 10060 1433 10085 1489
rect 10141 1433 10166 1489
rect 10222 1433 10229 1489
rect 10303 1433 10328 1489
rect 10384 1433 10409 1489
rect 10545 1433 10570 1489
rect 10626 1433 10651 1489
rect 10788 1433 10813 1489
rect 10869 1433 10894 1489
rect 10950 1433 10975 1489
rect 11031 1433 11055 1489
rect 11111 1433 11136 1489
rect 11192 1433 11217 1489
rect 11273 1433 11298 1489
rect 11354 1433 11379 1489
rect 11435 1433 11460 1489
rect 11516 1433 11541 1489
rect 11597 1433 11628 1489
rect 4760 1385 4801 1433
rect 4853 1385 5037 1433
rect 5089 1385 5273 1433
rect 5325 1385 5509 1433
rect 5561 1385 5745 1433
rect 5797 1385 5981 1433
rect 6033 1385 6217 1433
rect 6269 1385 6453 1433
rect 6505 1385 6689 1433
rect 6741 1385 6925 1433
rect 6977 1385 7161 1433
rect 7213 1385 7397 1433
rect 7449 1385 7633 1433
rect 7685 1385 7869 1433
rect 7921 1385 8105 1433
rect 8157 1385 8341 1433
rect 8393 1385 8577 1433
rect 8629 1385 8813 1433
rect 8865 1385 9049 1433
rect 9101 1385 9285 1433
rect 9337 1385 9521 1433
rect 9573 1385 9757 1433
rect 9809 1385 9993 1433
rect 10045 1385 10229 1433
rect 10281 1385 10465 1433
rect 10517 1385 10701 1433
rect 10753 1385 11628 1433
rect 4760 1329 4775 1385
rect 4853 1329 4856 1385
rect 4912 1329 4937 1385
rect 4993 1329 5018 1385
rect 5089 1329 5099 1385
rect 5155 1329 5180 1385
rect 5236 1329 5261 1385
rect 5325 1329 5363 1385
rect 5419 1329 5444 1385
rect 5500 1329 5509 1385
rect 5581 1329 5606 1385
rect 5662 1329 5687 1385
rect 5743 1329 5745 1385
rect 5824 1329 5849 1385
rect 5905 1329 5951 1385
rect 6088 1329 6113 1385
rect 6169 1329 6194 1385
rect 6269 1329 6275 1385
rect 6331 1329 6356 1385
rect 6412 1329 6437 1385
rect 6505 1329 6517 1385
rect 6573 1329 6598 1385
rect 6654 1329 6679 1385
rect 6741 1329 6760 1385
rect 6816 1329 6841 1385
rect 6897 1329 6922 1385
rect 6978 1329 7003 1385
rect 7059 1329 7090 1385
rect 7146 1329 7161 1385
rect 7227 1329 7252 1385
rect 7308 1329 7333 1385
rect 7389 1329 7397 1385
rect 7470 1329 7495 1385
rect 7551 1329 7576 1385
rect 7632 1329 7633 1385
rect 7712 1329 7737 1385
rect 7793 1329 7818 1385
rect 7955 1329 7980 1385
rect 8036 1329 8061 1385
rect 8198 1329 8222 1385
rect 8278 1329 8303 1385
rect 8440 1329 8465 1385
rect 8521 1329 8546 1385
rect 8683 1329 8708 1385
rect 8764 1329 8788 1385
rect 8865 1329 8869 1385
rect 8925 1329 8950 1385
rect 9006 1329 9031 1385
rect 9101 1329 9112 1385
rect 9168 1329 9193 1385
rect 9249 1329 9274 1385
rect 9337 1329 9357 1385
rect 9413 1329 9438 1385
rect 9494 1329 9519 1385
rect 9575 1329 9600 1385
rect 9656 1329 9681 1385
rect 9737 1329 9757 1385
rect 9818 1329 9843 1385
rect 9899 1329 9923 1385
rect 9979 1329 9993 1385
rect 10060 1329 10085 1385
rect 10141 1329 10166 1385
rect 10222 1329 10229 1385
rect 10303 1329 10328 1385
rect 10384 1329 10409 1385
rect 10545 1329 10570 1385
rect 10626 1329 10651 1385
rect 10788 1329 10813 1385
rect 10869 1329 10894 1385
rect 10950 1329 10975 1385
rect 11031 1329 11055 1385
rect 11111 1329 11136 1385
rect 11192 1329 11217 1385
rect 11273 1329 11298 1385
rect 11354 1329 11379 1385
rect 11435 1329 11460 1385
rect 11516 1329 11541 1385
rect 11597 1329 11628 1385
rect 4760 1319 4801 1329
rect 4853 1319 5037 1329
rect 5089 1319 5273 1329
rect 5325 1319 5509 1329
rect 5561 1319 5745 1329
rect 5797 1319 5981 1329
rect 6033 1319 6217 1329
rect 6269 1319 6453 1329
rect 6505 1319 6689 1329
rect 6741 1319 6925 1329
rect 6977 1319 7161 1329
rect 7213 1319 7397 1329
rect 7449 1319 7633 1329
rect 7685 1319 7869 1329
rect 7921 1319 8105 1329
rect 8157 1319 8341 1329
rect 8393 1319 8577 1329
rect 8629 1319 8813 1329
rect 8865 1319 9049 1329
rect 9101 1319 9285 1329
rect 9337 1319 9521 1329
rect 9573 1319 9757 1329
rect 9809 1319 9993 1329
rect 10045 1319 10229 1329
rect 10281 1319 10465 1329
rect 10517 1319 10701 1329
rect 10753 1319 11628 1329
rect 4801 1170 4853 1319
rect 4801 600 4853 610
rect 4915 1170 4971 1180
rect 4915 600 4971 610
rect 5037 1170 5089 1319
rect 5037 600 5089 610
rect 5151 1170 5207 1180
rect 5151 600 5207 610
rect 5273 1170 5325 1319
rect 5273 600 5325 610
rect 5387 1170 5443 1180
rect 5387 600 5443 610
rect 5509 1170 5561 1319
rect 5509 600 5561 610
rect 5623 1170 5679 1180
rect 5623 600 5679 610
rect 5745 1170 5797 1319
rect 5745 600 5797 610
rect 5859 1170 5915 1180
rect 5859 600 5915 610
rect 5981 1170 6033 1319
rect 5981 600 6033 610
rect 6095 1170 6151 1180
rect 6095 600 6151 610
rect 6217 1170 6269 1319
rect 6217 600 6269 610
rect 6331 1170 6387 1180
rect 6331 600 6387 610
rect 6453 1170 6505 1319
rect 6453 600 6505 610
rect 6567 1170 6623 1180
rect 6567 600 6623 610
rect 6689 1170 6741 1319
rect 6689 600 6741 610
rect 6803 1170 6859 1180
rect 6803 600 6859 610
rect 6925 1170 6977 1319
rect 6925 600 6977 610
rect 7039 1170 7095 1180
rect 7039 600 7095 610
rect 7161 1170 7213 1319
rect 7161 600 7213 610
rect 7275 1170 7331 1180
rect 7275 600 7331 610
rect 7397 1170 7449 1319
rect 7397 600 7449 610
rect 7511 1170 7567 1180
rect 7511 600 7567 610
rect 7633 1170 7685 1319
rect 7633 600 7685 610
rect 7747 1170 7803 1180
rect 7747 600 7803 610
rect 7869 1170 7921 1319
rect 7869 600 7921 610
rect 7983 1170 8039 1180
rect 7983 600 8039 610
rect 8105 1170 8157 1319
rect 8105 600 8157 610
rect 8219 1170 8275 1180
rect 8219 600 8275 610
rect 8341 1170 8393 1319
rect 8341 600 8393 610
rect 8455 1170 8511 1180
rect 8455 600 8511 610
rect 8577 1170 8629 1319
rect 8577 600 8629 610
rect 8691 1170 8747 1180
rect 8691 600 8747 610
rect 8813 1170 8865 1319
rect 8813 600 8865 610
rect 8927 1170 8983 1180
rect 8927 600 8983 610
rect 9049 1170 9101 1319
rect 9049 600 9101 610
rect 9163 1170 9219 1180
rect 9163 600 9219 610
rect 9285 1170 9337 1319
rect 9285 600 9337 610
rect 9399 1170 9455 1180
rect 9399 600 9455 610
rect 9521 1170 9573 1319
rect 9521 600 9573 610
rect 9635 1170 9691 1180
rect 9635 600 9691 610
rect 9757 1170 9809 1319
rect 9757 600 9809 610
rect 9871 1170 9927 1180
rect 9871 600 9927 610
rect 9993 1170 10045 1319
rect 9993 600 10045 610
rect 10107 1170 10163 1180
rect 10107 600 10163 610
rect 10229 1170 10281 1319
rect 10229 600 10281 610
rect 10343 1170 10399 1180
rect 10343 600 10399 610
rect 10465 1170 10517 1319
rect 10465 600 10517 610
rect 10579 1170 10635 1180
rect 10579 600 10635 610
rect 10701 1170 10753 1319
rect 10701 600 10753 610
rect 4136 556 4857 557
rect 4136 549 10697 556
rect 4136 395 4857 549
rect 4915 395 4975 549
rect 5033 395 5093 549
rect 5151 395 5211 549
rect 5269 395 5329 549
rect 5387 395 5447 549
rect 5505 395 5565 549
rect 5623 395 5683 549
rect 5741 395 5801 549
rect 5859 395 5919 549
rect 5977 395 6037 549
rect 6095 395 6155 549
rect 6213 395 6273 549
rect 6331 395 6391 549
rect 6449 395 6509 549
rect 6567 395 6627 549
rect 6685 395 6745 549
rect 6803 395 6863 549
rect 6921 395 6981 549
rect 7039 395 7099 549
rect 7157 395 7217 549
rect 7275 395 7335 549
rect 7393 395 7453 549
rect 7511 395 7571 549
rect 7629 395 7689 549
rect 7747 395 7807 549
rect 7865 395 7925 549
rect 7983 395 8043 549
rect 8101 395 8161 549
rect 8219 395 8279 549
rect 8337 395 8397 549
rect 8455 395 8515 549
rect 8573 395 8633 549
rect 8691 395 8751 549
rect 8809 395 8869 549
rect 8927 395 8987 549
rect 9045 395 9105 549
rect 9163 395 9223 549
rect 9281 395 9341 549
rect 9399 395 9459 549
rect 9517 395 9577 549
rect 9635 395 9695 549
rect 9753 395 9813 549
rect 9871 395 9931 549
rect 9989 395 10049 549
rect 10107 395 10167 549
rect 10225 395 10285 549
rect 10343 395 10403 549
rect 10461 395 10521 549
rect 10579 395 10639 549
rect 4136 389 10697 395
rect 4136 -429 4304 389
rect 4801 334 4853 344
rect 4801 -375 4853 -226
rect 4915 334 4971 344
rect 4915 -236 4971 -226
rect 5037 334 5089 344
rect 5037 -375 5089 -226
rect 5151 334 5207 344
rect 5151 -236 5207 -226
rect 5273 334 5325 344
rect 5273 -375 5325 -226
rect 5387 334 5443 344
rect 5387 -236 5443 -226
rect 5509 334 5561 344
rect 5509 -375 5561 -226
rect 5623 334 5679 344
rect 5623 -236 5679 -226
rect 5745 334 5797 344
rect 5745 -375 5797 -226
rect 5859 334 5915 344
rect 5859 -236 5915 -226
rect 5981 334 6033 344
rect 5981 -375 6033 -226
rect 6095 334 6151 344
rect 6095 -236 6151 -226
rect 6217 334 6269 344
rect 6217 -375 6269 -226
rect 6331 334 6387 344
rect 6331 -236 6387 -226
rect 6453 334 6505 344
rect 6453 -375 6505 -226
rect 6567 334 6623 344
rect 6567 -236 6623 -226
rect 6689 334 6741 344
rect 6689 -375 6741 -226
rect 6803 334 6859 344
rect 6803 -236 6859 -226
rect 6925 334 6977 344
rect 6925 -375 6977 -226
rect 7039 334 7095 344
rect 7039 -236 7095 -226
rect 7161 334 7213 344
rect 7161 -375 7213 -226
rect 7275 334 7331 344
rect 7275 -236 7331 -226
rect 7397 334 7449 344
rect 7397 -375 7449 -226
rect 7511 334 7567 344
rect 7511 -236 7567 -226
rect 7633 334 7685 344
rect 7633 -375 7685 -226
rect 7747 334 7803 344
rect 7747 -236 7803 -226
rect 7869 334 7921 344
rect 7869 -375 7921 -226
rect 7983 334 8039 344
rect 7983 -236 8039 -226
rect 8105 334 8157 344
rect 8105 -375 8157 -226
rect 8219 334 8275 344
rect 8219 -236 8275 -226
rect 8341 334 8393 344
rect 8341 -375 8393 -226
rect 8455 334 8511 344
rect 8455 -236 8511 -226
rect 8577 334 8629 344
rect 8577 -375 8629 -226
rect 8691 334 8747 344
rect 8691 -236 8747 -226
rect 8813 334 8865 344
rect 8813 -375 8865 -226
rect 8927 334 8983 344
rect 8927 -236 8983 -226
rect 9049 334 9101 344
rect 9049 -375 9101 -226
rect 9163 334 9219 344
rect 9163 -236 9219 -226
rect 9285 334 9337 344
rect 9285 -375 9337 -226
rect 9399 334 9455 344
rect 9399 -236 9455 -226
rect 9521 334 9573 344
rect 9521 -375 9573 -226
rect 9635 334 9691 344
rect 9635 -236 9691 -226
rect 9757 334 9809 344
rect 9757 -375 9809 -226
rect 9871 334 9927 344
rect 9871 -236 9927 -226
rect 9993 334 10045 344
rect 9993 -375 10045 -226
rect 10107 334 10163 344
rect 10107 -236 10163 -226
rect 10229 334 10281 344
rect 10229 -375 10281 -226
rect 10343 334 10399 344
rect 10343 -236 10399 -226
rect 10465 334 10517 344
rect 10465 -375 10517 -226
rect 10579 334 10635 344
rect 10579 -236 10635 -226
rect 10701 334 10753 344
rect 10701 -375 10753 -226
rect 10841 -375 11612 1319
rect 12491 1163 12543 1270
rect 12607 1830 12663 1840
rect 12607 1260 12663 1270
rect 12727 1830 12779 1840
rect 12727 1163 12779 1270
rect 12843 1830 12899 1840
rect 12843 1260 12899 1270
rect 12963 1830 13015 1840
rect 12963 1163 13015 1270
rect 13079 1830 13135 1840
rect 13079 1260 13135 1270
rect 13199 1830 13251 1840
rect 13199 1163 13251 1270
rect 13315 1830 13371 1840
rect 13315 1260 13371 1270
rect 13435 1830 13487 1840
rect 13435 1163 13487 1270
rect 13551 1830 13607 1840
rect 13551 1260 13607 1270
rect 13671 1830 13723 1840
rect 13671 1163 13723 1270
rect 13787 1830 13843 1840
rect 13787 1260 13843 1270
rect 13907 1830 13959 1840
rect 13907 1163 13959 1270
rect 14023 1830 14079 1840
rect 14023 1260 14079 1270
rect 14143 1830 14195 1840
rect 14143 1163 14195 1270
rect 14259 1830 14315 1840
rect 14259 1260 14315 1270
rect 14379 1830 14431 1840
rect 14379 1163 14431 1270
rect 14495 1830 14551 1840
rect 14495 1260 14551 1270
rect 14615 1830 14667 1840
rect 14615 1163 14667 1270
rect 14731 1830 14787 1840
rect 14731 1260 14787 1270
rect 14851 1830 14903 1840
rect 14851 1163 14903 1270
rect 14967 1830 15023 1840
rect 14967 1260 15023 1270
rect 15087 1830 15139 1840
rect 15087 1163 15139 1270
rect 15203 1830 15259 1840
rect 15203 1260 15259 1270
rect 15323 1830 15375 1840
rect 15323 1163 15375 1270
rect 15439 1830 15495 1840
rect 15439 1260 15495 1270
rect 16614 1830 16666 1840
rect 16614 1163 16666 1270
rect 16730 1830 16786 1840
rect 16730 1260 16786 1270
rect 16850 1830 16902 1840
rect 16850 1163 16902 1270
rect 16966 1830 17022 1840
rect 16966 1260 17022 1270
rect 17086 1830 17138 1840
rect 17086 1163 17138 1270
rect 17202 1830 17258 1840
rect 17202 1260 17258 1270
rect 17322 1830 17374 1840
rect 17322 1163 17374 1270
rect 17438 1830 17494 1840
rect 17438 1260 17494 1270
rect 17558 1830 17610 1840
rect 17558 1163 17610 1270
rect 17674 1830 17730 1840
rect 17674 1260 17730 1270
rect 17794 1830 17846 1840
rect 17794 1163 17846 1270
rect 17910 1830 17966 1840
rect 17910 1260 17966 1270
rect 18030 1830 18082 1840
rect 18030 1163 18082 1270
rect 18146 1830 18202 1840
rect 18146 1260 18202 1270
rect 18266 1830 18318 1840
rect 18266 1163 18318 1270
rect 18382 1830 18438 1840
rect 18382 1260 18438 1270
rect 18502 1830 18554 1840
rect 18502 1163 18554 1270
rect 18618 1830 18674 1840
rect 18618 1260 18674 1270
rect 18738 1830 18790 1840
rect 18738 1163 18790 1270
rect 18854 1830 18910 1840
rect 18854 1260 18910 1270
rect 18974 1830 19026 1840
rect 18974 1163 19026 1270
rect 19090 1830 19146 1840
rect 19090 1260 19146 1270
rect 19210 1830 19262 1840
rect 19210 1163 19262 1270
rect 19326 1830 19382 1840
rect 19326 1260 19382 1270
rect 19446 1830 19498 1840
rect 19446 1163 19498 1270
rect 19562 1830 19618 1840
rect 19562 1260 19618 1270
rect 20737 1830 20789 1840
rect 20737 1163 20789 1270
rect 20853 1830 20909 1840
rect 20853 1260 20909 1270
rect 20973 1830 21025 1840
rect 20973 1163 21025 1270
rect 21089 1830 21145 1840
rect 21089 1260 21145 1270
rect 21209 1830 21261 1840
rect 21209 1163 21261 1270
rect 21325 1830 21381 1840
rect 21325 1260 21381 1270
rect 21445 1830 21497 1840
rect 21445 1163 21497 1270
rect 21561 1830 21617 1840
rect 21561 1260 21617 1270
rect 21681 1830 21733 1840
rect 21681 1163 21733 1270
rect 21797 1830 21853 1840
rect 21797 1260 21853 1270
rect 21917 1830 21969 1840
rect 21917 1163 21969 1270
rect 22033 1830 22089 1840
rect 22033 1260 22089 1270
rect 22153 1830 22205 1840
rect 22153 1163 22205 1270
rect 22269 1830 22325 1840
rect 22269 1260 22325 1270
rect 22389 1830 22441 1840
rect 22389 1163 22441 1270
rect 22505 1830 22561 1840
rect 22505 1260 22561 1270
rect 22625 1830 22677 1840
rect 22625 1163 22677 1270
rect 22741 1830 22797 1840
rect 22741 1260 22797 1270
rect 22861 1830 22913 1840
rect 22861 1163 22913 1270
rect 22977 1830 23033 1840
rect 22977 1260 23033 1270
rect 23097 1830 23149 1840
rect 23097 1163 23149 1270
rect 23213 1830 23269 1840
rect 23213 1260 23269 1270
rect 23333 1830 23385 1840
rect 23333 1163 23385 1270
rect 23449 1830 23505 1840
rect 23449 1260 23505 1270
rect 23569 1830 23621 1840
rect 23569 1163 23621 1270
rect 23685 1830 23741 1840
rect 23685 1260 23741 1270
rect 23947 1801 23975 1853
rect 24027 1801 24055 1853
rect 24107 1801 24135 1853
rect 24187 1801 24215 1853
rect 24267 1801 24295 1853
rect 24347 1801 24375 1853
rect 24427 1801 24455 1853
rect 24507 1801 24535 1853
rect 24587 1801 24615 1853
rect 24667 1801 24695 1853
rect 24747 1801 24775 1853
rect 24827 1801 24855 1853
rect 24907 1801 24935 1853
rect 24987 1801 25015 1853
rect 23895 1773 25067 1801
rect 23947 1721 23975 1773
rect 24027 1721 24055 1773
rect 24107 1721 24135 1773
rect 24187 1721 24215 1773
rect 24267 1721 24295 1773
rect 24347 1721 24375 1773
rect 24427 1721 24455 1773
rect 24507 1721 24535 1773
rect 24587 1721 24615 1773
rect 24667 1721 24695 1773
rect 24747 1721 24775 1773
rect 24827 1721 24855 1773
rect 24907 1721 24935 1773
rect 24987 1721 25015 1773
rect 23895 1693 25067 1721
rect 23947 1641 23975 1693
rect 24027 1641 24055 1693
rect 24107 1641 24135 1693
rect 24187 1641 24215 1693
rect 24267 1641 24295 1693
rect 24347 1641 24375 1693
rect 24427 1641 24455 1693
rect 24507 1641 24535 1693
rect 24587 1641 24615 1693
rect 24667 1641 24695 1693
rect 24747 1641 24775 1693
rect 24827 1641 24855 1693
rect 24907 1641 24935 1693
rect 24987 1641 25015 1693
rect 23895 1613 25067 1641
rect 23947 1561 23975 1613
rect 24027 1561 24055 1613
rect 24107 1561 24135 1613
rect 24187 1561 24215 1613
rect 24267 1561 24295 1613
rect 24347 1561 24375 1613
rect 24427 1561 24455 1613
rect 24507 1561 24535 1613
rect 24587 1561 24615 1613
rect 24667 1561 24695 1613
rect 24747 1561 24775 1613
rect 24827 1561 24855 1613
rect 24907 1561 24935 1613
rect 24987 1561 25015 1613
rect 23895 1533 25067 1561
rect 23947 1481 23975 1533
rect 24027 1481 24055 1533
rect 24107 1481 24135 1533
rect 24187 1481 24215 1533
rect 24267 1481 24295 1533
rect 24347 1481 24375 1533
rect 24427 1481 24455 1533
rect 24507 1481 24535 1533
rect 24587 1481 24615 1533
rect 24667 1481 24695 1533
rect 24747 1481 24775 1533
rect 24827 1481 24855 1533
rect 24907 1481 24935 1533
rect 24987 1481 25015 1533
rect 23895 1453 25067 1481
rect 23947 1401 23975 1453
rect 24027 1401 24055 1453
rect 24107 1401 24135 1453
rect 24187 1401 24215 1453
rect 24267 1401 24295 1453
rect 24347 1401 24375 1453
rect 24427 1401 24455 1453
rect 24507 1401 24535 1453
rect 24587 1401 24615 1453
rect 24667 1401 24695 1453
rect 24747 1401 24775 1453
rect 24827 1401 24855 1453
rect 24907 1401 24935 1453
rect 24987 1401 25015 1453
rect 23895 1373 25067 1401
rect 23947 1321 23975 1373
rect 24027 1321 24055 1373
rect 24107 1321 24135 1373
rect 24187 1321 24215 1373
rect 24267 1321 24295 1373
rect 24347 1321 24375 1373
rect 24427 1321 24455 1373
rect 24507 1321 24535 1373
rect 24587 1321 24615 1373
rect 24667 1321 24695 1373
rect 24747 1321 24775 1373
rect 24827 1321 24855 1373
rect 24907 1321 24935 1373
rect 24987 1321 25015 1373
rect 23895 1293 25067 1321
rect 23947 1241 23975 1293
rect 24027 1241 24055 1293
rect 24107 1241 24135 1293
rect 24187 1241 24215 1293
rect 24267 1241 24295 1293
rect 24347 1241 24375 1293
rect 24427 1241 24455 1293
rect 24507 1241 24535 1293
rect 24587 1241 24615 1293
rect 24667 1241 24695 1293
rect 24747 1241 24775 1293
rect 24827 1241 24855 1293
rect 24907 1241 24935 1293
rect 24987 1241 25015 1293
rect 23895 1227 25067 1241
rect 23903 1163 25067 1227
rect 12485 1149 25067 1163
rect 12537 1097 12565 1149
rect 12617 1097 12645 1149
rect 12697 1097 12725 1149
rect 12777 1097 12805 1149
rect 12857 1097 12885 1149
rect 12937 1097 12965 1149
rect 13017 1097 13045 1149
rect 13097 1097 13125 1149
rect 13177 1097 13205 1149
rect 13257 1097 13285 1149
rect 13337 1097 13365 1149
rect 13417 1097 13445 1149
rect 13497 1097 13525 1149
rect 13577 1097 13605 1149
rect 13657 1097 13685 1149
rect 13737 1097 13765 1149
rect 13817 1097 13845 1149
rect 13897 1097 13925 1149
rect 13977 1097 14005 1149
rect 14057 1097 14085 1149
rect 14137 1097 14165 1149
rect 14217 1097 14245 1149
rect 14297 1097 14325 1149
rect 14377 1097 14405 1149
rect 14457 1097 14485 1149
rect 14537 1097 14565 1149
rect 14617 1097 14645 1149
rect 14697 1097 14725 1149
rect 14777 1097 14805 1149
rect 14857 1097 14885 1149
rect 14937 1097 14965 1149
rect 15017 1097 15045 1149
rect 15097 1097 15125 1149
rect 15177 1097 15205 1149
rect 15257 1097 15285 1149
rect 15337 1097 15365 1149
rect 15417 1097 15445 1149
rect 15497 1097 15525 1149
rect 15577 1097 15605 1149
rect 15657 1097 15685 1149
rect 15737 1097 15765 1149
rect 15817 1097 15845 1149
rect 15897 1097 15925 1149
rect 15977 1097 16005 1149
rect 16057 1097 16085 1149
rect 16137 1097 16165 1149
rect 16217 1097 16245 1149
rect 16297 1097 16325 1149
rect 16377 1097 16405 1149
rect 16457 1097 16485 1149
rect 16537 1097 16565 1149
rect 16617 1097 16645 1149
rect 16697 1097 16725 1149
rect 16777 1097 16805 1149
rect 16857 1097 16885 1149
rect 16937 1097 16965 1149
rect 17017 1097 17045 1149
rect 17097 1097 17125 1149
rect 17177 1097 17205 1149
rect 17257 1097 17285 1149
rect 17337 1097 17365 1149
rect 17417 1097 17445 1149
rect 17497 1097 17525 1149
rect 17577 1097 17605 1149
rect 17657 1097 17685 1149
rect 17737 1097 17765 1149
rect 17817 1097 17845 1149
rect 17897 1097 17925 1149
rect 17977 1097 18005 1149
rect 18057 1097 18085 1149
rect 18137 1097 18165 1149
rect 18217 1097 18245 1149
rect 18297 1097 18325 1149
rect 18377 1097 18405 1149
rect 18457 1097 18485 1149
rect 18537 1097 18565 1149
rect 18617 1097 18645 1149
rect 18697 1097 18725 1149
rect 18777 1097 18805 1149
rect 18857 1097 18885 1149
rect 18937 1097 18965 1149
rect 19017 1097 19045 1149
rect 19097 1097 19125 1149
rect 19177 1097 19205 1149
rect 19257 1097 19285 1149
rect 19337 1097 19365 1149
rect 19417 1097 19445 1149
rect 19497 1097 19525 1149
rect 19577 1097 19605 1149
rect 19657 1097 19685 1149
rect 19737 1097 19765 1149
rect 19817 1097 19845 1149
rect 19897 1097 19925 1149
rect 19977 1097 20005 1149
rect 20057 1097 20085 1149
rect 20137 1097 20165 1149
rect 20217 1097 20245 1149
rect 20297 1097 20325 1149
rect 20377 1097 20405 1149
rect 20457 1097 20485 1149
rect 20537 1097 20565 1149
rect 20617 1097 20645 1149
rect 20697 1097 20725 1149
rect 20777 1097 20805 1149
rect 20857 1097 20885 1149
rect 20937 1097 20965 1149
rect 21017 1097 21045 1149
rect 21097 1097 21125 1149
rect 21177 1097 21205 1149
rect 21257 1097 21285 1149
rect 21337 1097 21365 1149
rect 21417 1097 21445 1149
rect 21497 1097 21525 1149
rect 21577 1097 21605 1149
rect 21657 1097 21685 1149
rect 21737 1097 21765 1149
rect 21817 1097 21845 1149
rect 21897 1097 21925 1149
rect 21977 1097 22005 1149
rect 22057 1097 22085 1149
rect 22137 1097 22165 1149
rect 22217 1097 22245 1149
rect 22297 1097 22325 1149
rect 22377 1097 22405 1149
rect 22457 1097 22485 1149
rect 22537 1097 22565 1149
rect 22617 1097 22645 1149
rect 22697 1097 22725 1149
rect 22777 1097 22805 1149
rect 22857 1097 22885 1149
rect 22937 1097 22965 1149
rect 23017 1097 23045 1149
rect 23097 1097 23125 1149
rect 23177 1097 23205 1149
rect 23257 1097 23285 1149
rect 23337 1097 23365 1149
rect 23417 1097 23445 1149
rect 23497 1097 23525 1149
rect 23577 1097 23605 1149
rect 23657 1097 23685 1149
rect 23737 1097 23765 1149
rect 23817 1097 23845 1149
rect 23897 1097 23925 1149
rect 23977 1097 24005 1149
rect 24057 1097 24085 1149
rect 24137 1097 24165 1149
rect 24217 1097 24245 1149
rect 24297 1097 24325 1149
rect 24377 1097 24405 1149
rect 24457 1097 25067 1149
rect 12485 1069 25067 1097
rect 12537 1017 12565 1069
rect 12617 1017 12645 1069
rect 12697 1017 12725 1069
rect 12777 1017 12805 1069
rect 12857 1017 12885 1069
rect 12937 1017 12965 1069
rect 13017 1017 13045 1069
rect 13097 1017 13125 1069
rect 13177 1017 13205 1069
rect 13257 1017 13285 1069
rect 13337 1017 13365 1069
rect 13417 1017 13445 1069
rect 13497 1017 13525 1069
rect 13577 1017 13605 1069
rect 13657 1017 13685 1069
rect 13737 1017 13765 1069
rect 13817 1017 13845 1069
rect 13897 1017 13925 1069
rect 13977 1017 14005 1069
rect 14057 1017 14085 1069
rect 14137 1017 14165 1069
rect 14217 1017 14245 1069
rect 14297 1017 14325 1069
rect 14377 1017 14405 1069
rect 14457 1017 14485 1069
rect 14537 1017 14565 1069
rect 14617 1017 14645 1069
rect 14697 1017 14725 1069
rect 14777 1017 14805 1069
rect 14857 1017 14885 1069
rect 14937 1017 14965 1069
rect 15017 1017 15045 1069
rect 15097 1017 15125 1069
rect 15177 1017 15205 1069
rect 15257 1017 15285 1069
rect 15337 1017 15365 1069
rect 15417 1017 15445 1069
rect 15497 1017 15525 1069
rect 15577 1017 15605 1069
rect 15657 1017 15685 1069
rect 15737 1017 15765 1069
rect 15817 1017 15845 1069
rect 15897 1017 15925 1069
rect 15977 1017 16005 1069
rect 16057 1017 16085 1069
rect 16137 1017 16165 1069
rect 16217 1017 16245 1069
rect 16297 1017 16325 1069
rect 16377 1017 16405 1069
rect 16457 1017 16485 1069
rect 16537 1017 16565 1069
rect 16617 1017 16645 1069
rect 16697 1017 16725 1069
rect 16777 1017 16805 1069
rect 16857 1017 16885 1069
rect 16937 1017 16965 1069
rect 17017 1017 17045 1069
rect 17097 1017 17125 1069
rect 17177 1017 17205 1069
rect 17257 1017 17285 1069
rect 17337 1017 17365 1069
rect 17417 1017 17445 1069
rect 17497 1017 17525 1069
rect 17577 1017 17605 1069
rect 17657 1017 17685 1069
rect 17737 1017 17765 1069
rect 17817 1017 17845 1069
rect 17897 1017 17925 1069
rect 17977 1017 18005 1069
rect 18057 1017 18085 1069
rect 18137 1017 18165 1069
rect 18217 1017 18245 1069
rect 18297 1017 18325 1069
rect 18377 1017 18405 1069
rect 18457 1017 18485 1069
rect 18537 1017 18565 1069
rect 18617 1017 18645 1069
rect 18697 1017 18725 1069
rect 18777 1017 18805 1069
rect 18857 1017 18885 1069
rect 18937 1017 18965 1069
rect 19017 1017 19045 1069
rect 19097 1017 19125 1069
rect 19177 1017 19205 1069
rect 19257 1017 19285 1069
rect 19337 1017 19365 1069
rect 19417 1017 19445 1069
rect 19497 1017 19525 1069
rect 19577 1017 19605 1069
rect 19657 1017 19685 1069
rect 19737 1017 19765 1069
rect 19817 1017 19845 1069
rect 19897 1017 19925 1069
rect 19977 1017 20005 1069
rect 20057 1017 20085 1069
rect 20137 1017 20165 1069
rect 20217 1017 20245 1069
rect 20297 1017 20325 1069
rect 20377 1017 20405 1069
rect 20457 1017 20485 1069
rect 20537 1017 20565 1069
rect 20617 1017 20645 1069
rect 20697 1017 20725 1069
rect 20777 1017 20805 1069
rect 20857 1017 20885 1069
rect 20937 1017 20965 1069
rect 21017 1017 21045 1069
rect 21097 1017 21125 1069
rect 21177 1017 21205 1069
rect 21257 1017 21285 1069
rect 21337 1017 21365 1069
rect 21417 1017 21445 1069
rect 21497 1017 21525 1069
rect 21577 1017 21605 1069
rect 21657 1017 21685 1069
rect 21737 1017 21765 1069
rect 21817 1017 21845 1069
rect 21897 1017 21925 1069
rect 21977 1017 22005 1069
rect 22057 1017 22085 1069
rect 22137 1017 22165 1069
rect 22217 1017 22245 1069
rect 22297 1017 22325 1069
rect 22377 1017 22405 1069
rect 22457 1017 22485 1069
rect 22537 1017 22565 1069
rect 22617 1017 22645 1069
rect 22697 1017 22725 1069
rect 22777 1017 22805 1069
rect 22857 1017 22885 1069
rect 22937 1017 22965 1069
rect 23017 1017 23045 1069
rect 23097 1017 23125 1069
rect 23177 1017 23205 1069
rect 23257 1017 23285 1069
rect 23337 1017 23365 1069
rect 23417 1017 23445 1069
rect 23497 1017 23525 1069
rect 23577 1017 23605 1069
rect 23657 1017 23685 1069
rect 23737 1017 23765 1069
rect 23817 1017 23845 1069
rect 23897 1017 23925 1069
rect 23977 1017 24005 1069
rect 24057 1017 24085 1069
rect 24137 1017 24165 1069
rect 24217 1017 24245 1069
rect 24297 1017 24325 1069
rect 24377 1017 24405 1069
rect 24457 1017 25067 1069
rect 12485 1004 25067 1017
rect 12485 1003 24457 1004
rect 3032 -677 4304 -429
rect 4746 -625 4801 -375
rect 4853 -625 5037 -375
rect 5089 -625 5273 -375
rect 5325 -625 5509 -375
rect 5561 -625 5745 -375
rect 5797 -625 5981 -375
rect 6033 -625 6217 -375
rect 6269 -625 6453 -375
rect 6505 -625 6689 -375
rect 6741 -625 6925 -375
rect 6977 -625 7161 -375
rect 7213 -625 7397 -375
rect 7449 -625 7633 -375
rect 7685 -625 7869 -375
rect 7921 -625 8105 -375
rect 8157 -625 8341 -375
rect 8393 -625 8577 -375
rect 8629 -625 8813 -375
rect 8865 -625 9049 -375
rect 9101 -625 9285 -375
rect 9337 -625 9521 -375
rect 9573 -625 9757 -375
rect 9809 -625 9993 -375
rect 10045 -625 10229 -375
rect 10281 -625 10465 -375
rect 10517 -625 10701 -375
rect 10753 -625 11612 -375
rect 4746 -626 11612 -625
rect 4136 -1493 4304 -677
rect 4801 -880 4853 -626
rect 4801 -1450 4853 -1440
rect 4915 -880 4971 -870
rect 4915 -1450 4971 -1440
rect 5037 -880 5089 -626
rect 5037 -1450 5089 -1440
rect 5151 -880 5207 -870
rect 5151 -1450 5207 -1440
rect 5273 -880 5325 -626
rect 5273 -1450 5325 -1440
rect 5387 -880 5443 -870
rect 5387 -1450 5443 -1440
rect 5509 -880 5561 -626
rect 5509 -1450 5561 -1440
rect 5623 -880 5679 -870
rect 5623 -1450 5679 -1440
rect 5745 -880 5797 -626
rect 5745 -1450 5797 -1440
rect 5859 -880 5915 -870
rect 5859 -1450 5915 -1440
rect 5981 -880 6033 -626
rect 5981 -1450 6033 -1440
rect 6095 -880 6151 -870
rect 6095 -1450 6151 -1440
rect 6217 -880 6269 -626
rect 6217 -1450 6269 -1440
rect 6331 -880 6387 -870
rect 6331 -1450 6387 -1440
rect 6453 -880 6505 -626
rect 6453 -1450 6505 -1440
rect 6567 -880 6623 -870
rect 6567 -1450 6623 -1440
rect 6689 -880 6741 -626
rect 6689 -1450 6741 -1440
rect 6803 -880 6859 -870
rect 6803 -1450 6859 -1440
rect 6925 -880 6977 -626
rect 6925 -1450 6977 -1440
rect 7039 -880 7095 -870
rect 7039 -1450 7095 -1440
rect 7161 -880 7213 -626
rect 7161 -1450 7213 -1440
rect 7275 -880 7331 -870
rect 7275 -1450 7331 -1440
rect 7397 -880 7449 -626
rect 7397 -1450 7449 -1440
rect 7511 -880 7567 -870
rect 7511 -1450 7567 -1440
rect 7633 -880 7685 -626
rect 7633 -1450 7685 -1440
rect 7747 -880 7803 -870
rect 7747 -1450 7803 -1440
rect 7869 -880 7921 -626
rect 7869 -1450 7921 -1440
rect 7983 -880 8039 -870
rect 7983 -1450 8039 -1440
rect 8105 -880 8157 -626
rect 8105 -1450 8157 -1440
rect 8219 -880 8275 -870
rect 8219 -1450 8275 -1440
rect 8341 -880 8393 -626
rect 8341 -1450 8393 -1440
rect 8455 -880 8511 -870
rect 8455 -1450 8511 -1440
rect 8577 -880 8629 -626
rect 8577 -1450 8629 -1440
rect 8691 -880 8747 -870
rect 8691 -1450 8747 -1440
rect 8813 -880 8865 -626
rect 8813 -1450 8865 -1440
rect 8927 -880 8983 -870
rect 8927 -1450 8983 -1440
rect 9049 -880 9101 -626
rect 9049 -1450 9101 -1440
rect 9163 -880 9219 -870
rect 9163 -1450 9219 -1440
rect 9285 -880 9337 -626
rect 9285 -1450 9337 -1440
rect 9399 -880 9455 -870
rect 9399 -1450 9455 -1440
rect 9521 -880 9573 -626
rect 9521 -1450 9573 -1440
rect 9635 -880 9691 -870
rect 9635 -1450 9691 -1440
rect 9757 -880 9809 -626
rect 9757 -1450 9809 -1440
rect 9871 -880 9927 -870
rect 9871 -1450 9927 -1440
rect 9993 -880 10045 -626
rect 9993 -1450 10045 -1440
rect 10107 -880 10163 -870
rect 10107 -1450 10163 -1440
rect 10229 -880 10281 -626
rect 10229 -1450 10281 -1440
rect 10343 -880 10399 -870
rect 10343 -1450 10399 -1440
rect 10465 -880 10517 -626
rect 10465 -1450 10517 -1440
rect 10579 -880 10635 -870
rect 10579 -1450 10635 -1440
rect 10701 -880 10753 -626
rect 10701 -1450 10753 -1440
rect 4136 -1494 4857 -1493
rect 4136 -1501 10697 -1494
rect 4136 -1655 4857 -1501
rect 4915 -1655 4975 -1501
rect 5033 -1655 5093 -1501
rect 5151 -1655 5211 -1501
rect 5269 -1655 5329 -1501
rect 5387 -1655 5447 -1501
rect 5505 -1655 5565 -1501
rect 5623 -1655 5683 -1501
rect 5741 -1655 5801 -1501
rect 5859 -1655 5919 -1501
rect 5977 -1655 6037 -1501
rect 6095 -1655 6155 -1501
rect 6213 -1655 6273 -1501
rect 6331 -1655 6391 -1501
rect 6449 -1655 6509 -1501
rect 6567 -1655 6627 -1501
rect 6685 -1655 6745 -1501
rect 6803 -1655 6863 -1501
rect 6921 -1655 6981 -1501
rect 7039 -1655 7099 -1501
rect 7157 -1655 7217 -1501
rect 7275 -1655 7335 -1501
rect 7393 -1655 7453 -1501
rect 7511 -1655 7571 -1501
rect 7629 -1655 7689 -1501
rect 7747 -1655 7807 -1501
rect 7865 -1655 7925 -1501
rect 7983 -1655 8043 -1501
rect 8101 -1655 8161 -1501
rect 8219 -1655 8279 -1501
rect 8337 -1655 8397 -1501
rect 8455 -1655 8515 -1501
rect 8573 -1655 8633 -1501
rect 8691 -1655 8751 -1501
rect 8809 -1655 8869 -1501
rect 8927 -1655 8987 -1501
rect 9045 -1655 9105 -1501
rect 9163 -1655 9223 -1501
rect 9281 -1655 9341 -1501
rect 9399 -1655 9459 -1501
rect 9517 -1655 9577 -1501
rect 9635 -1655 9695 -1501
rect 9753 -1655 9813 -1501
rect 9871 -1655 9931 -1501
rect 9989 -1655 10049 -1501
rect 10107 -1655 10167 -1501
rect 10225 -1655 10285 -1501
rect 10343 -1655 10403 -1501
rect 10461 -1655 10521 -1501
rect 10579 -1655 10639 -1501
rect 4136 -1661 10697 -1655
rect 4801 -1716 4853 -1706
rect 4801 -2424 4853 -2276
rect 4915 -1716 4971 -1706
rect 4915 -2286 4971 -2276
rect 5037 -1716 5089 -1706
rect 5037 -2424 5089 -2276
rect 5151 -1716 5207 -1706
rect 5151 -2286 5207 -2276
rect 5273 -1716 5325 -1706
rect 5273 -2424 5325 -2276
rect 5387 -1716 5443 -1706
rect 5387 -2286 5443 -2276
rect 5509 -1716 5561 -1706
rect 5509 -2424 5561 -2276
rect 5623 -1716 5679 -1706
rect 5623 -2286 5679 -2276
rect 5745 -1716 5797 -1706
rect 5745 -2424 5797 -2276
rect 5859 -1716 5915 -1706
rect 5859 -2286 5915 -2276
rect 5981 -1716 6033 -1706
rect 5981 -2424 6033 -2276
rect 6095 -1716 6151 -1706
rect 6095 -2286 6151 -2276
rect 6217 -1716 6269 -1706
rect 6217 -2424 6269 -2276
rect 6331 -1716 6387 -1706
rect 6331 -2286 6387 -2276
rect 6453 -1716 6505 -1706
rect 6453 -2424 6505 -2276
rect 6567 -1716 6623 -1706
rect 6567 -2286 6623 -2276
rect 6689 -1716 6741 -1706
rect 6689 -2424 6741 -2276
rect 6803 -1716 6859 -1706
rect 6803 -2286 6859 -2276
rect 6925 -1716 6977 -1706
rect 6925 -2424 6977 -2276
rect 7039 -1716 7095 -1706
rect 7039 -2286 7095 -2276
rect 7161 -1716 7213 -1706
rect 7161 -2424 7213 -2276
rect 7275 -1716 7331 -1706
rect 7275 -2286 7331 -2276
rect 7397 -1716 7449 -1706
rect 7397 -2424 7449 -2276
rect 7511 -1716 7567 -1706
rect 7511 -2286 7567 -2276
rect 7633 -1716 7685 -1706
rect 7633 -2424 7685 -2276
rect 7747 -1716 7803 -1706
rect 7747 -2286 7803 -2276
rect 7869 -1716 7921 -1706
rect 7869 -2424 7921 -2276
rect 7983 -1716 8039 -1706
rect 7983 -2286 8039 -2276
rect 8105 -1716 8157 -1706
rect 8105 -2424 8157 -2276
rect 8219 -1716 8275 -1706
rect 8219 -2286 8275 -2276
rect 8341 -1716 8393 -1706
rect 8341 -2424 8393 -2276
rect 8455 -1716 8511 -1706
rect 8455 -2286 8511 -2276
rect 8577 -1716 8629 -1706
rect 8577 -2424 8629 -2276
rect 8691 -1716 8747 -1706
rect 8691 -2286 8747 -2276
rect 8813 -1716 8865 -1706
rect 8813 -2424 8865 -2276
rect 8927 -1716 8983 -1706
rect 8927 -2286 8983 -2276
rect 9049 -1716 9101 -1706
rect 9049 -2424 9101 -2276
rect 9163 -1716 9219 -1706
rect 9163 -2286 9219 -2276
rect 9285 -1716 9337 -1706
rect 9285 -2424 9337 -2276
rect 9399 -1716 9455 -1706
rect 9399 -2286 9455 -2276
rect 9521 -1716 9573 -1706
rect 9521 -2424 9573 -2276
rect 9635 -1716 9691 -1706
rect 9635 -2286 9691 -2276
rect 9757 -1716 9809 -1706
rect 9757 -2424 9809 -2276
rect 9871 -1716 9927 -1706
rect 9871 -2286 9927 -2276
rect 9993 -1716 10045 -1706
rect 9993 -2424 10045 -2276
rect 10107 -1716 10163 -1706
rect 10107 -2286 10163 -2276
rect 10229 -1716 10281 -1706
rect 10229 -2424 10281 -2276
rect 10343 -1716 10399 -1706
rect 10343 -2286 10399 -2276
rect 10465 -1716 10517 -1706
rect 10465 -2424 10517 -2276
rect 10579 -1716 10635 -1706
rect 10579 -2286 10635 -2276
rect 10701 -1716 10753 -1706
rect 10701 -2424 10753 -2276
rect 10841 -2424 11612 -626
rect 4746 -2425 11612 -2424
rect 4746 -2675 4801 -2425
rect 4853 -2675 5037 -2425
rect 5089 -2675 5273 -2425
rect 5325 -2675 5509 -2425
rect 5561 -2675 5745 -2425
rect 5797 -2675 5981 -2425
rect 6033 -2675 6217 -2425
rect 6269 -2675 6453 -2425
rect 6505 -2675 6689 -2425
rect 6741 -2675 6925 -2425
rect 6977 -2675 7161 -2425
rect 7213 -2675 7397 -2425
rect 7449 -2675 7633 -2425
rect 7685 -2675 7869 -2425
rect 7921 -2675 8105 -2425
rect 8157 -2675 8341 -2425
rect 8393 -2675 8577 -2425
rect 8629 -2675 8813 -2425
rect 8865 -2675 9049 -2425
rect 9101 -2675 9285 -2425
rect 9337 -2675 9521 -2425
rect 9573 -2675 9757 -2425
rect 9809 -2675 9993 -2425
rect 10045 -2675 10229 -2425
rect 10281 -2675 10465 -2425
rect 10517 -2675 10701 -2425
rect 10753 -2675 11612 -2425
rect 4801 -2930 4853 -2675
rect 4801 -3500 4853 -3490
rect 4919 -2930 4975 -2920
rect 4919 -3500 4975 -3490
rect 5037 -2930 5089 -2675
rect 5037 -3500 5089 -3490
rect 5155 -2930 5211 -2920
rect 5155 -3500 5211 -3490
rect 5273 -2930 5325 -2675
rect 5273 -3500 5325 -3490
rect 5391 -2930 5447 -2920
rect 5391 -3500 5447 -3490
rect 5509 -2930 5561 -2675
rect 5509 -3500 5561 -3490
rect 5627 -2930 5683 -2920
rect 5627 -3500 5683 -3490
rect 5745 -2930 5797 -2675
rect 5745 -3500 5797 -3490
rect 5863 -2930 5919 -2920
rect 5863 -3500 5919 -3490
rect 5981 -2930 6033 -2675
rect 5981 -3500 6033 -3490
rect 6099 -2930 6155 -2920
rect 6099 -3500 6155 -3490
rect 6217 -2930 6269 -2675
rect 6217 -3500 6269 -3490
rect 6335 -2930 6391 -2920
rect 6335 -3500 6391 -3490
rect 6453 -2930 6505 -2675
rect 6453 -3500 6505 -3490
rect 6571 -2930 6627 -2920
rect 6571 -3500 6627 -3490
rect 6689 -2930 6741 -2675
rect 6689 -3500 6741 -3490
rect 6807 -2930 6863 -2920
rect 6807 -3500 6863 -3490
rect 6925 -2930 6977 -2675
rect 6925 -3500 6977 -3490
rect 7043 -2930 7099 -2920
rect 7043 -3500 7099 -3490
rect 7161 -2930 7213 -2675
rect 7161 -3500 7213 -3490
rect 7279 -2930 7335 -2920
rect 7279 -3500 7335 -3490
rect 7397 -2930 7449 -2675
rect 7397 -3500 7449 -3490
rect 7515 -2930 7571 -2920
rect 7515 -3500 7571 -3490
rect 7633 -2930 7685 -2675
rect 7633 -3500 7685 -3490
rect 7751 -2930 7807 -2920
rect 7751 -3500 7807 -3490
rect 7869 -2930 7921 -2675
rect 7869 -3500 7921 -3490
rect 7987 -2930 8043 -2920
rect 7987 -3500 8043 -3490
rect 8105 -2930 8157 -2675
rect 8105 -3500 8157 -3490
rect 8223 -2930 8279 -2920
rect 8223 -3500 8279 -3490
rect 8341 -2930 8393 -2675
rect 8341 -3500 8393 -3490
rect 8459 -2930 8515 -2920
rect 8459 -3500 8515 -3490
rect 8577 -2930 8629 -2675
rect 8577 -3500 8629 -3490
rect 8695 -2930 8751 -2920
rect 8695 -3500 8751 -3490
rect 8813 -2930 8865 -2675
rect 8813 -3500 8865 -3490
rect 8931 -2930 8987 -2920
rect 8931 -3500 8987 -3490
rect 9049 -2930 9101 -2675
rect 9049 -3500 9101 -3490
rect 9167 -2930 9223 -2920
rect 9167 -3500 9223 -3490
rect 9285 -2930 9337 -2675
rect 9285 -3500 9337 -3490
rect 9403 -2930 9459 -2920
rect 9403 -3500 9459 -3490
rect 9521 -2930 9573 -2675
rect 9521 -3500 9573 -3490
rect 9639 -2930 9695 -2920
rect 9639 -3500 9695 -3490
rect 9757 -2930 9809 -2675
rect 9757 -3500 9809 -3490
rect 9875 -2930 9931 -2920
rect 9875 -3500 9931 -3490
rect 9993 -2930 10045 -2675
rect 9993 -3500 10045 -3490
rect 10111 -2930 10167 -2920
rect 10111 -3500 10167 -3490
rect 10229 -2930 10281 -2675
rect 10229 -3500 10281 -3490
rect 10347 -2930 10403 -2920
rect 10347 -3500 10403 -3490
rect 10465 -2930 10517 -2675
rect 10465 -3500 10517 -3490
rect 10583 -2930 10639 -2920
rect 10583 -3500 10639 -3490
rect 10701 -2930 10753 -2675
rect 10701 -3500 10753 -3490
rect 4136 -3544 4857 -3543
rect 4136 -3551 10697 -3544
rect 4136 -3705 4857 -3551
rect 4915 -3705 4975 -3551
rect 5033 -3705 5093 -3551
rect 5151 -3705 5211 -3551
rect 5269 -3705 5329 -3551
rect 5387 -3705 5447 -3551
rect 5505 -3705 5565 -3551
rect 5623 -3705 5683 -3551
rect 5741 -3705 5801 -3551
rect 5859 -3705 5919 -3551
rect 5977 -3705 6037 -3551
rect 6095 -3705 6155 -3551
rect 6213 -3705 6273 -3551
rect 6331 -3705 6391 -3551
rect 6449 -3705 6509 -3551
rect 6567 -3705 6627 -3551
rect 6685 -3705 6745 -3551
rect 6803 -3705 6863 -3551
rect 6921 -3705 6981 -3551
rect 7039 -3705 7099 -3551
rect 7157 -3705 7217 -3551
rect 7275 -3705 7335 -3551
rect 7393 -3705 7453 -3551
rect 7511 -3705 7571 -3551
rect 7629 -3705 7689 -3551
rect 7747 -3705 7807 -3551
rect 7865 -3705 7925 -3551
rect 7983 -3705 8043 -3551
rect 8101 -3705 8161 -3551
rect 8219 -3705 8279 -3551
rect 8337 -3705 8397 -3551
rect 8455 -3705 8515 -3551
rect 8573 -3705 8633 -3551
rect 8691 -3705 8751 -3551
rect 8809 -3705 8869 -3551
rect 8927 -3705 8987 -3551
rect 9045 -3705 9105 -3551
rect 9163 -3705 9223 -3551
rect 9281 -3705 9341 -3551
rect 9399 -3705 9459 -3551
rect 9517 -3705 9577 -3551
rect 9635 -3705 9695 -3551
rect 9753 -3705 9813 -3551
rect 9871 -3705 9931 -3551
rect 9989 -3705 10049 -3551
rect 10107 -3705 10167 -3551
rect 10225 -3705 10285 -3551
rect 10343 -3705 10403 -3551
rect 10461 -3705 10521 -3551
rect 10579 -3705 10639 -3551
rect 4136 -3711 10697 -3705
rect 4136 -4529 4304 -3711
rect 4801 -3766 4853 -3756
rect 4801 -4475 4853 -4326
rect 4919 -3766 4975 -3756
rect 4919 -4336 4975 -4326
rect 5037 -3766 5089 -3756
rect 5037 -4475 5089 -4326
rect 5155 -3766 5211 -3756
rect 5155 -4336 5211 -4326
rect 5273 -3766 5325 -3756
rect 5273 -4475 5325 -4326
rect 5391 -3766 5447 -3756
rect 5391 -4336 5447 -4326
rect 5509 -3766 5561 -3756
rect 5509 -4475 5561 -4326
rect 5627 -3766 5683 -3756
rect 5627 -4336 5683 -4326
rect 5745 -3766 5797 -3756
rect 5745 -4475 5797 -4326
rect 5863 -3766 5919 -3756
rect 5863 -4336 5919 -4326
rect 5981 -3766 6033 -3756
rect 5981 -4475 6033 -4326
rect 6099 -3766 6155 -3756
rect 6099 -4336 6155 -4326
rect 6217 -3766 6269 -3756
rect 6217 -4475 6269 -4326
rect 6335 -3766 6391 -3756
rect 6335 -4336 6391 -4326
rect 6453 -3766 6505 -3756
rect 6453 -4475 6505 -4326
rect 6571 -3766 6627 -3756
rect 6571 -4336 6627 -4326
rect 6689 -3766 6741 -3756
rect 6689 -4475 6741 -4326
rect 6807 -3766 6863 -3756
rect 6807 -4336 6863 -4326
rect 6925 -3766 6977 -3756
rect 6925 -4475 6977 -4326
rect 7043 -3766 7099 -3756
rect 7043 -4336 7099 -4326
rect 7161 -3766 7213 -3756
rect 7161 -4475 7213 -4326
rect 7279 -3766 7335 -3756
rect 7279 -4336 7335 -4326
rect 7397 -3766 7449 -3756
rect 7397 -4475 7449 -4326
rect 7515 -3766 7571 -3756
rect 7515 -4336 7571 -4326
rect 7633 -3766 7685 -3756
rect 7633 -4475 7685 -4326
rect 7751 -3766 7807 -3756
rect 7751 -4336 7807 -4326
rect 7869 -3766 7921 -3756
rect 7869 -4475 7921 -4326
rect 7987 -3766 8043 -3756
rect 7987 -4336 8043 -4326
rect 8105 -3766 8157 -3756
rect 8105 -4475 8157 -4326
rect 8223 -3766 8279 -3756
rect 8223 -4336 8279 -4326
rect 8341 -3766 8393 -3756
rect 8341 -4475 8393 -4326
rect 8459 -3766 8515 -3756
rect 8459 -4336 8515 -4326
rect 8577 -3766 8629 -3756
rect 8577 -4475 8629 -4326
rect 8695 -3766 8751 -3756
rect 8695 -4336 8751 -4326
rect 8813 -3766 8865 -3756
rect 8813 -4475 8865 -4326
rect 8931 -3766 8987 -3756
rect 8931 -4336 8987 -4326
rect 9049 -3766 9101 -3756
rect 9049 -4475 9101 -4326
rect 9167 -3766 9223 -3756
rect 9167 -4336 9223 -4326
rect 9285 -3766 9337 -3756
rect 9285 -4475 9337 -4326
rect 9403 -3766 9459 -3756
rect 9403 -4336 9459 -4326
rect 9521 -3766 9573 -3756
rect 9521 -4475 9573 -4326
rect 9639 -3766 9695 -3756
rect 9639 -4336 9695 -4326
rect 9757 -3766 9809 -3756
rect 9757 -4475 9809 -4326
rect 9875 -3766 9931 -3756
rect 9875 -4336 9931 -4326
rect 9993 -3766 10045 -3756
rect 9993 -4475 10045 -4326
rect 10111 -3766 10167 -3756
rect 10111 -4336 10167 -4326
rect 10229 -3766 10281 -3756
rect 10229 -4475 10281 -4326
rect 10347 -3766 10403 -3756
rect 10347 -4336 10403 -4326
rect 10465 -3766 10517 -3756
rect 10465 -4475 10517 -4326
rect 10583 -3766 10639 -3756
rect 10583 -4336 10639 -4326
rect 10701 -3766 10753 -3756
rect 10701 -4475 10753 -4326
rect 10841 -4475 11612 -2675
rect 3032 -4777 4304 -4529
rect 4760 -4725 4801 -4475
rect 4853 -4725 5037 -4475
rect 5089 -4725 5273 -4475
rect 5325 -4725 5509 -4475
rect 5561 -4725 5745 -4475
rect 5797 -4725 5981 -4475
rect 6033 -4725 6217 -4475
rect 6269 -4725 6453 -4475
rect 6505 -4725 6689 -4475
rect 6741 -4725 6925 -4475
rect 6977 -4725 7161 -4475
rect 7213 -4725 7397 -4475
rect 7449 -4725 7633 -4475
rect 7685 -4725 7869 -4475
rect 7921 -4725 8105 -4475
rect 8157 -4725 8341 -4475
rect 8393 -4725 8577 -4475
rect 8629 -4725 8813 -4475
rect 8865 -4725 9049 -4475
rect 9101 -4725 9285 -4475
rect 9337 -4725 9521 -4475
rect 9573 -4725 9757 -4475
rect 9809 -4725 9993 -4475
rect 10045 -4725 10229 -4475
rect 10281 -4725 10465 -4475
rect 10517 -4725 10701 -4475
rect 10753 -4725 11612 -4475
rect 4136 -5593 4304 -4777
rect 4801 -4980 4853 -4725
rect 4801 -5550 4853 -5540
rect 4919 -4980 4975 -4970
rect 4919 -5550 4975 -5540
rect 5037 -4980 5089 -4725
rect 5037 -5550 5089 -5540
rect 5155 -4980 5211 -4970
rect 5155 -5550 5211 -5540
rect 5273 -4980 5325 -4725
rect 5273 -5550 5325 -5540
rect 5391 -4980 5447 -4970
rect 5391 -5550 5447 -5540
rect 5509 -4980 5561 -4725
rect 5509 -5550 5561 -5540
rect 5627 -4980 5683 -4970
rect 5627 -5550 5683 -5540
rect 5745 -4980 5797 -4725
rect 5745 -5550 5797 -5540
rect 5863 -4980 5919 -4970
rect 5863 -5550 5919 -5540
rect 5981 -4980 6033 -4725
rect 5981 -5550 6033 -5540
rect 6099 -4980 6155 -4970
rect 6099 -5550 6155 -5540
rect 6217 -4980 6269 -4725
rect 6217 -5550 6269 -5540
rect 6335 -4980 6391 -4970
rect 6335 -5550 6391 -5540
rect 6453 -4980 6505 -4725
rect 6453 -5550 6505 -5540
rect 6571 -4980 6627 -4970
rect 6571 -5550 6627 -5540
rect 6689 -4980 6741 -4725
rect 6689 -5550 6741 -5540
rect 6807 -4980 6863 -4970
rect 6807 -5550 6863 -5540
rect 6925 -4980 6977 -4725
rect 6925 -5550 6977 -5540
rect 7043 -4980 7099 -4970
rect 7043 -5550 7099 -5540
rect 7161 -4980 7213 -4725
rect 7161 -5550 7213 -5540
rect 7279 -4980 7335 -4970
rect 7279 -5550 7335 -5540
rect 7397 -4980 7449 -4725
rect 7397 -5550 7449 -5540
rect 7515 -4980 7571 -4970
rect 7515 -5550 7571 -5540
rect 7633 -4980 7685 -4725
rect 7633 -5550 7685 -5540
rect 7751 -4980 7807 -4970
rect 7751 -5550 7807 -5540
rect 7869 -4980 7921 -4725
rect 7869 -5550 7921 -5540
rect 7987 -4980 8043 -4970
rect 7987 -5550 8043 -5540
rect 8105 -4980 8157 -4725
rect 8105 -5550 8157 -5540
rect 8223 -4980 8279 -4970
rect 8223 -5550 8279 -5540
rect 8341 -4980 8393 -4725
rect 8341 -5550 8393 -5540
rect 8459 -4980 8515 -4970
rect 8459 -5550 8515 -5540
rect 8577 -4980 8629 -4725
rect 8577 -5550 8629 -5540
rect 8695 -4980 8751 -4970
rect 8695 -5550 8751 -5540
rect 8813 -4980 8865 -4725
rect 8813 -5550 8865 -5540
rect 8931 -4980 8987 -4970
rect 8931 -5550 8987 -5540
rect 9049 -4980 9101 -4725
rect 9049 -5550 9101 -5540
rect 9167 -4980 9223 -4970
rect 9167 -5550 9223 -5540
rect 9285 -4980 9337 -4725
rect 9285 -5550 9337 -5540
rect 9403 -4980 9459 -4970
rect 9403 -5550 9459 -5540
rect 9521 -4980 9573 -4725
rect 9521 -5550 9573 -5540
rect 9639 -4980 9695 -4970
rect 9639 -5550 9695 -5540
rect 9757 -4980 9809 -4725
rect 9757 -5550 9809 -5540
rect 9875 -4980 9931 -4970
rect 9875 -5550 9931 -5540
rect 9993 -4980 10045 -4725
rect 9993 -5550 10045 -5540
rect 10111 -4980 10167 -4970
rect 10111 -5550 10167 -5540
rect 10229 -4980 10281 -4725
rect 10229 -5550 10281 -5540
rect 10347 -4980 10403 -4970
rect 10347 -5550 10403 -5540
rect 10465 -4980 10517 -4725
rect 10465 -5550 10517 -5540
rect 10583 -4980 10639 -4970
rect 10583 -5550 10639 -5540
rect 10701 -4980 10753 -4725
rect 10701 -5550 10753 -5540
rect 4136 -5594 5029 -5593
rect 4136 -5601 10697 -5594
rect 4136 -5755 4857 -5601
rect 4915 -5755 4975 -5601
rect 5033 -5755 5093 -5601
rect 5151 -5755 5211 -5601
rect 5269 -5755 5329 -5601
rect 5387 -5755 5447 -5601
rect 5505 -5755 5565 -5601
rect 5623 -5755 5683 -5601
rect 5741 -5755 5801 -5601
rect 5859 -5755 5919 -5601
rect 5977 -5755 6037 -5601
rect 6095 -5755 6155 -5601
rect 6213 -5755 6273 -5601
rect 6331 -5755 6391 -5601
rect 6449 -5755 6509 -5601
rect 6567 -5755 6627 -5601
rect 6685 -5755 6745 -5601
rect 6803 -5755 6863 -5601
rect 6921 -5755 6981 -5601
rect 7039 -5755 7099 -5601
rect 7157 -5755 7217 -5601
rect 7275 -5755 7335 -5601
rect 7393 -5755 7453 -5601
rect 7511 -5755 7571 -5601
rect 7629 -5755 7689 -5601
rect 7747 -5755 7807 -5601
rect 7865 -5755 7925 -5601
rect 7983 -5755 8043 -5601
rect 8101 -5755 8161 -5601
rect 8219 -5755 8279 -5601
rect 8337 -5755 8397 -5601
rect 8455 -5755 8515 -5601
rect 8573 -5755 8633 -5601
rect 8691 -5755 8751 -5601
rect 8809 -5755 8869 -5601
rect 8927 -5755 8987 -5601
rect 9045 -5755 9105 -5601
rect 9163 -5755 9223 -5601
rect 9281 -5755 9341 -5601
rect 9399 -5755 9459 -5601
rect 9517 -5755 9577 -5601
rect 9635 -5755 9695 -5601
rect 9753 -5755 9813 -5601
rect 9871 -5755 9931 -5601
rect 9989 -5755 10049 -5601
rect 10107 -5755 10167 -5601
rect 10225 -5755 10285 -5601
rect 10343 -5755 10403 -5601
rect 10461 -5755 10521 -5601
rect 10579 -5755 10639 -5601
rect 4136 -5761 10697 -5755
rect 4801 -5816 4853 -5806
rect 4801 -6525 4853 -6376
rect 4919 -5816 4975 -5806
rect 4919 -6386 4975 -6376
rect 5037 -5816 5089 -5806
rect 5037 -6525 5089 -6376
rect 5155 -5816 5211 -5806
rect 5155 -6386 5211 -6376
rect 5273 -5816 5325 -5806
rect 5273 -6525 5325 -6376
rect 5391 -5816 5447 -5806
rect 5391 -6386 5447 -6376
rect 5509 -5816 5561 -5806
rect 5509 -6525 5561 -6376
rect 5627 -5816 5683 -5806
rect 5627 -6386 5683 -6376
rect 5745 -5816 5797 -5806
rect 5745 -6525 5797 -6376
rect 5863 -5816 5919 -5806
rect 5863 -6386 5919 -6376
rect 5981 -5816 6033 -5806
rect 5981 -6525 6033 -6376
rect 6099 -5816 6155 -5806
rect 6099 -6386 6155 -6376
rect 6217 -5816 6269 -5806
rect 6217 -6525 6269 -6376
rect 6335 -5816 6391 -5806
rect 6335 -6386 6391 -6376
rect 6453 -5816 6505 -5806
rect 6453 -6525 6505 -6376
rect 6571 -5816 6627 -5806
rect 6571 -6386 6627 -6376
rect 6689 -5816 6741 -5806
rect 6689 -6525 6741 -6376
rect 6807 -5816 6863 -5806
rect 6807 -6386 6863 -6376
rect 6925 -5816 6977 -5806
rect 6925 -6525 6977 -6376
rect 7043 -5816 7099 -5806
rect 7043 -6386 7099 -6376
rect 7161 -5816 7213 -5806
rect 7161 -6525 7213 -6376
rect 7279 -5816 7335 -5806
rect 7279 -6386 7335 -6376
rect 7397 -5816 7449 -5806
rect 7397 -6525 7449 -6376
rect 7515 -5816 7571 -5806
rect 7515 -6386 7571 -6376
rect 7633 -5816 7685 -5806
rect 7633 -6525 7685 -6376
rect 7751 -5816 7807 -5806
rect 7751 -6386 7807 -6376
rect 7869 -5816 7921 -5806
rect 7869 -6525 7921 -6376
rect 7987 -5816 8043 -5806
rect 7987 -6386 8043 -6376
rect 8105 -5816 8157 -5806
rect 8105 -6525 8157 -6376
rect 8223 -5816 8279 -5806
rect 8223 -6386 8279 -6376
rect 8341 -5816 8393 -5806
rect 8341 -6525 8393 -6376
rect 8459 -5816 8515 -5806
rect 8459 -6386 8515 -6376
rect 8577 -5816 8629 -5806
rect 8577 -6525 8629 -6376
rect 8695 -5816 8751 -5806
rect 8695 -6386 8751 -6376
rect 8813 -5816 8865 -5806
rect 8813 -6525 8865 -6376
rect 8931 -5816 8987 -5806
rect 8931 -6386 8987 -6376
rect 9049 -5816 9101 -5806
rect 9049 -6525 9101 -6376
rect 9167 -5816 9223 -5806
rect 9167 -6386 9223 -6376
rect 9285 -5816 9337 -5806
rect 9285 -6525 9337 -6376
rect 9403 -5816 9459 -5806
rect 9403 -6386 9459 -6376
rect 9521 -5816 9573 -5806
rect 9521 -6525 9573 -6376
rect 9639 -5816 9695 -5806
rect 9639 -6386 9695 -6376
rect 9757 -5816 9809 -5806
rect 9757 -6525 9809 -6376
rect 9875 -5816 9931 -5806
rect 9875 -6386 9931 -6376
rect 9993 -5816 10045 -5806
rect 9993 -6525 10045 -6376
rect 10111 -5816 10167 -5806
rect 10111 -6386 10167 -6376
rect 10229 -5816 10281 -5806
rect 10229 -6525 10281 -6376
rect 10347 -5816 10403 -5806
rect 10347 -6386 10403 -6376
rect 10465 -5816 10517 -5806
rect 10465 -6525 10517 -6376
rect 10583 -5816 10639 -5806
rect 10583 -6386 10639 -6376
rect 10701 -5816 10753 -5806
rect 10701 -6525 10753 -6376
rect 10841 -6525 11612 -4725
rect 4760 -6775 4801 -6525
rect 4853 -6775 5037 -6525
rect 5089 -6775 5273 -6525
rect 5325 -6775 5509 -6525
rect 5561 -6775 5745 -6525
rect 5797 -6775 5981 -6525
rect 6033 -6775 6217 -6525
rect 6269 -6775 6453 -6525
rect 6505 -6775 6689 -6525
rect 6741 -6775 6925 -6525
rect 6977 -6775 7161 -6525
rect 7213 -6775 7397 -6525
rect 7449 -6775 7633 -6525
rect 7685 -6775 7869 -6525
rect 7921 -6775 8105 -6525
rect 8157 -6775 8341 -6525
rect 8393 -6775 8577 -6525
rect 8629 -6775 8813 -6525
rect 8865 -6775 9049 -6525
rect 9101 -6775 9285 -6525
rect 9337 -6775 9521 -6525
rect 9573 -6775 9757 -6525
rect 9809 -6775 9993 -6525
rect 10045 -6775 10229 -6525
rect 10281 -6775 10465 -6525
rect 10517 -6775 10701 -6525
rect 10753 -6625 11612 -6525
rect 10753 -6628 10903 -6625
rect 11463 -6628 11612 -6625
rect 10753 -6775 10902 -6628
rect 4760 -6776 10902 -6775
rect 11057 -6698 11617 -6690
rect 11057 -6754 11066 -6698
rect 11122 -6754 11147 -6698
rect 11203 -6754 11228 -6698
rect 11284 -6754 11309 -6698
rect 11365 -6754 11390 -6698
rect 11446 -6754 11471 -6698
rect 11527 -6754 11552 -6698
rect 11608 -6754 11617 -6698
rect 4801 -6785 4853 -6776
rect 5037 -6785 5089 -6776
rect 5273 -6785 5325 -6776
rect 5509 -6785 5561 -6776
rect 5745 -6785 5797 -6776
rect 5981 -6785 6033 -6776
rect 6217 -6785 6269 -6776
rect 6453 -6785 6505 -6776
rect 6689 -6785 6741 -6776
rect 6925 -6785 6977 -6776
rect 7161 -6785 7213 -6776
rect 7397 -6785 7449 -6776
rect 7633 -6785 7685 -6776
rect 7869 -6785 7921 -6776
rect 8105 -6785 8157 -6776
rect 8341 -6785 8393 -6776
rect 8577 -6785 8629 -6776
rect 8813 -6785 8865 -6776
rect 9049 -6785 9101 -6776
rect 9285 -6785 9337 -6776
rect 9521 -6785 9573 -6776
rect 9757 -6785 9809 -6776
rect 9993 -6785 10045 -6776
rect 10229 -6785 10281 -6776
rect 10465 -6785 10517 -6776
rect 10701 -6785 10753 -6776
rect 11057 -6802 11617 -6754
rect 11057 -6858 11066 -6802
rect 11122 -6858 11147 -6802
rect 11203 -6858 11228 -6802
rect 11284 -6858 11309 -6802
rect 11365 -6858 11390 -6802
rect 11446 -6858 11471 -6802
rect 11527 -6858 11552 -6802
rect 11608 -6858 11617 -6802
rect 11057 -6906 11617 -6858
rect 4083 -6942 10851 -6928
rect 4083 -6994 5759 -6942
rect 5811 -6994 5839 -6942
rect 5891 -6994 5919 -6942
rect 5971 -6994 5999 -6942
rect 6051 -6994 6079 -6942
rect 6131 -6994 6159 -6942
rect 6211 -6994 6239 -6942
rect 6291 -6994 6319 -6942
rect 6371 -6994 6399 -6942
rect 6451 -6994 6479 -6942
rect 6531 -6994 6559 -6942
rect 6611 -6994 6639 -6942
rect 6691 -6994 6719 -6942
rect 6771 -6994 6799 -6942
rect 6851 -6994 6879 -6942
rect 6931 -6994 6959 -6942
rect 7011 -6994 7039 -6942
rect 7091 -6994 7119 -6942
rect 7171 -6994 7199 -6942
rect 7251 -6994 7279 -6942
rect 7331 -6994 7359 -6942
rect 7411 -6994 7439 -6942
rect 7491 -6994 7519 -6942
rect 7571 -6994 7599 -6942
rect 7651 -6994 7679 -6942
rect 7731 -6994 7759 -6942
rect 7811 -6994 7839 -6942
rect 7891 -6994 7919 -6942
rect 7971 -6994 7999 -6942
rect 8051 -6994 8079 -6942
rect 8131 -6994 8159 -6942
rect 8211 -6994 8239 -6942
rect 8291 -6994 8319 -6942
rect 8371 -6994 8399 -6942
rect 8451 -6994 8479 -6942
rect 8531 -6994 8559 -6942
rect 8611 -6994 8639 -6942
rect 8691 -6994 8719 -6942
rect 8771 -6994 8799 -6942
rect 8851 -6994 8879 -6942
rect 8931 -6994 8959 -6942
rect 9011 -6994 9039 -6942
rect 9091 -6994 9119 -6942
rect 9171 -6994 9199 -6942
rect 9251 -6994 9279 -6942
rect 9331 -6994 9359 -6942
rect 9411 -6994 9439 -6942
rect 9491 -6994 9519 -6942
rect 9571 -6994 9599 -6942
rect 9651 -6994 9679 -6942
rect 9731 -6994 9759 -6942
rect 9811 -6994 9839 -6942
rect 9891 -6994 9919 -6942
rect 9971 -6994 9999 -6942
rect 10051 -6994 10079 -6942
rect 10131 -6994 10159 -6942
rect 10211 -6994 10239 -6942
rect 10291 -6994 10319 -6942
rect 10371 -6994 10399 -6942
rect 10451 -6994 10479 -6942
rect 10531 -6994 10559 -6942
rect 10611 -6994 10639 -6942
rect 10691 -6994 10719 -6942
rect 10771 -6994 10799 -6942
rect 11057 -6962 11066 -6906
rect 11122 -6962 11147 -6906
rect 11203 -6962 11228 -6906
rect 11284 -6962 11309 -6906
rect 11365 -6962 11390 -6906
rect 11446 -6962 11471 -6906
rect 11527 -6962 11552 -6906
rect 11608 -6962 11617 -6906
rect 11057 -6972 11617 -6962
rect 4083 -7022 10851 -6994
rect 4083 -7061 5759 -7022
rect 4083 -7117 4092 -7061
rect 4148 -7117 4173 -7061
rect 4229 -7117 4254 -7061
rect 4310 -7117 4335 -7061
rect 4391 -7117 4416 -7061
rect 4472 -7117 4497 -7061
rect 4553 -7117 4578 -7061
rect 4634 -7117 4660 -7061
rect 4716 -7117 4741 -7061
rect 4797 -7117 4822 -7061
rect 4878 -7117 4903 -7061
rect 4959 -7117 4984 -7061
rect 5040 -7117 5065 -7061
rect 5121 -7117 5146 -7061
rect 5202 -7117 5228 -7061
rect 5284 -7117 5309 -7061
rect 5365 -7117 5390 -7061
rect 5446 -7074 5759 -7061
rect 5811 -7074 5839 -7022
rect 5891 -7074 5919 -7022
rect 5971 -7074 5999 -7022
rect 6051 -7074 6079 -7022
rect 6131 -7074 6159 -7022
rect 6211 -7074 6239 -7022
rect 6291 -7074 6319 -7022
rect 6371 -7074 6399 -7022
rect 6451 -7074 6479 -7022
rect 6531 -7074 6559 -7022
rect 6611 -7074 6639 -7022
rect 6691 -7074 6719 -7022
rect 6771 -7074 6799 -7022
rect 6851 -7074 6879 -7022
rect 6931 -7074 6959 -7022
rect 7011 -7074 7039 -7022
rect 7091 -7074 7119 -7022
rect 7171 -7074 7199 -7022
rect 7251 -7074 7279 -7022
rect 7331 -7074 7359 -7022
rect 7411 -7074 7439 -7022
rect 7491 -7074 7519 -7022
rect 7571 -7074 7599 -7022
rect 7651 -7074 7679 -7022
rect 7731 -7074 7759 -7022
rect 7811 -7074 7839 -7022
rect 7891 -7074 7919 -7022
rect 7971 -7074 7999 -7022
rect 8051 -7074 8079 -7022
rect 8131 -7074 8159 -7022
rect 8211 -7074 8239 -7022
rect 8291 -7074 8319 -7022
rect 8371 -7074 8399 -7022
rect 8451 -7074 8479 -7022
rect 8531 -7074 8559 -7022
rect 8611 -7074 8639 -7022
rect 8691 -7074 8719 -7022
rect 8771 -7074 8799 -7022
rect 8851 -7074 8879 -7022
rect 8931 -7074 8959 -7022
rect 9011 -7074 9039 -7022
rect 9091 -7074 9119 -7022
rect 9171 -7074 9199 -7022
rect 9251 -7074 9279 -7022
rect 9331 -7074 9359 -7022
rect 9411 -7074 9439 -7022
rect 9491 -7074 9519 -7022
rect 9571 -7074 9599 -7022
rect 9651 -7074 9679 -7022
rect 9731 -7074 9759 -7022
rect 9811 -7074 9839 -7022
rect 9891 -7074 9919 -7022
rect 9971 -7074 9999 -7022
rect 10051 -7074 10079 -7022
rect 10131 -7074 10159 -7022
rect 10211 -7074 10239 -7022
rect 10291 -7074 10319 -7022
rect 10371 -7074 10399 -7022
rect 10451 -7074 10479 -7022
rect 10531 -7074 10559 -7022
rect 10611 -7074 10639 -7022
rect 10691 -7074 10719 -7022
rect 10771 -7074 10799 -7022
rect 5446 -7088 10851 -7074
rect 5446 -7100 5766 -7088
rect 5446 -7117 5471 -7100
rect 4083 -7165 5471 -7117
rect 4083 -7221 4092 -7165
rect 4148 -7221 4173 -7165
rect 4229 -7221 4254 -7165
rect 4310 -7221 4335 -7165
rect 4391 -7221 4416 -7165
rect 4472 -7221 4497 -7165
rect 4553 -7221 4578 -7165
rect 4634 -7221 4660 -7165
rect 4716 -7221 4741 -7165
rect 4797 -7221 4822 -7165
rect 4878 -7221 4903 -7165
rect 4959 -7221 4984 -7165
rect 5040 -7221 5065 -7165
rect 5121 -7221 5146 -7165
rect 5202 -7221 5228 -7165
rect 5284 -7221 5309 -7165
rect 5365 -7221 5390 -7165
rect 5446 -7221 5471 -7165
rect 4083 -7269 5471 -7221
rect 4083 -7325 4092 -7269
rect 4148 -7325 4173 -7269
rect 4229 -7325 4254 -7269
rect 4310 -7325 4335 -7269
rect 4391 -7325 4416 -7269
rect 4472 -7325 4497 -7269
rect 4553 -7325 4578 -7269
rect 4634 -7325 4660 -7269
rect 4716 -7325 4741 -7269
rect 4797 -7325 4822 -7269
rect 4878 -7325 4903 -7269
rect 4959 -7325 4984 -7269
rect 5040 -7325 5065 -7269
rect 5121 -7325 5146 -7269
rect 5202 -7325 5228 -7269
rect 5284 -7325 5309 -7269
rect 5365 -7325 5390 -7269
rect 5446 -7325 5471 -7269
rect 4083 -7373 5471 -7325
rect 4083 -7429 4092 -7373
rect 4148 -7429 4173 -7373
rect 4229 -7429 4254 -7373
rect 4310 -7429 4335 -7373
rect 4391 -7429 4416 -7373
rect 4472 -7429 4497 -7373
rect 4553 -7429 4578 -7373
rect 4634 -7429 4660 -7373
rect 4716 -7429 4741 -7373
rect 4797 -7429 4822 -7373
rect 4878 -7429 4903 -7373
rect 4959 -7429 4984 -7373
rect 5040 -7429 5065 -7373
rect 5121 -7429 5146 -7373
rect 5202 -7429 5228 -7373
rect 5284 -7429 5309 -7373
rect 5365 -7429 5390 -7373
rect 5446 -7429 5471 -7373
rect 4083 -7477 5471 -7429
rect 4083 -7533 4092 -7477
rect 4148 -7533 4173 -7477
rect 4229 -7533 4254 -7477
rect 4310 -7533 4335 -7477
rect 4391 -7533 4416 -7477
rect 4472 -7533 4497 -7477
rect 4553 -7533 4578 -7477
rect 4634 -7533 4660 -7477
rect 4716 -7533 4741 -7477
rect 4797 -7533 4822 -7477
rect 4878 -7533 4903 -7477
rect 4959 -7533 4984 -7477
rect 5040 -7533 5065 -7477
rect 5121 -7533 5146 -7477
rect 5202 -7533 5228 -7477
rect 5284 -7533 5309 -7477
rect 5365 -7533 5390 -7477
rect 5446 -7533 5471 -7477
rect 4083 -7581 5471 -7533
rect 4083 -7637 4092 -7581
rect 4148 -7637 4173 -7581
rect 4229 -7637 4254 -7581
rect 4310 -7637 4335 -7581
rect 4391 -7637 4416 -7581
rect 4472 -7637 4497 -7581
rect 4553 -7637 4578 -7581
rect 4634 -7637 4660 -7581
rect 4716 -7637 4741 -7581
rect 4797 -7637 4822 -7581
rect 4878 -7637 4903 -7581
rect 4959 -7637 4984 -7581
rect 5040 -7637 5065 -7581
rect 5121 -7637 5146 -7581
rect 5202 -7637 5228 -7581
rect 5284 -7637 5309 -7581
rect 5365 -7637 5390 -7581
rect 5446 -7637 5471 -7581
rect 4083 -7685 5471 -7637
rect 4083 -7741 4092 -7685
rect 4148 -7741 4173 -7685
rect 4229 -7741 4254 -7685
rect 4310 -7741 4335 -7685
rect 4391 -7741 4416 -7685
rect 4472 -7741 4497 -7685
rect 4553 -7741 4578 -7685
rect 4634 -7741 4660 -7685
rect 4716 -7741 4741 -7685
rect 4797 -7741 4822 -7685
rect 4878 -7741 4903 -7685
rect 4959 -7741 4984 -7685
rect 5040 -7741 5065 -7685
rect 5121 -7741 5146 -7685
rect 5202 -7741 5228 -7685
rect 5284 -7741 5309 -7685
rect 5365 -7741 5390 -7685
rect 5446 -7741 5471 -7685
rect 4083 -7789 5471 -7741
rect 4083 -7845 4092 -7789
rect 4148 -7845 4173 -7789
rect 4229 -7845 4254 -7789
rect 4310 -7845 4335 -7789
rect 4391 -7845 4416 -7789
rect 4472 -7845 4497 -7789
rect 4553 -7845 4578 -7789
rect 4634 -7845 4660 -7789
rect 4716 -7845 4741 -7789
rect 4797 -7845 4822 -7789
rect 4878 -7845 4903 -7789
rect 4959 -7845 4984 -7789
rect 5040 -7845 5065 -7789
rect 5121 -7845 5146 -7789
rect 5202 -7845 5228 -7789
rect 5284 -7845 5309 -7789
rect 5365 -7845 5390 -7789
rect 5446 -7845 5471 -7789
rect 5867 -7223 5919 -7088
rect 5867 -7793 5919 -7783
rect 5983 -7223 6039 -7213
rect 5983 -7825 6039 -7783
rect 6103 -7223 6155 -7088
rect 6103 -7793 6155 -7783
rect 6219 -7223 6275 -7213
rect 6219 -7825 6275 -7783
rect 6339 -7223 6391 -7088
rect 6339 -7793 6391 -7783
rect 6455 -7223 6511 -7213
rect 6455 -7825 6511 -7783
rect 6575 -7223 6627 -7088
rect 6575 -7793 6627 -7783
rect 6691 -7223 6747 -7213
rect 6691 -7825 6747 -7783
rect 6811 -7223 6863 -7088
rect 6811 -7793 6863 -7783
rect 6927 -7223 6983 -7213
rect 6927 -7825 6983 -7783
rect 7047 -7223 7099 -7088
rect 7047 -7793 7099 -7783
rect 7163 -7223 7219 -7213
rect 7163 -7825 7219 -7783
rect 7283 -7223 7335 -7088
rect 7283 -7793 7335 -7783
rect 7399 -7223 7455 -7213
rect 7399 -7825 7455 -7783
rect 7519 -7223 7571 -7088
rect 7519 -7793 7571 -7783
rect 7635 -7223 7691 -7213
rect 7635 -7825 7691 -7783
rect 7865 -7223 7917 -7088
rect 7865 -7793 7917 -7783
rect 7981 -7223 8037 -7213
rect 7981 -7793 8037 -7783
rect 8101 -7223 8153 -7088
rect 8101 -7793 8153 -7783
rect 8217 -7223 8273 -7213
rect 8217 -7793 8273 -7783
rect 8337 -7223 8389 -7088
rect 8337 -7793 8389 -7783
rect 8453 -7223 8509 -7213
rect 8453 -7793 8509 -7783
rect 8573 -7223 8625 -7088
rect 8573 -7793 8625 -7783
rect 8689 -7223 8745 -7213
rect 8689 -7793 8745 -7783
rect 8809 -7223 8861 -7088
rect 8809 -7793 8861 -7783
rect 8925 -7223 8981 -7213
rect 8925 -7793 8981 -7783
rect 9045 -7223 9097 -7088
rect 9045 -7793 9097 -7783
rect 9161 -7223 9217 -7213
rect 9161 -7793 9217 -7783
rect 9281 -7223 9333 -7088
rect 9281 -7793 9333 -7783
rect 9397 -7223 9453 -7213
rect 9397 -7793 9453 -7783
rect 9517 -7223 9569 -7088
rect 9828 -7206 10401 -7088
rect 9517 -7793 9569 -7783
rect 9633 -7223 9689 -7213
rect 9828 -7258 9839 -7206
rect 9891 -7258 9919 -7206
rect 9971 -7258 9999 -7206
rect 10051 -7258 10079 -7206
rect 10131 -7258 10159 -7206
rect 10211 -7258 10239 -7206
rect 10291 -7258 10319 -7206
rect 10371 -7258 10401 -7206
rect 9828 -7285 10401 -7258
rect 11173 -7261 11602 -6972
rect 12523 -7219 12579 -7209
rect 9828 -7337 9839 -7285
rect 9891 -7337 9919 -7285
rect 9971 -7337 9999 -7285
rect 10051 -7337 10079 -7285
rect 10131 -7337 10159 -7285
rect 10211 -7337 10239 -7285
rect 10291 -7337 10319 -7285
rect 10371 -7337 10401 -7285
rect 10616 -7333 12209 -7261
rect 11173 -7335 11283 -7333
rect 9828 -7354 10401 -7337
rect 9828 -7406 9839 -7354
rect 9891 -7406 9919 -7354
rect 9971 -7406 9999 -7354
rect 10051 -7406 10079 -7354
rect 10131 -7406 10159 -7354
rect 10211 -7406 10239 -7354
rect 10291 -7406 10319 -7354
rect 10371 -7406 10401 -7354
rect 9828 -7433 10401 -7406
rect 9828 -7485 9839 -7433
rect 9891 -7485 9919 -7433
rect 9971 -7485 9999 -7433
rect 10051 -7485 10079 -7433
rect 10131 -7485 10159 -7433
rect 10211 -7485 10239 -7433
rect 10291 -7485 10319 -7433
rect 10371 -7485 10401 -7433
rect 9828 -7581 10401 -7485
rect 10513 -7395 10565 -7385
rect 9633 -7793 9689 -7783
rect 4083 -7893 5471 -7845
rect 4083 -7949 4092 -7893
rect 4148 -7949 4173 -7893
rect 4229 -7949 4254 -7893
rect 4310 -7949 4335 -7893
rect 4391 -7949 4416 -7893
rect 4472 -7949 4497 -7893
rect 4553 -7949 4578 -7893
rect 4634 -7949 4660 -7893
rect 4716 -7949 4741 -7893
rect 4797 -7949 4822 -7893
rect 4878 -7949 4903 -7893
rect 4959 -7949 4984 -7893
rect 5040 -7949 5065 -7893
rect 5121 -7949 5146 -7893
rect 5202 -7949 5228 -7893
rect 5284 -7949 5309 -7893
rect 5365 -7949 5390 -7893
rect 5446 -7949 5471 -7893
rect 4083 -7997 5471 -7949
rect 4083 -8053 4092 -7997
rect 4148 -8053 4173 -7997
rect 4229 -8053 4254 -7997
rect 4310 -8053 4335 -7997
rect 4391 -8053 4416 -7997
rect 4472 -8053 4497 -7997
rect 4553 -8053 4578 -7997
rect 4634 -8053 4660 -7997
rect 4716 -8053 4741 -7997
rect 4797 -8053 4822 -7997
rect 4878 -8053 4903 -7997
rect 4959 -8053 4984 -7997
rect 5040 -8053 5065 -7997
rect 5121 -8053 5146 -7997
rect 5202 -8053 5228 -7997
rect 5284 -8053 5309 -7997
rect 5365 -8053 5390 -7997
rect 5446 -8053 5471 -7997
rect 5923 -7835 9689 -7825
rect 5981 -7989 6041 -7835
rect 6099 -7989 6159 -7835
rect 6217 -7989 6277 -7835
rect 6335 -7989 6395 -7835
rect 6453 -7989 6513 -7835
rect 6571 -7989 6631 -7835
rect 6689 -7989 6749 -7835
rect 6807 -7989 6867 -7835
rect 6925 -7989 6985 -7835
rect 7043 -7989 7103 -7835
rect 7161 -7989 7221 -7835
rect 7279 -7989 7339 -7835
rect 7397 -7989 7457 -7835
rect 7515 -7989 7575 -7835
rect 7633 -7989 7921 -7835
rect 7979 -7989 8039 -7835
rect 8097 -7989 8157 -7835
rect 8215 -7989 8275 -7835
rect 8333 -7989 8393 -7835
rect 8451 -7989 8511 -7835
rect 8569 -7989 8629 -7835
rect 8687 -7989 8747 -7835
rect 8805 -7989 8865 -7835
rect 8923 -7989 8983 -7835
rect 9041 -7989 9101 -7835
rect 9159 -7989 9219 -7835
rect 9277 -7989 9337 -7835
rect 9395 -7989 9455 -7835
rect 9513 -7989 9573 -7835
rect 9631 -7989 9689 -7835
rect 5923 -7999 9689 -7989
rect 4083 -8101 5471 -8053
rect 4083 -8157 4092 -8101
rect 4148 -8157 4173 -8101
rect 4229 -8157 4254 -8101
rect 4310 -8157 4335 -8101
rect 4391 -8157 4416 -8101
rect 4472 -8157 4497 -8101
rect 4553 -8157 4578 -8101
rect 4634 -8157 4660 -8101
rect 4716 -8157 4741 -8101
rect 4797 -8157 4822 -8101
rect 4878 -8157 4903 -8101
rect 4959 -8157 4984 -8101
rect 5040 -8157 5065 -8101
rect 5121 -8157 5146 -8101
rect 5202 -8157 5228 -8101
rect 5284 -8157 5309 -8101
rect 5365 -8157 5390 -8101
rect 5446 -8157 5471 -8101
rect 4083 -8205 5471 -8157
rect 4083 -8261 4092 -8205
rect 4148 -8261 4173 -8205
rect 4229 -8261 4254 -8205
rect 4310 -8261 4335 -8205
rect 4391 -8261 4416 -8205
rect 4472 -8261 4497 -8205
rect 4553 -8261 4578 -8205
rect 4634 -8261 4660 -8205
rect 4716 -8261 4741 -8205
rect 4797 -8261 4822 -8205
rect 4878 -8261 4903 -8205
rect 4959 -8261 4984 -8205
rect 5040 -8261 5065 -8205
rect 5121 -8261 5146 -8205
rect 5202 -8261 5228 -8205
rect 5284 -8261 5309 -8205
rect 5365 -8261 5390 -8205
rect 5446 -8261 5471 -8205
rect 4083 -8309 5471 -8261
rect 4083 -8365 4092 -8309
rect 4148 -8365 4173 -8309
rect 4229 -8365 4254 -8309
rect 4310 -8365 4335 -8309
rect 4391 -8365 4416 -8309
rect 4472 -8365 4497 -8309
rect 4553 -8365 4578 -8309
rect 4634 -8365 4660 -8309
rect 4716 -8365 4741 -8309
rect 4797 -8365 4822 -8309
rect 4878 -8365 4903 -8309
rect 4959 -8365 4984 -8309
rect 5040 -8365 5065 -8309
rect 5121 -8365 5146 -8309
rect 5202 -8365 5228 -8309
rect 5284 -8365 5309 -8309
rect 5365 -8365 5390 -8309
rect 5446 -8365 5471 -8309
rect 4083 -8413 5471 -8365
rect 4083 -8469 4092 -8413
rect 4148 -8469 4173 -8413
rect 4229 -8469 4254 -8413
rect 4310 -8469 4335 -8413
rect 4391 -8469 4416 -8413
rect 4472 -8469 4497 -8413
rect 4553 -8469 4578 -8413
rect 4634 -8469 4660 -8413
rect 4716 -8469 4741 -8413
rect 4797 -8469 4822 -8413
rect 4878 -8469 4903 -8413
rect 4959 -8469 4984 -8413
rect 5040 -8469 5065 -8413
rect 5121 -8469 5146 -8413
rect 5202 -8469 5228 -8413
rect 5284 -8469 5309 -8413
rect 5365 -8469 5390 -8413
rect 5446 -8469 5471 -8413
rect 4083 -8517 5471 -8469
rect 4083 -8573 4092 -8517
rect 4148 -8573 4173 -8517
rect 4229 -8573 4254 -8517
rect 4310 -8573 4335 -8517
rect 4391 -8573 4416 -8517
rect 4472 -8573 4497 -8517
rect 4553 -8573 4578 -8517
rect 4634 -8573 4660 -8517
rect 4716 -8573 4741 -8517
rect 4797 -8573 4822 -8517
rect 4878 -8573 4903 -8517
rect 4959 -8573 4984 -8517
rect 5040 -8573 5065 -8517
rect 5121 -8573 5146 -8517
rect 5202 -8573 5228 -8517
rect 5284 -8573 5309 -8517
rect 5365 -8573 5390 -8517
rect 5446 -8573 5471 -8517
rect 4083 -8606 5471 -8573
rect 5867 -8041 5919 -8031
rect 5867 -8815 5919 -8601
rect 5983 -8041 6039 -7999
rect 5983 -8611 6039 -8601
rect 6103 -8041 6155 -8031
rect 6103 -8815 6155 -8601
rect 6219 -8041 6275 -7999
rect 6219 -8611 6275 -8601
rect 6339 -8041 6391 -8031
rect 6339 -8815 6391 -8601
rect 6455 -8041 6511 -7999
rect 6455 -8611 6511 -8601
rect 6575 -8041 6627 -8031
rect 6575 -8815 6627 -8601
rect 6691 -8041 6747 -7999
rect 6691 -8611 6747 -8601
rect 6811 -8041 6863 -8031
rect 6811 -8815 6863 -8601
rect 6927 -8041 6983 -7999
rect 6927 -8611 6983 -8601
rect 7047 -8041 7099 -8031
rect 7047 -8815 7099 -8601
rect 7163 -8041 7219 -7999
rect 7163 -8611 7219 -8601
rect 7283 -8041 7335 -8031
rect 7283 -8815 7335 -8601
rect 7399 -8041 7455 -7999
rect 7399 -8611 7455 -8601
rect 7519 -8041 7571 -8031
rect 7519 -8815 7571 -8601
rect 7635 -8041 7691 -7999
rect 10513 -8031 10565 -7515
rect 10625 -7395 10681 -7385
rect 10625 -7525 10681 -7515
rect 10829 -7395 10881 -7385
rect 10829 -8012 10881 -7515
rect 10941 -7395 10997 -7385
rect 10941 -7525 10997 -7515
rect 11145 -7395 11197 -7385
rect 11145 -8012 11197 -7515
rect 11257 -7395 11313 -7385
rect 11257 -7525 11313 -7515
rect 11461 -7395 11513 -7385
rect 11461 -8012 11513 -7515
rect 11573 -7395 11629 -7385
rect 11573 -7525 11629 -7515
rect 11777 -7395 11829 -7385
rect 11777 -8012 11829 -7515
rect 11889 -7395 11945 -7385
rect 11889 -7525 11945 -7515
rect 12093 -7395 12145 -7385
rect 10829 -8020 11914 -8012
rect 10825 -8031 10834 -8020
rect 7635 -8611 7691 -8601
rect 7865 -8041 7917 -8031
rect 7865 -8815 7917 -8601
rect 7981 -8041 8037 -8031
rect 7981 -8611 8037 -8601
rect 8101 -8041 8153 -8031
rect 8101 -8815 8153 -8601
rect 8217 -8041 8273 -8031
rect 8217 -8611 8273 -8601
rect 8337 -8041 8389 -8031
rect 8337 -8815 8389 -8601
rect 8453 -8041 8509 -8031
rect 8453 -8611 8509 -8601
rect 8573 -8041 8625 -8031
rect 8573 -8815 8625 -8601
rect 8689 -8041 8745 -8031
rect 8689 -8611 8745 -8601
rect 8809 -8041 8861 -8031
rect 8809 -8815 8861 -8601
rect 8925 -8041 8981 -8031
rect 8925 -8611 8981 -8601
rect 9045 -8041 9097 -8031
rect 9045 -8815 9097 -8601
rect 9161 -8041 9217 -8031
rect 9161 -8611 9217 -8601
rect 9281 -8041 9333 -8031
rect 9281 -8815 9333 -8601
rect 9397 -8041 9453 -8031
rect 9397 -8611 9453 -8601
rect 9517 -8041 9569 -8031
rect 9517 -8815 9569 -8601
rect 9633 -8041 9689 -8031
rect 10513 -8076 10834 -8031
rect 10890 -8076 10915 -8020
rect 10971 -8076 10996 -8020
rect 11052 -8076 11077 -8020
rect 11133 -8076 11158 -8020
rect 11214 -8076 11239 -8020
rect 11295 -8076 11320 -8020
rect 11376 -8076 11401 -8020
rect 11457 -8076 11482 -8020
rect 11538 -8076 11563 -8020
rect 11619 -8076 11644 -8020
rect 11700 -8076 11725 -8020
rect 11781 -8076 11806 -8020
rect 11862 -8076 11914 -8020
rect 10513 -8083 11914 -8076
rect 10825 -8124 11914 -8083
rect 10825 -8180 10834 -8124
rect 10890 -8180 10915 -8124
rect 10971 -8180 10996 -8124
rect 11052 -8180 11077 -8124
rect 11133 -8180 11158 -8124
rect 11214 -8180 11239 -8124
rect 11295 -8180 11320 -8124
rect 11376 -8180 11401 -8124
rect 11457 -8180 11482 -8124
rect 11538 -8180 11563 -8124
rect 11619 -8180 11644 -8124
rect 11700 -8180 11725 -8124
rect 11781 -8180 11806 -8124
rect 11862 -8126 11914 -8124
rect 12093 -8126 12145 -7515
rect 12205 -7395 12261 -7385
rect 12205 -7525 12261 -7515
rect 12523 -8069 12579 -8059
rect 12671 -7219 12727 -7209
rect 12671 -8069 12727 -8059
rect 12819 -7219 12875 -7209
rect 12819 -8069 12875 -8059
rect 12967 -7219 13023 -7209
rect 12967 -8069 13023 -8059
rect 13115 -7219 13171 -7209
rect 13115 -8069 13171 -8059
rect 13263 -7219 13319 -7209
rect 13263 -8069 13319 -8059
rect 13411 -7219 13467 -7209
rect 13411 -8069 13467 -8059
rect 13559 -7219 13615 -7209
rect 13559 -8069 13615 -8059
rect 13707 -7219 13763 -7209
rect 13707 -8069 13763 -8059
rect 13855 -7219 13911 -7209
rect 13855 -8069 13911 -8059
rect 14003 -7219 14059 -7209
rect 14003 -8069 14059 -8059
rect 14151 -7219 14207 -7209
rect 14151 -8069 14207 -8059
rect 14299 -7219 14355 -7209
rect 14299 -8069 14355 -8059
rect 14447 -7219 14503 -7209
rect 14447 -8069 14503 -8059
rect 14595 -7219 14651 -7209
rect 14595 -8069 14651 -8059
rect 14743 -7219 14799 -7209
rect 14743 -8069 14799 -8059
rect 14891 -7219 14947 -7209
rect 14891 -8069 14947 -8059
rect 15039 -7219 15095 -7209
rect 15039 -8069 15095 -8059
rect 15187 -7219 15243 -7209
rect 15187 -8069 15243 -8059
rect 15335 -7219 15391 -7209
rect 15335 -8069 15391 -8059
rect 15483 -7219 15539 -7209
rect 15483 -8069 15539 -8059
rect 15631 -7219 15687 -7209
rect 15631 -8069 15687 -8059
rect 15779 -7219 15835 -7209
rect 15779 -8069 15835 -8059
rect 15927 -7219 15983 -7209
rect 15927 -8069 15983 -8059
rect 16075 -7219 16131 -7209
rect 16075 -8069 16131 -8059
rect 16223 -7219 16279 -7209
rect 16223 -8069 16279 -8059
rect 16371 -7219 16427 -7209
rect 16371 -8069 16427 -8059
rect 16519 -7219 16575 -7209
rect 16519 -8069 16575 -8059
rect 16667 -7219 16723 -7209
rect 16667 -8069 16723 -8059
rect 16815 -7219 16871 -7209
rect 16815 -8069 16871 -8059
rect 16963 -7219 17019 -7209
rect 16963 -8069 17019 -8059
rect 17111 -7219 17167 -7209
rect 17111 -8069 17167 -8059
rect 17259 -7219 17315 -7209
rect 17259 -8069 17315 -8059
rect 17407 -7219 17463 -7209
rect 17407 -8069 17463 -8059
rect 17555 -7219 17611 -7209
rect 17555 -8069 17611 -8059
rect 17703 -7219 17759 -7209
rect 17703 -8069 17759 -8059
rect 17851 -7219 17907 -7209
rect 17851 -8069 17907 -8059
rect 17999 -7219 18055 -7209
rect 17999 -8069 18055 -8059
rect 18147 -7219 18203 -7209
rect 18147 -8069 18203 -8059
rect 18295 -7219 18351 -7209
rect 18295 -8069 18351 -8059
rect 18443 -7219 18499 -7209
rect 18443 -8069 18499 -8059
rect 18591 -7219 18647 -7209
rect 18591 -8069 18647 -8059
rect 18739 -7219 18795 -7209
rect 18739 -8069 18795 -8059
rect 18887 -7219 18943 -7209
rect 18887 -8069 18943 -8059
rect 19035 -7219 19091 -7209
rect 19035 -8069 19091 -8059
rect 19183 -7219 19239 -7209
rect 19183 -8069 19239 -8059
rect 19331 -7219 19387 -7209
rect 19331 -8069 19387 -8059
rect 19479 -7219 19535 -7209
rect 19479 -8069 19535 -8059
rect 19627 -7219 19683 -7209
rect 19627 -8069 19683 -8059
rect 19775 -7219 19831 -7209
rect 19775 -8069 19831 -8059
rect 19923 -7219 19979 -7209
rect 19923 -8069 19979 -8059
rect 20071 -7219 20127 -7209
rect 20071 -8069 20127 -8059
rect 20219 -7219 20275 -7209
rect 20219 -8069 20275 -8059
rect 20367 -7219 20423 -7209
rect 20367 -8069 20423 -8059
rect 20515 -7219 20571 -7209
rect 20515 -8069 20571 -8059
rect 20663 -7219 20719 -7209
rect 20663 -8069 20719 -8059
rect 20811 -7219 20867 -7209
rect 20811 -8069 20867 -8059
rect 20959 -7219 21015 -7209
rect 20959 -8069 21015 -8059
rect 21107 -7219 21163 -7209
rect 21107 -8069 21163 -8059
rect 21255 -7219 21311 -7209
rect 21255 -8069 21311 -8059
rect 21403 -7219 21459 -7209
rect 21403 -8069 21459 -8059
rect 21551 -7219 21607 -7209
rect 21551 -8069 21607 -8059
rect 21699 -7219 21755 -7209
rect 21699 -8069 21755 -8059
rect 21847 -7219 21903 -7209
rect 21847 -8069 21903 -8059
rect 21995 -7219 22051 -7209
rect 21995 -8069 22051 -8059
rect 22143 -7219 22199 -7209
rect 22143 -8069 22199 -8059
rect 22291 -7219 22347 -7209
rect 22291 -8069 22347 -8059
rect 22439 -7219 22495 -7209
rect 22439 -8069 22495 -8059
rect 22587 -7219 22643 -7209
rect 22587 -8069 22643 -8059
rect 22735 -7219 22791 -7209
rect 22735 -8069 22791 -8059
rect 22883 -7219 22939 -7209
rect 22883 -8069 22939 -8059
rect 23031 -7219 23087 -7209
rect 23031 -8069 23087 -8059
rect 23179 -7219 23235 -7209
rect 23179 -8069 23235 -8059
rect 23327 -7219 23383 -7209
rect 23327 -8069 23383 -8059
rect 23475 -7219 23531 -7209
rect 23475 -8069 23531 -8059
rect 23623 -7219 23679 -7209
rect 23623 -8069 23679 -8059
rect 12580 -8126 23632 -8125
rect 11862 -8135 23632 -8126
rect 11862 -8180 12580 -8135
rect 10825 -8228 12580 -8180
rect 10825 -8284 10834 -8228
rect 10890 -8284 10915 -8228
rect 10971 -8284 10996 -8228
rect 11052 -8284 11077 -8228
rect 11133 -8284 11158 -8228
rect 11214 -8284 11239 -8228
rect 11295 -8284 11320 -8228
rect 11376 -8284 11401 -8228
rect 11457 -8284 11482 -8228
rect 11538 -8284 11563 -8228
rect 11619 -8284 11644 -8228
rect 11700 -8284 11725 -8228
rect 11781 -8284 11806 -8228
rect 11862 -8284 12580 -8228
rect 10825 -8289 12580 -8284
rect 12670 -8289 12728 -8135
rect 12818 -8289 12876 -8135
rect 12966 -8289 13024 -8135
rect 13114 -8289 13172 -8135
rect 13262 -8289 13320 -8135
rect 13410 -8289 13468 -8135
rect 13558 -8289 13616 -8135
rect 13706 -8289 13764 -8135
rect 13854 -8289 13912 -8135
rect 14002 -8289 14060 -8135
rect 14150 -8289 14208 -8135
rect 14298 -8289 14356 -8135
rect 14446 -8289 14504 -8135
rect 14594 -8289 14652 -8135
rect 14742 -8289 14800 -8135
rect 14890 -8289 14948 -8135
rect 15038 -8289 15096 -8135
rect 15186 -8289 15244 -8135
rect 15334 -8289 15392 -8135
rect 15482 -8289 15540 -8135
rect 15630 -8289 15688 -8135
rect 15778 -8289 15836 -8135
rect 15926 -8289 15984 -8135
rect 16074 -8289 16132 -8135
rect 16222 -8289 16280 -8135
rect 16370 -8289 16428 -8135
rect 16518 -8289 16576 -8135
rect 16666 -8289 16724 -8135
rect 16814 -8289 16872 -8135
rect 16962 -8289 17020 -8135
rect 17110 -8289 17168 -8135
rect 17258 -8289 17316 -8135
rect 17406 -8289 17464 -8135
rect 17554 -8289 17612 -8135
rect 17702 -8289 17760 -8135
rect 17850 -8289 17908 -8135
rect 17998 -8289 18056 -8135
rect 18146 -8289 18204 -8135
rect 18294 -8289 18352 -8135
rect 18442 -8289 18500 -8135
rect 18590 -8289 18648 -8135
rect 18738 -8289 18796 -8135
rect 18886 -8289 18944 -8135
rect 19034 -8289 19092 -8135
rect 19182 -8289 19240 -8135
rect 19330 -8289 19388 -8135
rect 19478 -8289 19536 -8135
rect 19626 -8289 19684 -8135
rect 19774 -8289 19832 -8135
rect 19922 -8289 19980 -8135
rect 20070 -8289 20128 -8135
rect 20218 -8289 20276 -8135
rect 20366 -8289 20424 -8135
rect 20514 -8289 20572 -8135
rect 20662 -8289 20720 -8135
rect 20810 -8289 20868 -8135
rect 20958 -8289 21016 -8135
rect 21106 -8289 21164 -8135
rect 21254 -8289 21312 -8135
rect 21402 -8289 21460 -8135
rect 21550 -8289 21608 -8135
rect 21698 -8289 21756 -8135
rect 21846 -8289 21904 -8135
rect 21994 -8289 22052 -8135
rect 22142 -8289 22200 -8135
rect 22290 -8289 22348 -8135
rect 22438 -8289 22496 -8135
rect 22586 -8289 22644 -8135
rect 22734 -8289 22792 -8135
rect 22882 -8289 22940 -8135
rect 23030 -8289 23088 -8135
rect 23178 -8289 23236 -8135
rect 23326 -8289 23384 -8135
rect 23474 -8289 23532 -8135
rect 23622 -8289 23632 -8135
rect 10825 -8299 23632 -8289
rect 10825 -8332 11914 -8299
rect 10825 -8388 10834 -8332
rect 10890 -8388 10915 -8332
rect 10971 -8388 10996 -8332
rect 11052 -8388 11077 -8332
rect 11133 -8388 11158 -8332
rect 11214 -8388 11239 -8332
rect 11295 -8388 11320 -8332
rect 11376 -8388 11401 -8332
rect 11457 -8388 11482 -8332
rect 11538 -8388 11563 -8332
rect 11619 -8388 11644 -8332
rect 11700 -8388 11725 -8332
rect 11781 -8388 11806 -8332
rect 11862 -8388 11914 -8332
rect 10825 -8403 11914 -8388
rect 12523 -8365 12579 -8355
rect 9633 -8611 9689 -8601
rect 9828 -8538 10620 -8524
rect 9828 -8590 9839 -8538
rect 9891 -8590 9919 -8538
rect 9971 -8590 9999 -8538
rect 10051 -8590 10079 -8538
rect 10131 -8590 10159 -8538
rect 10211 -8590 10239 -8538
rect 10291 -8590 10319 -8538
rect 10371 -8590 10399 -8538
rect 10451 -8590 10479 -8538
rect 10531 -8590 10559 -8538
rect 10611 -8590 10620 -8538
rect 9828 -8617 10620 -8590
rect 9828 -8669 9839 -8617
rect 9891 -8669 9919 -8617
rect 9971 -8669 9999 -8617
rect 10051 -8669 10079 -8617
rect 10131 -8669 10159 -8617
rect 10211 -8669 10239 -8617
rect 10291 -8669 10319 -8617
rect 10371 -8669 10399 -8617
rect 10451 -8669 10479 -8617
rect 10531 -8669 10559 -8617
rect 10611 -8669 10620 -8617
rect 9828 -8815 10620 -8669
rect 5759 -8829 10851 -8815
rect 5811 -8881 5839 -8829
rect 5891 -8881 5919 -8829
rect 5971 -8881 5999 -8829
rect 6051 -8881 6079 -8829
rect 6131 -8881 6159 -8829
rect 6211 -8881 6239 -8829
rect 6291 -8881 6319 -8829
rect 6371 -8881 6399 -8829
rect 6451 -8881 6479 -8829
rect 6531 -8881 6559 -8829
rect 6611 -8881 6639 -8829
rect 6691 -8881 6719 -8829
rect 6771 -8881 6799 -8829
rect 6851 -8881 6879 -8829
rect 6931 -8881 6959 -8829
rect 7011 -8881 7039 -8829
rect 7091 -8881 7119 -8829
rect 7171 -8881 7199 -8829
rect 7251 -8881 7279 -8829
rect 7331 -8881 7359 -8829
rect 7411 -8881 7439 -8829
rect 7491 -8881 7519 -8829
rect 7571 -8881 7599 -8829
rect 7651 -8881 7679 -8829
rect 7731 -8881 7759 -8829
rect 7811 -8881 7839 -8829
rect 7891 -8881 7919 -8829
rect 7971 -8881 7999 -8829
rect 8051 -8881 8079 -8829
rect 8131 -8881 8159 -8829
rect 8211 -8881 8239 -8829
rect 8291 -8881 8319 -8829
rect 8371 -8881 8399 -8829
rect 8451 -8881 8479 -8829
rect 8531 -8881 8559 -8829
rect 8611 -8881 8639 -8829
rect 8691 -8881 8719 -8829
rect 8771 -8881 8799 -8829
rect 8851 -8881 8879 -8829
rect 8931 -8881 8959 -8829
rect 9011 -8881 9039 -8829
rect 9091 -8881 9119 -8829
rect 9171 -8881 9199 -8829
rect 9251 -8881 9279 -8829
rect 9331 -8881 9359 -8829
rect 9411 -8881 9439 -8829
rect 9491 -8881 9519 -8829
rect 9571 -8881 9599 -8829
rect 9651 -8881 9679 -8829
rect 9731 -8881 9759 -8829
rect 9811 -8881 9839 -8829
rect 9891 -8881 9919 -8829
rect 9971 -8881 9999 -8829
rect 10051 -8881 10079 -8829
rect 10131 -8881 10159 -8829
rect 10211 -8881 10239 -8829
rect 10291 -8881 10319 -8829
rect 10371 -8881 10399 -8829
rect 10451 -8881 10479 -8829
rect 10531 -8881 10559 -8829
rect 10611 -8881 10639 -8829
rect 10691 -8881 10719 -8829
rect 10771 -8881 10799 -8829
rect 5759 -8909 10851 -8881
rect 5811 -8961 5839 -8909
rect 5891 -8961 5919 -8909
rect 5971 -8961 5999 -8909
rect 6051 -8961 6079 -8909
rect 6131 -8961 6159 -8909
rect 6211 -8961 6239 -8909
rect 6291 -8961 6319 -8909
rect 6371 -8961 6399 -8909
rect 6451 -8961 6479 -8909
rect 6531 -8961 6559 -8909
rect 6611 -8961 6639 -8909
rect 6691 -8961 6719 -8909
rect 6771 -8961 6799 -8909
rect 6851 -8961 6879 -8909
rect 6931 -8961 6959 -8909
rect 7011 -8961 7039 -8909
rect 7091 -8961 7119 -8909
rect 7171 -8961 7199 -8909
rect 7251 -8961 7279 -8909
rect 7331 -8961 7359 -8909
rect 7411 -8961 7439 -8909
rect 7491 -8961 7519 -8909
rect 7571 -8961 7599 -8909
rect 7651 -8961 7679 -8909
rect 7731 -8961 7759 -8909
rect 7811 -8961 7839 -8909
rect 7891 -8961 7919 -8909
rect 7971 -8961 7999 -8909
rect 8051 -8961 8079 -8909
rect 8131 -8961 8159 -8909
rect 8211 -8961 8239 -8909
rect 8291 -8961 8319 -8909
rect 8371 -8961 8399 -8909
rect 8451 -8961 8479 -8909
rect 8531 -8961 8559 -8909
rect 8611 -8961 8639 -8909
rect 8691 -8961 8719 -8909
rect 8771 -8961 8799 -8909
rect 8851 -8961 8879 -8909
rect 8931 -8961 8959 -8909
rect 9011 -8961 9039 -8909
rect 9091 -8961 9119 -8909
rect 9171 -8961 9199 -8909
rect 9251 -8961 9279 -8909
rect 9331 -8961 9359 -8909
rect 9411 -8961 9439 -8909
rect 9491 -8961 9519 -8909
rect 9571 -8961 9599 -8909
rect 9651 -8961 9679 -8909
rect 9731 -8961 9759 -8909
rect 9811 -8961 9839 -8909
rect 9891 -8961 9919 -8909
rect 9971 -8961 9999 -8909
rect 10051 -8961 10079 -8909
rect 10131 -8961 10159 -8909
rect 10211 -8961 10239 -8909
rect 10291 -8961 10319 -8909
rect 10371 -8961 10399 -8909
rect 10451 -8961 10479 -8909
rect 10531 -8961 10559 -8909
rect 10611 -8961 10639 -8909
rect 10691 -8961 10719 -8909
rect 10771 -8961 10799 -8909
rect 5759 -8975 10851 -8961
rect 12523 -9215 12579 -9205
rect 12671 -8365 12727 -8355
rect 12671 -9215 12727 -9205
rect 12819 -8365 12875 -8355
rect 12819 -9215 12875 -9205
rect 12967 -8365 13023 -8355
rect 12967 -9215 13023 -9205
rect 13115 -8365 13171 -8355
rect 13115 -9215 13171 -9205
rect 13263 -8365 13319 -8355
rect 13263 -9215 13319 -9205
rect 13411 -8365 13467 -8355
rect 13411 -9215 13467 -9205
rect 13559 -8365 13615 -8355
rect 13559 -9215 13615 -9205
rect 13707 -8365 13763 -8355
rect 13707 -9215 13763 -9205
rect 13855 -8365 13911 -8355
rect 13855 -9215 13911 -9205
rect 14003 -8365 14059 -8355
rect 14003 -9215 14059 -9205
rect 14151 -8365 14207 -8355
rect 14151 -9215 14207 -9205
rect 14299 -8365 14355 -8355
rect 14299 -9215 14355 -9205
rect 14447 -8365 14503 -8355
rect 14447 -9215 14503 -9205
rect 14595 -8365 14651 -8355
rect 14595 -9215 14651 -9205
rect 14743 -8365 14799 -8355
rect 14743 -9215 14799 -9205
rect 14891 -8365 14947 -8355
rect 14891 -9215 14947 -9205
rect 15039 -8365 15095 -8355
rect 15039 -9215 15095 -9205
rect 15187 -8365 15243 -8355
rect 15187 -9215 15243 -9205
rect 15335 -8365 15391 -8355
rect 15335 -9215 15391 -9205
rect 15483 -8365 15539 -8355
rect 15483 -9215 15539 -9205
rect 15631 -8365 15687 -8355
rect 15631 -9215 15687 -9205
rect 15779 -8365 15835 -8355
rect 15779 -9215 15835 -9205
rect 15927 -8365 15983 -8355
rect 15927 -9215 15983 -9205
rect 16075 -8365 16131 -8355
rect 16075 -9215 16131 -9205
rect 16223 -8365 16279 -8355
rect 16223 -9215 16279 -9205
rect 16371 -8365 16427 -8355
rect 16371 -9215 16427 -9205
rect 16519 -8365 16575 -8355
rect 16519 -9215 16575 -9205
rect 16667 -8365 16723 -8355
rect 16667 -9215 16723 -9205
rect 16815 -8365 16871 -8355
rect 16815 -9215 16871 -9205
rect 16963 -8365 17019 -8355
rect 16963 -9215 17019 -9205
rect 17111 -8365 17167 -8355
rect 17111 -9215 17167 -9205
rect 17259 -8365 17315 -8355
rect 17259 -9215 17315 -9205
rect 17407 -8365 17463 -8355
rect 17407 -9215 17463 -9205
rect 17555 -8365 17611 -8355
rect 17555 -9215 17611 -9205
rect 17703 -8365 17759 -8355
rect 17703 -9215 17759 -9205
rect 17851 -8365 17907 -8355
rect 17851 -9215 17907 -9205
rect 17999 -8365 18055 -8355
rect 17999 -9215 18055 -9205
rect 18147 -8365 18203 -8355
rect 18147 -9215 18203 -9205
rect 18295 -8365 18351 -8355
rect 18295 -9215 18351 -9205
rect 18443 -8365 18499 -8355
rect 18443 -9215 18499 -9205
rect 18591 -8365 18647 -8355
rect 18591 -9215 18647 -9205
rect 18739 -8365 18795 -8355
rect 18739 -9215 18795 -9205
rect 18887 -8365 18943 -8355
rect 18887 -9215 18943 -9205
rect 19035 -8365 19091 -8355
rect 19035 -9215 19091 -9205
rect 19183 -8365 19239 -8355
rect 19183 -9215 19239 -9205
rect 19331 -8365 19387 -8355
rect 19331 -9215 19387 -9205
rect 19479 -8365 19535 -8355
rect 19479 -9215 19535 -9205
rect 19627 -8365 19683 -8355
rect 19627 -9215 19683 -9205
rect 19775 -8365 19831 -8355
rect 19775 -9215 19831 -9205
rect 19923 -8365 19979 -8355
rect 19923 -9215 19979 -9205
rect 20071 -8365 20127 -8355
rect 20071 -9215 20127 -9205
rect 20219 -8365 20275 -8355
rect 20219 -9215 20275 -9205
rect 20367 -8365 20423 -8355
rect 20367 -9215 20423 -9205
rect 20515 -8365 20571 -8355
rect 20515 -9215 20571 -9205
rect 20663 -8365 20719 -8355
rect 20663 -9215 20719 -9205
rect 20811 -8365 20867 -8355
rect 20811 -9215 20867 -9205
rect 20959 -8365 21015 -8355
rect 20959 -9215 21015 -9205
rect 21107 -8365 21163 -8355
rect 21107 -9215 21163 -9205
rect 21255 -8365 21311 -8355
rect 21255 -9215 21311 -9205
rect 21403 -8365 21459 -8355
rect 21403 -9215 21459 -9205
rect 21551 -8365 21607 -8355
rect 21551 -9215 21607 -9205
rect 21699 -8365 21755 -8355
rect 21699 -9215 21755 -9205
rect 21847 -8365 21903 -8355
rect 21847 -9215 21903 -9205
rect 21995 -8365 22051 -8355
rect 21995 -9215 22051 -9205
rect 22143 -8365 22199 -8355
rect 22143 -9215 22199 -9205
rect 22291 -8365 22347 -8355
rect 22291 -9215 22347 -9205
rect 22439 -8365 22495 -8355
rect 22439 -9215 22495 -9205
rect 22587 -8365 22643 -8355
rect 22587 -9215 22643 -9205
rect 22735 -8365 22791 -8355
rect 22735 -9215 22791 -9205
rect 22883 -8365 22939 -8355
rect 22883 -9215 22939 -9205
rect 23031 -8365 23087 -8355
rect 23031 -9215 23087 -9205
rect 23179 -8365 23235 -8355
rect 23179 -9215 23235 -9205
rect 23327 -8365 23383 -8355
rect 23327 -9215 23383 -9205
rect 23475 -8365 23531 -8355
rect 23475 -9215 23531 -9205
rect 23623 -8365 23679 -8355
rect 23623 -9215 23679 -9205
rect 4044 -9681 26275 -9673
rect 4044 -9737 4053 -9681
rect 4109 -9737 4134 -9681
rect 4190 -9737 4215 -9681
rect 4271 -9737 4296 -9681
rect 4352 -9737 4377 -9681
rect 4433 -9737 4458 -9681
rect 4514 -9737 4539 -9681
rect 4595 -9737 4621 -9681
rect 4677 -9737 4702 -9681
rect 4758 -9737 4783 -9681
rect 4839 -9737 4864 -9681
rect 4920 -9737 4945 -9681
rect 5001 -9737 5026 -9681
rect 5082 -9737 5107 -9681
rect 5163 -9737 5189 -9681
rect 5245 -9737 5270 -9681
rect 5326 -9737 5351 -9681
rect 5407 -9737 5432 -9681
rect 5488 -9737 5513 -9681
rect 5569 -9737 5594 -9681
rect 5650 -9737 5675 -9681
rect 5731 -9737 5757 -9681
rect 5813 -9737 5838 -9681
rect 5894 -9737 5919 -9681
rect 5975 -9737 6000 -9681
rect 6056 -9737 6081 -9681
rect 6137 -9737 6162 -9681
rect 6218 -9737 6243 -9681
rect 6299 -9737 6325 -9681
rect 6381 -9737 6406 -9681
rect 6462 -9737 6487 -9681
rect 6543 -9737 6568 -9681
rect 6624 -9737 6649 -9681
rect 6705 -9737 6730 -9681
rect 6786 -9737 6811 -9681
rect 6867 -9737 6893 -9681
rect 6949 -9737 6974 -9681
rect 7030 -9737 7055 -9681
rect 7111 -9737 7136 -9681
rect 7192 -9737 7217 -9681
rect 7273 -9737 7298 -9681
rect 7354 -9737 7379 -9681
rect 7435 -9737 7461 -9681
rect 7517 -9737 7542 -9681
rect 7598 -9737 7623 -9681
rect 7679 -9737 7704 -9681
rect 7760 -9737 7785 -9681
rect 7841 -9737 7866 -9681
rect 7922 -9737 7947 -9681
rect 8003 -9737 8029 -9681
rect 8085 -9737 8110 -9681
rect 8166 -9737 8191 -9681
rect 8247 -9737 8272 -9681
rect 8328 -9737 8353 -9681
rect 8409 -9737 8434 -9681
rect 8490 -9737 8515 -9681
rect 8571 -9737 8597 -9681
rect 8653 -9737 8678 -9681
rect 8734 -9737 8759 -9681
rect 8815 -9737 8840 -9681
rect 8896 -9737 8921 -9681
rect 8977 -9737 9002 -9681
rect 9058 -9737 9083 -9681
rect 9139 -9737 9165 -9681
rect 9221 -9737 9246 -9681
rect 9302 -9737 9327 -9681
rect 9383 -9737 9408 -9681
rect 9464 -9737 9489 -9681
rect 9545 -9737 9570 -9681
rect 9626 -9737 9651 -9681
rect 9707 -9737 9733 -9681
rect 9789 -9737 9814 -9681
rect 9870 -9737 9895 -9681
rect 9951 -9737 9976 -9681
rect 10032 -9737 10057 -9681
rect 10113 -9737 10138 -9681
rect 10194 -9737 10219 -9681
rect 10275 -9737 10301 -9681
rect 10357 -9737 10382 -9681
rect 10438 -9737 10463 -9681
rect 10519 -9737 10544 -9681
rect 10600 -9737 10625 -9681
rect 10681 -9737 10706 -9681
rect 10762 -9737 10787 -9681
rect 10843 -9737 10869 -9681
rect 10925 -9737 10950 -9681
rect 11006 -9737 11031 -9681
rect 11087 -9737 11112 -9681
rect 11168 -9737 11193 -9681
rect 11249 -9737 11274 -9681
rect 11330 -9737 11355 -9681
rect 11411 -9737 11437 -9681
rect 11493 -9737 11518 -9681
rect 11574 -9737 11599 -9681
rect 11655 -9737 11680 -9681
rect 11736 -9737 11761 -9681
rect 11817 -9737 11842 -9681
rect 11898 -9737 11923 -9681
rect 11979 -9737 12005 -9681
rect 12061 -9737 12086 -9681
rect 12142 -9737 12167 -9681
rect 12223 -9737 12248 -9681
rect 12304 -9737 12329 -9681
rect 12385 -9737 12410 -9681
rect 12466 -9737 12491 -9681
rect 12547 -9737 12573 -9681
rect 12629 -9737 12654 -9681
rect 12710 -9737 12735 -9681
rect 12791 -9737 12816 -9681
rect 12872 -9737 12897 -9681
rect 12953 -9737 12978 -9681
rect 13034 -9737 13059 -9681
rect 13115 -9737 13141 -9681
rect 13197 -9737 13222 -9681
rect 13278 -9737 13303 -9681
rect 13359 -9737 13384 -9681
rect 13440 -9737 13465 -9681
rect 13521 -9737 13546 -9681
rect 13602 -9737 13627 -9681
rect 13683 -9737 13709 -9681
rect 13765 -9737 13790 -9681
rect 13846 -9737 13871 -9681
rect 13927 -9737 13952 -9681
rect 14008 -9737 14033 -9681
rect 14089 -9737 14114 -9681
rect 14170 -9737 14195 -9681
rect 14251 -9737 14277 -9681
rect 14333 -9737 14358 -9681
rect 14414 -9737 14439 -9681
rect 14495 -9737 14520 -9681
rect 14576 -9737 14601 -9681
rect 14657 -9737 14682 -9681
rect 14738 -9737 14763 -9681
rect 14819 -9737 14845 -9681
rect 14901 -9737 14926 -9681
rect 14982 -9737 15007 -9681
rect 15063 -9737 15088 -9681
rect 15144 -9737 15169 -9681
rect 15225 -9737 15250 -9681
rect 15306 -9737 15331 -9681
rect 15387 -9737 15413 -9681
rect 15469 -9737 15494 -9681
rect 15550 -9737 15575 -9681
rect 15631 -9737 15656 -9681
rect 15712 -9737 15737 -9681
rect 15793 -9737 15818 -9681
rect 15874 -9737 15899 -9681
rect 15955 -9737 15981 -9681
rect 16037 -9737 16062 -9681
rect 16118 -9737 16143 -9681
rect 16199 -9737 16224 -9681
rect 16280 -9737 16305 -9681
rect 16361 -9737 16386 -9681
rect 16442 -9737 16467 -9681
rect 16523 -9737 16549 -9681
rect 16605 -9737 16630 -9681
rect 16686 -9737 16711 -9681
rect 16767 -9737 16792 -9681
rect 16848 -9737 16873 -9681
rect 16929 -9737 16954 -9681
rect 17010 -9737 17035 -9681
rect 17091 -9737 17117 -9681
rect 17173 -9737 17198 -9681
rect 17254 -9737 17279 -9681
rect 17335 -9737 17360 -9681
rect 17416 -9737 17441 -9681
rect 17497 -9737 17522 -9681
rect 17578 -9737 17603 -9681
rect 17659 -9737 17684 -9681
rect 17740 -9737 17765 -9681
rect 17821 -9737 17846 -9681
rect 17902 -9737 17927 -9681
rect 17983 -9737 18008 -9681
rect 18064 -9737 18089 -9681
rect 18145 -9737 18171 -9681
rect 18227 -9737 18252 -9681
rect 18308 -9737 18333 -9681
rect 18389 -9737 18414 -9681
rect 18470 -9737 18495 -9681
rect 18551 -9737 18576 -9681
rect 18632 -9737 18657 -9681
rect 18713 -9737 18739 -9681
rect 18795 -9737 18820 -9681
rect 18876 -9737 18901 -9681
rect 18957 -9737 18982 -9681
rect 19038 -9737 19063 -9681
rect 19119 -9737 19144 -9681
rect 19200 -9737 19225 -9681
rect 19281 -9737 19307 -9681
rect 19363 -9737 19388 -9681
rect 19444 -9737 19469 -9681
rect 19525 -9737 19550 -9681
rect 19606 -9737 19631 -9681
rect 19687 -9737 19712 -9681
rect 19768 -9737 19793 -9681
rect 19849 -9737 19875 -9681
rect 19931 -9737 19956 -9681
rect 20012 -9737 20037 -9681
rect 20093 -9737 20118 -9681
rect 20174 -9737 20199 -9681
rect 20255 -9737 20280 -9681
rect 20336 -9737 20361 -9681
rect 20417 -9737 20443 -9681
rect 20499 -9737 20524 -9681
rect 20580 -9737 20605 -9681
rect 20661 -9737 20686 -9681
rect 20742 -9737 20767 -9681
rect 20823 -9737 20848 -9681
rect 20904 -9737 20929 -9681
rect 20985 -9737 21011 -9681
rect 21067 -9737 21092 -9681
rect 21148 -9737 21173 -9681
rect 21229 -9737 21254 -9681
rect 21310 -9737 21335 -9681
rect 21391 -9737 21416 -9681
rect 21472 -9737 21497 -9681
rect 21553 -9737 21579 -9681
rect 21635 -9737 21660 -9681
rect 21716 -9737 21741 -9681
rect 21797 -9737 21822 -9681
rect 21878 -9737 21903 -9681
rect 21959 -9737 21984 -9681
rect 22040 -9737 22065 -9681
rect 22121 -9737 22147 -9681
rect 22203 -9737 22228 -9681
rect 22284 -9737 22309 -9681
rect 22365 -9737 22390 -9681
rect 22446 -9737 22471 -9681
rect 22527 -9737 22552 -9681
rect 22608 -9737 22633 -9681
rect 22689 -9737 22715 -9681
rect 22771 -9737 22796 -9681
rect 22852 -9737 22877 -9681
rect 22933 -9737 22958 -9681
rect 23014 -9737 23039 -9681
rect 23095 -9737 23120 -9681
rect 23176 -9737 23201 -9681
rect 23257 -9737 23283 -9681
rect 23339 -9737 23364 -9681
rect 23420 -9737 23445 -9681
rect 23501 -9737 23526 -9681
rect 23582 -9737 23607 -9681
rect 23663 -9737 23688 -9681
rect 23744 -9737 23769 -9681
rect 23825 -9737 23851 -9681
rect 23907 -9737 23932 -9681
rect 23988 -9737 24013 -9681
rect 24069 -9737 24094 -9681
rect 24150 -9737 24175 -9681
rect 24231 -9737 24256 -9681
rect 24312 -9737 24337 -9681
rect 24393 -9737 24419 -9681
rect 24475 -9737 24500 -9681
rect 24556 -9737 24581 -9681
rect 24637 -9737 24662 -9681
rect 24718 -9737 24743 -9681
rect 24799 -9737 24824 -9681
rect 24880 -9737 24905 -9681
rect 24961 -9737 24987 -9681
rect 25043 -9737 25068 -9681
rect 25124 -9737 25149 -9681
rect 25205 -9737 25230 -9681
rect 25286 -9737 25311 -9681
rect 25367 -9737 25392 -9681
rect 25448 -9737 25473 -9681
rect 25529 -9737 25555 -9681
rect 25611 -9737 25636 -9681
rect 25692 -9737 25717 -9681
rect 25773 -9737 25798 -9681
rect 25854 -9737 25879 -9681
rect 25935 -9737 25960 -9681
rect 26016 -9737 26041 -9681
rect 26097 -9737 26123 -9681
rect 26179 -9737 26204 -9681
rect 26260 -9737 26275 -9681
rect 4044 -9785 26275 -9737
rect 4044 -9841 4053 -9785
rect 4109 -9841 4134 -9785
rect 4190 -9841 4215 -9785
rect 4271 -9841 4296 -9785
rect 4352 -9841 4377 -9785
rect 4433 -9841 4458 -9785
rect 4514 -9841 4539 -9785
rect 4595 -9841 4621 -9785
rect 4677 -9841 4702 -9785
rect 4758 -9841 4783 -9785
rect 4839 -9841 4864 -9785
rect 4920 -9841 4945 -9785
rect 5001 -9841 5026 -9785
rect 5082 -9841 5107 -9785
rect 5163 -9841 5189 -9785
rect 5245 -9841 5270 -9785
rect 5326 -9841 5351 -9785
rect 5407 -9841 5432 -9785
rect 5488 -9841 5513 -9785
rect 5569 -9841 5594 -9785
rect 5650 -9841 5675 -9785
rect 5731 -9841 5757 -9785
rect 5813 -9841 5838 -9785
rect 5894 -9841 5919 -9785
rect 5975 -9841 6000 -9785
rect 6056 -9841 6081 -9785
rect 6137 -9841 6162 -9785
rect 6218 -9841 6243 -9785
rect 6299 -9841 6325 -9785
rect 6381 -9841 6406 -9785
rect 6462 -9841 6487 -9785
rect 6543 -9841 6568 -9785
rect 6624 -9841 6649 -9785
rect 6705 -9841 6730 -9785
rect 6786 -9841 6811 -9785
rect 6867 -9841 6893 -9785
rect 6949 -9841 6974 -9785
rect 7030 -9841 7055 -9785
rect 7111 -9841 7136 -9785
rect 7192 -9841 7217 -9785
rect 7273 -9841 7298 -9785
rect 7354 -9841 7379 -9785
rect 7435 -9841 7461 -9785
rect 7517 -9841 7542 -9785
rect 7598 -9841 7623 -9785
rect 7679 -9841 7704 -9785
rect 7760 -9841 7785 -9785
rect 7841 -9841 7866 -9785
rect 7922 -9841 7947 -9785
rect 8003 -9841 8029 -9785
rect 8085 -9841 8110 -9785
rect 8166 -9841 8191 -9785
rect 8247 -9841 8272 -9785
rect 8328 -9841 8353 -9785
rect 8409 -9841 8434 -9785
rect 8490 -9841 8515 -9785
rect 8571 -9841 8597 -9785
rect 8653 -9841 8678 -9785
rect 8734 -9841 8759 -9785
rect 8815 -9841 8840 -9785
rect 8896 -9841 8921 -9785
rect 8977 -9841 9002 -9785
rect 9058 -9841 9083 -9785
rect 9139 -9841 9165 -9785
rect 9221 -9841 9246 -9785
rect 9302 -9841 9327 -9785
rect 9383 -9841 9408 -9785
rect 9464 -9841 9489 -9785
rect 9545 -9841 9570 -9785
rect 9626 -9841 9651 -9785
rect 9707 -9841 9733 -9785
rect 9789 -9841 9814 -9785
rect 9870 -9841 9895 -9785
rect 9951 -9841 9976 -9785
rect 10032 -9841 10057 -9785
rect 10113 -9841 10138 -9785
rect 10194 -9841 10219 -9785
rect 10275 -9841 10301 -9785
rect 10357 -9841 10382 -9785
rect 10438 -9841 10463 -9785
rect 10519 -9841 10544 -9785
rect 10600 -9841 10625 -9785
rect 10681 -9841 10706 -9785
rect 10762 -9841 10787 -9785
rect 10843 -9841 10869 -9785
rect 10925 -9841 10950 -9785
rect 11006 -9841 11031 -9785
rect 11087 -9841 11112 -9785
rect 11168 -9841 11193 -9785
rect 11249 -9841 11274 -9785
rect 11330 -9841 11355 -9785
rect 11411 -9841 11437 -9785
rect 11493 -9841 11518 -9785
rect 11574 -9841 11599 -9785
rect 11655 -9841 11680 -9785
rect 11736 -9841 11761 -9785
rect 11817 -9841 11842 -9785
rect 11898 -9841 11923 -9785
rect 11979 -9841 12005 -9785
rect 12061 -9841 12086 -9785
rect 12142 -9841 12167 -9785
rect 12223 -9841 12248 -9785
rect 12304 -9841 12329 -9785
rect 12385 -9841 12410 -9785
rect 12466 -9841 12491 -9785
rect 12547 -9841 12573 -9785
rect 12629 -9841 12654 -9785
rect 12710 -9841 12735 -9785
rect 12791 -9841 12816 -9785
rect 12872 -9841 12897 -9785
rect 12953 -9841 12978 -9785
rect 13034 -9841 13059 -9785
rect 13115 -9841 13141 -9785
rect 13197 -9841 13222 -9785
rect 13278 -9841 13303 -9785
rect 13359 -9841 13384 -9785
rect 13440 -9841 13465 -9785
rect 13521 -9841 13546 -9785
rect 13602 -9841 13627 -9785
rect 13683 -9841 13709 -9785
rect 13765 -9841 13790 -9785
rect 13846 -9841 13871 -9785
rect 13927 -9841 13952 -9785
rect 14008 -9841 14033 -9785
rect 14089 -9841 14114 -9785
rect 14170 -9841 14195 -9785
rect 14251 -9841 14277 -9785
rect 14333 -9841 14358 -9785
rect 14414 -9841 14439 -9785
rect 14495 -9841 14520 -9785
rect 14576 -9841 14601 -9785
rect 14657 -9841 14682 -9785
rect 14738 -9841 14763 -9785
rect 14819 -9841 14845 -9785
rect 14901 -9841 14926 -9785
rect 14982 -9841 15007 -9785
rect 15063 -9841 15088 -9785
rect 15144 -9841 15169 -9785
rect 15225 -9841 15250 -9785
rect 15306 -9841 15331 -9785
rect 15387 -9841 15413 -9785
rect 15469 -9841 15494 -9785
rect 15550 -9841 15575 -9785
rect 15631 -9841 15656 -9785
rect 15712 -9841 15737 -9785
rect 15793 -9841 15818 -9785
rect 15874 -9841 15899 -9785
rect 15955 -9841 15981 -9785
rect 16037 -9841 16062 -9785
rect 16118 -9841 16143 -9785
rect 16199 -9841 16224 -9785
rect 16280 -9841 16305 -9785
rect 16361 -9841 16386 -9785
rect 16442 -9841 16467 -9785
rect 16523 -9841 16549 -9785
rect 16605 -9841 16630 -9785
rect 16686 -9841 16711 -9785
rect 16767 -9841 16792 -9785
rect 16848 -9841 16873 -9785
rect 16929 -9841 16954 -9785
rect 17010 -9841 17035 -9785
rect 17091 -9841 17117 -9785
rect 17173 -9841 17198 -9785
rect 17254 -9841 17279 -9785
rect 17335 -9841 17360 -9785
rect 17416 -9841 17441 -9785
rect 17497 -9841 17522 -9785
rect 17578 -9841 17603 -9785
rect 17659 -9841 17684 -9785
rect 17740 -9841 17765 -9785
rect 17821 -9841 17846 -9785
rect 17902 -9841 17927 -9785
rect 17983 -9841 18008 -9785
rect 18064 -9841 18089 -9785
rect 18145 -9841 18171 -9785
rect 18227 -9841 18252 -9785
rect 18308 -9841 18333 -9785
rect 18389 -9841 18414 -9785
rect 18470 -9841 18495 -9785
rect 18551 -9841 18576 -9785
rect 18632 -9841 18657 -9785
rect 18713 -9841 18739 -9785
rect 18795 -9841 18820 -9785
rect 18876 -9841 18901 -9785
rect 18957 -9841 18982 -9785
rect 19038 -9841 19063 -9785
rect 19119 -9841 19144 -9785
rect 19200 -9841 19225 -9785
rect 19281 -9841 19307 -9785
rect 19363 -9841 19388 -9785
rect 19444 -9841 19469 -9785
rect 19525 -9841 19550 -9785
rect 19606 -9841 19631 -9785
rect 19687 -9841 19712 -9785
rect 19768 -9841 19793 -9785
rect 19849 -9841 19875 -9785
rect 19931 -9841 19956 -9785
rect 20012 -9841 20037 -9785
rect 20093 -9841 20118 -9785
rect 20174 -9841 20199 -9785
rect 20255 -9841 20280 -9785
rect 20336 -9841 20361 -9785
rect 20417 -9841 20443 -9785
rect 20499 -9841 20524 -9785
rect 20580 -9841 20605 -9785
rect 20661 -9841 20686 -9785
rect 20742 -9841 20767 -9785
rect 20823 -9841 20848 -9785
rect 20904 -9841 20929 -9785
rect 20985 -9841 21011 -9785
rect 21067 -9841 21092 -9785
rect 21148 -9841 21173 -9785
rect 21229 -9841 21254 -9785
rect 21310 -9841 21335 -9785
rect 21391 -9841 21416 -9785
rect 21472 -9841 21497 -9785
rect 21553 -9841 21579 -9785
rect 21635 -9841 21660 -9785
rect 21716 -9841 21741 -9785
rect 21797 -9841 21822 -9785
rect 21878 -9841 21903 -9785
rect 21959 -9841 21984 -9785
rect 22040 -9841 22065 -9785
rect 22121 -9841 22147 -9785
rect 22203 -9841 22228 -9785
rect 22284 -9841 22309 -9785
rect 22365 -9841 22390 -9785
rect 22446 -9841 22471 -9785
rect 22527 -9841 22552 -9785
rect 22608 -9841 22633 -9785
rect 22689 -9841 22715 -9785
rect 22771 -9841 22796 -9785
rect 22852 -9841 22877 -9785
rect 22933 -9841 22958 -9785
rect 23014 -9841 23039 -9785
rect 23095 -9841 23120 -9785
rect 23176 -9841 23201 -9785
rect 23257 -9841 23283 -9785
rect 23339 -9841 23364 -9785
rect 23420 -9841 23445 -9785
rect 23501 -9841 23526 -9785
rect 23582 -9841 23607 -9785
rect 23663 -9841 23688 -9785
rect 23744 -9841 23769 -9785
rect 23825 -9841 23851 -9785
rect 23907 -9841 23932 -9785
rect 23988 -9841 24013 -9785
rect 24069 -9841 24094 -9785
rect 24150 -9841 24175 -9785
rect 24231 -9841 24256 -9785
rect 24312 -9841 24337 -9785
rect 24393 -9841 24419 -9785
rect 24475 -9841 24500 -9785
rect 24556 -9841 24581 -9785
rect 24637 -9841 24662 -9785
rect 24718 -9841 24743 -9785
rect 24799 -9841 24824 -9785
rect 24880 -9841 24905 -9785
rect 24961 -9841 24987 -9785
rect 25043 -9841 25068 -9785
rect 25124 -9841 25149 -9785
rect 25205 -9841 25230 -9785
rect 25286 -9841 25311 -9785
rect 25367 -9841 25392 -9785
rect 25448 -9841 25473 -9785
rect 25529 -9841 25555 -9785
rect 25611 -9841 25636 -9785
rect 25692 -9841 25717 -9785
rect 25773 -9841 25798 -9785
rect 25854 -9841 25879 -9785
rect 25935 -9841 25960 -9785
rect 26016 -9841 26041 -9785
rect 26097 -9841 26123 -9785
rect 26179 -9841 26204 -9785
rect 26260 -9841 26275 -9785
rect 4044 -9889 26275 -9841
rect 4044 -9945 4053 -9889
rect 4109 -9945 4134 -9889
rect 4190 -9945 4215 -9889
rect 4271 -9945 4296 -9889
rect 4352 -9945 4377 -9889
rect 4433 -9945 4458 -9889
rect 4514 -9945 4539 -9889
rect 4595 -9945 4621 -9889
rect 4677 -9945 4702 -9889
rect 4758 -9945 4783 -9889
rect 4839 -9945 4864 -9889
rect 4920 -9945 4945 -9889
rect 5001 -9945 5026 -9889
rect 5082 -9945 5107 -9889
rect 5163 -9945 5189 -9889
rect 5245 -9945 5270 -9889
rect 5326 -9945 5351 -9889
rect 5407 -9945 5432 -9889
rect 5488 -9945 5513 -9889
rect 5569 -9945 5594 -9889
rect 5650 -9945 5675 -9889
rect 5731 -9945 5757 -9889
rect 5813 -9945 5838 -9889
rect 5894 -9945 5919 -9889
rect 5975 -9945 6000 -9889
rect 6056 -9945 6081 -9889
rect 6137 -9945 6162 -9889
rect 6218 -9945 6243 -9889
rect 6299 -9945 6325 -9889
rect 6381 -9945 6406 -9889
rect 6462 -9945 6487 -9889
rect 6543 -9945 6568 -9889
rect 6624 -9945 6649 -9889
rect 6705 -9945 6730 -9889
rect 6786 -9945 6811 -9889
rect 6867 -9945 6893 -9889
rect 6949 -9945 6974 -9889
rect 7030 -9945 7055 -9889
rect 7111 -9945 7136 -9889
rect 7192 -9945 7217 -9889
rect 7273 -9945 7298 -9889
rect 7354 -9945 7379 -9889
rect 7435 -9945 7461 -9889
rect 7517 -9945 7542 -9889
rect 7598 -9945 7623 -9889
rect 7679 -9945 7704 -9889
rect 7760 -9945 7785 -9889
rect 7841 -9945 7866 -9889
rect 7922 -9945 7947 -9889
rect 8003 -9945 8029 -9889
rect 8085 -9945 8110 -9889
rect 8166 -9945 8191 -9889
rect 8247 -9945 8272 -9889
rect 8328 -9945 8353 -9889
rect 8409 -9945 8434 -9889
rect 8490 -9945 8515 -9889
rect 8571 -9945 8597 -9889
rect 8653 -9945 8678 -9889
rect 8734 -9945 8759 -9889
rect 8815 -9945 8840 -9889
rect 8896 -9945 8921 -9889
rect 8977 -9945 9002 -9889
rect 9058 -9945 9083 -9889
rect 9139 -9945 9165 -9889
rect 9221 -9945 9246 -9889
rect 9302 -9945 9327 -9889
rect 9383 -9945 9408 -9889
rect 9464 -9945 9489 -9889
rect 9545 -9945 9570 -9889
rect 9626 -9945 9651 -9889
rect 9707 -9945 9733 -9889
rect 9789 -9945 9814 -9889
rect 9870 -9945 9895 -9889
rect 9951 -9945 9976 -9889
rect 10032 -9945 10057 -9889
rect 10113 -9945 10138 -9889
rect 10194 -9945 10219 -9889
rect 10275 -9945 10301 -9889
rect 10357 -9945 10382 -9889
rect 10438 -9945 10463 -9889
rect 10519 -9945 10544 -9889
rect 10600 -9945 10625 -9889
rect 10681 -9945 10706 -9889
rect 10762 -9945 10787 -9889
rect 10843 -9945 10869 -9889
rect 10925 -9945 10950 -9889
rect 11006 -9945 11031 -9889
rect 11087 -9945 11112 -9889
rect 11168 -9945 11193 -9889
rect 11249 -9945 11274 -9889
rect 11330 -9945 11355 -9889
rect 11411 -9945 11437 -9889
rect 11493 -9945 11518 -9889
rect 11574 -9945 11599 -9889
rect 11655 -9945 11680 -9889
rect 11736 -9945 11761 -9889
rect 11817 -9945 11842 -9889
rect 11898 -9945 11923 -9889
rect 11979 -9945 12005 -9889
rect 12061 -9945 12086 -9889
rect 12142 -9945 12167 -9889
rect 12223 -9945 12248 -9889
rect 12304 -9945 12329 -9889
rect 12385 -9945 12410 -9889
rect 12466 -9945 12491 -9889
rect 12547 -9945 12573 -9889
rect 12629 -9945 12654 -9889
rect 12710 -9945 12735 -9889
rect 12791 -9945 12816 -9889
rect 12872 -9945 12897 -9889
rect 12953 -9945 12978 -9889
rect 13034 -9945 13059 -9889
rect 13115 -9945 13141 -9889
rect 13197 -9945 13222 -9889
rect 13278 -9945 13303 -9889
rect 13359 -9945 13384 -9889
rect 13440 -9945 13465 -9889
rect 13521 -9945 13546 -9889
rect 13602 -9945 13627 -9889
rect 13683 -9945 13709 -9889
rect 13765 -9945 13790 -9889
rect 13846 -9945 13871 -9889
rect 13927 -9945 13952 -9889
rect 14008 -9945 14033 -9889
rect 14089 -9945 14114 -9889
rect 14170 -9945 14195 -9889
rect 14251 -9945 14277 -9889
rect 14333 -9945 14358 -9889
rect 14414 -9945 14439 -9889
rect 14495 -9945 14520 -9889
rect 14576 -9945 14601 -9889
rect 14657 -9945 14682 -9889
rect 14738 -9945 14763 -9889
rect 14819 -9945 14845 -9889
rect 14901 -9945 14926 -9889
rect 14982 -9945 15007 -9889
rect 15063 -9945 15088 -9889
rect 15144 -9945 15169 -9889
rect 15225 -9945 15250 -9889
rect 15306 -9945 15331 -9889
rect 15387 -9945 15413 -9889
rect 15469 -9945 15494 -9889
rect 15550 -9945 15575 -9889
rect 15631 -9945 15656 -9889
rect 15712 -9945 15737 -9889
rect 15793 -9945 15818 -9889
rect 15874 -9945 15899 -9889
rect 15955 -9945 15981 -9889
rect 16037 -9945 16062 -9889
rect 16118 -9945 16143 -9889
rect 16199 -9945 16224 -9889
rect 16280 -9945 16305 -9889
rect 16361 -9945 16386 -9889
rect 16442 -9945 16467 -9889
rect 16523 -9945 16549 -9889
rect 16605 -9945 16630 -9889
rect 16686 -9945 16711 -9889
rect 16767 -9945 16792 -9889
rect 16848 -9945 16873 -9889
rect 16929 -9945 16954 -9889
rect 17010 -9945 17035 -9889
rect 17091 -9945 17117 -9889
rect 17173 -9945 17198 -9889
rect 17254 -9945 17279 -9889
rect 17335 -9945 17360 -9889
rect 17416 -9945 17441 -9889
rect 17497 -9945 17522 -9889
rect 17578 -9945 17603 -9889
rect 17659 -9945 17684 -9889
rect 17740 -9945 17765 -9889
rect 17821 -9945 17846 -9889
rect 17902 -9945 17927 -9889
rect 17983 -9945 18008 -9889
rect 18064 -9945 18089 -9889
rect 18145 -9945 18171 -9889
rect 18227 -9945 18252 -9889
rect 18308 -9945 18333 -9889
rect 18389 -9945 18414 -9889
rect 18470 -9945 18495 -9889
rect 18551 -9945 18576 -9889
rect 18632 -9945 18657 -9889
rect 18713 -9945 18739 -9889
rect 18795 -9945 18820 -9889
rect 18876 -9945 18901 -9889
rect 18957 -9945 18982 -9889
rect 19038 -9945 19063 -9889
rect 19119 -9945 19144 -9889
rect 19200 -9945 19225 -9889
rect 19281 -9945 19307 -9889
rect 19363 -9945 19388 -9889
rect 19444 -9945 19469 -9889
rect 19525 -9945 19550 -9889
rect 19606 -9945 19631 -9889
rect 19687 -9945 19712 -9889
rect 19768 -9945 19793 -9889
rect 19849 -9945 19875 -9889
rect 19931 -9945 19956 -9889
rect 20012 -9945 20037 -9889
rect 20093 -9945 20118 -9889
rect 20174 -9945 20199 -9889
rect 20255 -9945 20280 -9889
rect 20336 -9945 20361 -9889
rect 20417 -9945 20443 -9889
rect 20499 -9945 20524 -9889
rect 20580 -9945 20605 -9889
rect 20661 -9945 20686 -9889
rect 20742 -9945 20767 -9889
rect 20823 -9945 20848 -9889
rect 20904 -9945 20929 -9889
rect 20985 -9945 21011 -9889
rect 21067 -9945 21092 -9889
rect 21148 -9945 21173 -9889
rect 21229 -9945 21254 -9889
rect 21310 -9945 21335 -9889
rect 21391 -9945 21416 -9889
rect 21472 -9945 21497 -9889
rect 21553 -9945 21579 -9889
rect 21635 -9945 21660 -9889
rect 21716 -9945 21741 -9889
rect 21797 -9945 21822 -9889
rect 21878 -9945 21903 -9889
rect 21959 -9945 21984 -9889
rect 22040 -9945 22065 -9889
rect 22121 -9945 22147 -9889
rect 22203 -9945 22228 -9889
rect 22284 -9945 22309 -9889
rect 22365 -9945 22390 -9889
rect 22446 -9945 22471 -9889
rect 22527 -9945 22552 -9889
rect 22608 -9945 22633 -9889
rect 22689 -9945 22715 -9889
rect 22771 -9945 22796 -9889
rect 22852 -9945 22877 -9889
rect 22933 -9945 22958 -9889
rect 23014 -9945 23039 -9889
rect 23095 -9945 23120 -9889
rect 23176 -9945 23201 -9889
rect 23257 -9945 23283 -9889
rect 23339 -9945 23364 -9889
rect 23420 -9945 23445 -9889
rect 23501 -9945 23526 -9889
rect 23582 -9945 23607 -9889
rect 23663 -9945 23688 -9889
rect 23744 -9945 23769 -9889
rect 23825 -9945 23851 -9889
rect 23907 -9945 23932 -9889
rect 23988 -9945 24013 -9889
rect 24069 -9945 24094 -9889
rect 24150 -9945 24175 -9889
rect 24231 -9945 24256 -9889
rect 24312 -9945 24337 -9889
rect 24393 -9945 24419 -9889
rect 24475 -9945 24500 -9889
rect 24556 -9945 24581 -9889
rect 24637 -9945 24662 -9889
rect 24718 -9945 24743 -9889
rect 24799 -9945 24824 -9889
rect 24880 -9945 24905 -9889
rect 24961 -9945 24987 -9889
rect 25043 -9945 25068 -9889
rect 25124 -9945 25149 -9889
rect 25205 -9945 25230 -9889
rect 25286 -9945 25311 -9889
rect 25367 -9945 25392 -9889
rect 25448 -9945 25473 -9889
rect 25529 -9945 25555 -9889
rect 25611 -9945 25636 -9889
rect 25692 -9945 25717 -9889
rect 25773 -9945 25798 -9889
rect 25854 -9945 25879 -9889
rect 25935 -9945 25960 -9889
rect 26016 -9945 26041 -9889
rect 26097 -9945 26123 -9889
rect 26179 -9945 26204 -9889
rect 26260 -9945 26275 -9889
rect 4044 -9950 26275 -9945
<< via2 >>
rect 3036 3172 3092 3174
rect 3036 3120 3038 3172
rect 3038 3120 3090 3172
rect 3090 3120 3092 3172
rect 3036 3118 3092 3120
rect 3118 3172 3174 3174
rect 3118 3120 3120 3172
rect 3120 3120 3172 3172
rect 3172 3120 3174 3172
rect 3118 3118 3174 3120
rect 3199 3172 3255 3174
rect 3199 3120 3201 3172
rect 3201 3120 3253 3172
rect 3253 3120 3255 3172
rect 3199 3118 3255 3120
rect 3280 3172 3336 3174
rect 3280 3120 3282 3172
rect 3282 3120 3334 3172
rect 3334 3120 3336 3172
rect 3280 3118 3336 3120
rect 3361 3172 3417 3174
rect 3361 3120 3363 3172
rect 3363 3120 3415 3172
rect 3415 3120 3417 3172
rect 3361 3118 3417 3120
rect 3442 3172 3498 3174
rect 3442 3120 3444 3172
rect 3444 3120 3496 3172
rect 3496 3120 3498 3172
rect 3442 3118 3498 3120
rect 3523 3172 3579 3174
rect 3523 3120 3525 3172
rect 3525 3120 3577 3172
rect 3577 3120 3579 3172
rect 3523 3118 3579 3120
rect 3604 3172 3660 3174
rect 3604 3120 3606 3172
rect 3606 3120 3658 3172
rect 3658 3120 3660 3172
rect 3604 3118 3660 3120
rect 3686 3172 3742 3174
rect 3686 3120 3688 3172
rect 3688 3120 3740 3172
rect 3740 3120 3742 3172
rect 3686 3118 3742 3120
rect 3767 3172 3823 3174
rect 3767 3120 3769 3172
rect 3769 3120 3821 3172
rect 3821 3120 3823 3172
rect 3767 3118 3823 3120
rect 3848 3172 3904 3174
rect 3848 3120 3850 3172
rect 3850 3120 3902 3172
rect 3902 3120 3904 3172
rect 3848 3118 3904 3120
rect 3929 3172 3985 3174
rect 3929 3120 3931 3172
rect 3931 3120 3983 3172
rect 3983 3120 3985 3172
rect 3929 3118 3985 3120
rect 4010 3172 4066 3174
rect 4010 3120 4012 3172
rect 4012 3120 4064 3172
rect 4064 3120 4066 3172
rect 4010 3118 4066 3120
rect 4091 3172 4147 3174
rect 4091 3120 4093 3172
rect 4093 3120 4145 3172
rect 4145 3120 4147 3172
rect 4091 3118 4147 3120
rect 4172 3172 4228 3174
rect 4172 3120 4174 3172
rect 4174 3120 4226 3172
rect 4226 3120 4228 3172
rect 4172 3118 4228 3120
rect 4254 3172 4310 3174
rect 4254 3120 4256 3172
rect 4256 3120 4308 3172
rect 4308 3120 4310 3172
rect 4254 3118 4310 3120
rect 4335 3172 4391 3174
rect 4335 3120 4337 3172
rect 4337 3120 4389 3172
rect 4389 3120 4391 3172
rect 4335 3118 4391 3120
rect 4416 3172 4472 3174
rect 4416 3120 4418 3172
rect 4418 3120 4470 3172
rect 4470 3120 4472 3172
rect 4416 3118 4472 3120
rect 4497 3172 4553 3174
rect 4497 3120 4499 3172
rect 4499 3120 4551 3172
rect 4551 3120 4553 3172
rect 4497 3118 4553 3120
rect 4578 3172 4634 3174
rect 4578 3120 4580 3172
rect 4580 3120 4632 3172
rect 4632 3120 4634 3172
rect 4578 3118 4634 3120
rect 4659 3172 4715 3174
rect 4659 3120 4661 3172
rect 4661 3120 4713 3172
rect 4713 3120 4715 3172
rect 4659 3118 4715 3120
rect 4740 3172 4796 3174
rect 4740 3120 4742 3172
rect 4742 3120 4794 3172
rect 4794 3120 4796 3172
rect 4740 3118 4796 3120
rect 4822 3172 4878 3174
rect 4822 3120 4824 3172
rect 4824 3120 4876 3172
rect 4876 3120 4878 3172
rect 4822 3118 4878 3120
rect 4903 3172 4959 3174
rect 4903 3120 4905 3172
rect 4905 3120 4957 3172
rect 4957 3120 4959 3172
rect 4903 3118 4959 3120
rect 4984 3172 5040 3174
rect 4984 3120 4986 3172
rect 4986 3120 5038 3172
rect 5038 3120 5040 3172
rect 4984 3118 5040 3120
rect 5065 3172 5121 3174
rect 5065 3120 5067 3172
rect 5067 3120 5119 3172
rect 5119 3120 5121 3172
rect 5065 3118 5121 3120
rect 5146 3172 5202 3174
rect 5146 3120 5148 3172
rect 5148 3120 5200 3172
rect 5200 3120 5202 3172
rect 5146 3118 5202 3120
rect 5227 3172 5283 3174
rect 5227 3120 5229 3172
rect 5229 3120 5281 3172
rect 5281 3120 5283 3172
rect 5227 3118 5283 3120
rect 5308 3172 5364 3174
rect 5308 3120 5310 3172
rect 5310 3120 5362 3172
rect 5362 3120 5364 3172
rect 5308 3118 5364 3120
rect 5390 3172 5446 3174
rect 5390 3120 5392 3172
rect 5392 3120 5444 3172
rect 5444 3120 5446 3172
rect 5390 3118 5446 3120
rect 5471 3172 5527 3174
rect 5471 3120 5473 3172
rect 5473 3120 5525 3172
rect 5525 3120 5527 3172
rect 5471 3118 5527 3120
rect 5552 3172 5608 3174
rect 5552 3120 5554 3172
rect 5554 3120 5606 3172
rect 5606 3120 5608 3172
rect 5552 3118 5608 3120
rect 5633 3172 5689 3174
rect 5633 3120 5635 3172
rect 5635 3120 5687 3172
rect 5687 3120 5689 3172
rect 5633 3118 5689 3120
rect 5714 3172 5770 3174
rect 5714 3120 5716 3172
rect 5716 3120 5768 3172
rect 5768 3120 5770 3172
rect 5714 3118 5770 3120
rect 5795 3172 5851 3174
rect 5795 3120 5797 3172
rect 5797 3120 5849 3172
rect 5849 3120 5851 3172
rect 5795 3118 5851 3120
rect 5876 3172 5932 3174
rect 5876 3120 5878 3172
rect 5878 3120 5930 3172
rect 5930 3120 5932 3172
rect 5876 3118 5932 3120
rect 5958 3172 6014 3174
rect 5958 3120 5960 3172
rect 5960 3120 6012 3172
rect 6012 3120 6014 3172
rect 5958 3118 6014 3120
rect 6039 3172 6095 3174
rect 6039 3120 6041 3172
rect 6041 3120 6093 3172
rect 6093 3120 6095 3172
rect 6039 3118 6095 3120
rect 6120 3172 6176 3174
rect 6120 3120 6122 3172
rect 6122 3120 6174 3172
rect 6174 3120 6176 3172
rect 6120 3118 6176 3120
rect 6201 3172 6257 3174
rect 6201 3120 6203 3172
rect 6203 3120 6255 3172
rect 6255 3120 6257 3172
rect 6201 3118 6257 3120
rect 6282 3172 6338 3174
rect 6282 3120 6284 3172
rect 6284 3120 6336 3172
rect 6336 3120 6338 3172
rect 6282 3118 6338 3120
rect 6363 3172 6419 3174
rect 6363 3120 6365 3172
rect 6365 3120 6417 3172
rect 6417 3120 6419 3172
rect 6363 3118 6419 3120
rect 6444 3172 6500 3174
rect 6444 3120 6446 3172
rect 6446 3120 6498 3172
rect 6498 3120 6500 3172
rect 6444 3118 6500 3120
rect 6526 3172 6582 3174
rect 6526 3120 6528 3172
rect 6528 3120 6580 3172
rect 6580 3120 6582 3172
rect 6526 3118 6582 3120
rect 6607 3172 6663 3174
rect 6607 3120 6609 3172
rect 6609 3120 6661 3172
rect 6661 3120 6663 3172
rect 6607 3118 6663 3120
rect 6688 3172 6744 3174
rect 6688 3120 6690 3172
rect 6690 3120 6742 3172
rect 6742 3120 6744 3172
rect 6688 3118 6744 3120
rect 6769 3172 6825 3174
rect 6769 3120 6771 3172
rect 6771 3120 6823 3172
rect 6823 3120 6825 3172
rect 6769 3118 6825 3120
rect 6850 3172 6906 3174
rect 6850 3120 6852 3172
rect 6852 3120 6904 3172
rect 6904 3120 6906 3172
rect 6850 3118 6906 3120
rect 6931 3172 6987 3174
rect 6931 3120 6933 3172
rect 6933 3120 6985 3172
rect 6985 3120 6987 3172
rect 6931 3118 6987 3120
rect 7012 3172 7068 3174
rect 7012 3120 7014 3172
rect 7014 3120 7066 3172
rect 7066 3120 7068 3172
rect 7012 3118 7068 3120
rect 7094 3172 7150 3174
rect 7094 3120 7096 3172
rect 7096 3120 7148 3172
rect 7148 3120 7150 3172
rect 7094 3118 7150 3120
rect 7175 3172 7231 3174
rect 7175 3120 7177 3172
rect 7177 3120 7229 3172
rect 7229 3120 7231 3172
rect 7175 3118 7231 3120
rect 7256 3172 7312 3174
rect 7256 3120 7258 3172
rect 7258 3120 7310 3172
rect 7310 3120 7312 3172
rect 7256 3118 7312 3120
rect 7337 3172 7393 3174
rect 7337 3120 7339 3172
rect 7339 3120 7391 3172
rect 7391 3120 7393 3172
rect 7337 3118 7393 3120
rect 7418 3172 7474 3174
rect 7418 3120 7420 3172
rect 7420 3120 7472 3172
rect 7472 3120 7474 3172
rect 7418 3118 7474 3120
rect 7499 3172 7555 3174
rect 7499 3120 7501 3172
rect 7501 3120 7553 3172
rect 7553 3120 7555 3172
rect 7499 3118 7555 3120
rect 7580 3172 7636 3174
rect 7580 3120 7582 3172
rect 7582 3120 7634 3172
rect 7634 3120 7636 3172
rect 7580 3118 7636 3120
rect 7662 3172 7718 3174
rect 7662 3120 7664 3172
rect 7664 3120 7716 3172
rect 7716 3120 7718 3172
rect 7662 3118 7718 3120
rect 7743 3172 7799 3174
rect 7743 3120 7745 3172
rect 7745 3120 7797 3172
rect 7797 3120 7799 3172
rect 7743 3118 7799 3120
rect 7824 3172 7880 3174
rect 7824 3120 7826 3172
rect 7826 3120 7878 3172
rect 7878 3120 7880 3172
rect 7824 3118 7880 3120
rect 7905 3172 7961 3174
rect 7905 3120 7907 3172
rect 7907 3120 7959 3172
rect 7959 3120 7961 3172
rect 7905 3118 7961 3120
rect 7986 3172 8042 3174
rect 7986 3120 7988 3172
rect 7988 3120 8040 3172
rect 8040 3120 8042 3172
rect 7986 3118 8042 3120
rect 8067 3172 8123 3174
rect 8067 3120 8069 3172
rect 8069 3120 8121 3172
rect 8121 3120 8123 3172
rect 8067 3118 8123 3120
rect 8148 3172 8204 3174
rect 8148 3120 8150 3172
rect 8150 3120 8202 3172
rect 8202 3120 8204 3172
rect 8148 3118 8204 3120
rect 8230 3172 8286 3174
rect 8230 3120 8232 3172
rect 8232 3120 8284 3172
rect 8284 3120 8286 3172
rect 8230 3118 8286 3120
rect 8311 3172 8367 3174
rect 8311 3120 8313 3172
rect 8313 3120 8365 3172
rect 8365 3120 8367 3172
rect 8311 3118 8367 3120
rect 8392 3172 8448 3174
rect 8392 3120 8394 3172
rect 8394 3120 8446 3172
rect 8446 3120 8448 3172
rect 8392 3118 8448 3120
rect 8473 3172 8529 3174
rect 8473 3120 8475 3172
rect 8475 3120 8527 3172
rect 8527 3120 8529 3172
rect 8473 3118 8529 3120
rect 8554 3172 8610 3174
rect 8554 3120 8556 3172
rect 8556 3120 8608 3172
rect 8608 3120 8610 3172
rect 8554 3118 8610 3120
rect 8635 3172 8691 3174
rect 8635 3120 8637 3172
rect 8637 3120 8689 3172
rect 8689 3120 8691 3172
rect 8635 3118 8691 3120
rect 8716 3172 8772 3174
rect 8716 3120 8718 3172
rect 8718 3120 8770 3172
rect 8770 3120 8772 3172
rect 8716 3118 8772 3120
rect 8798 3172 8854 3174
rect 8798 3120 8800 3172
rect 8800 3120 8852 3172
rect 8852 3120 8854 3172
rect 8798 3118 8854 3120
rect 8879 3172 8935 3174
rect 8879 3120 8881 3172
rect 8881 3120 8933 3172
rect 8933 3120 8935 3172
rect 8879 3118 8935 3120
rect 8960 3172 9016 3174
rect 8960 3120 8962 3172
rect 8962 3120 9014 3172
rect 9014 3120 9016 3172
rect 8960 3118 9016 3120
rect 9041 3172 9097 3174
rect 9041 3120 9043 3172
rect 9043 3120 9095 3172
rect 9095 3120 9097 3172
rect 9041 3118 9097 3120
rect 9122 3172 9178 3174
rect 9122 3120 9124 3172
rect 9124 3120 9176 3172
rect 9176 3120 9178 3172
rect 9122 3118 9178 3120
rect 9203 3172 9259 3174
rect 9203 3120 9205 3172
rect 9205 3120 9257 3172
rect 9257 3120 9259 3172
rect 9203 3118 9259 3120
rect 9284 3172 9340 3174
rect 9284 3120 9286 3172
rect 9286 3120 9338 3172
rect 9338 3120 9340 3172
rect 9284 3118 9340 3120
rect 9366 3172 9422 3174
rect 9366 3120 9368 3172
rect 9368 3120 9420 3172
rect 9420 3120 9422 3172
rect 9366 3118 9422 3120
rect 9447 3172 9503 3174
rect 9447 3120 9449 3172
rect 9449 3120 9501 3172
rect 9501 3120 9503 3172
rect 9447 3118 9503 3120
rect 9528 3172 9584 3174
rect 9528 3120 9530 3172
rect 9530 3120 9582 3172
rect 9582 3120 9584 3172
rect 9528 3118 9584 3120
rect 9609 3172 9665 3174
rect 9609 3120 9611 3172
rect 9611 3120 9663 3172
rect 9663 3120 9665 3172
rect 9609 3118 9665 3120
rect 9690 3172 9746 3174
rect 9690 3120 9692 3172
rect 9692 3120 9744 3172
rect 9744 3120 9746 3172
rect 9690 3118 9746 3120
rect 9771 3172 9827 3174
rect 9771 3120 9773 3172
rect 9773 3120 9825 3172
rect 9825 3120 9827 3172
rect 9771 3118 9827 3120
rect 9852 3172 9908 3174
rect 9852 3120 9854 3172
rect 9854 3120 9906 3172
rect 9906 3120 9908 3172
rect 9852 3118 9908 3120
rect 9934 3172 9990 3174
rect 9934 3120 9936 3172
rect 9936 3120 9988 3172
rect 9988 3120 9990 3172
rect 9934 3118 9990 3120
rect 10015 3172 10071 3174
rect 10015 3120 10017 3172
rect 10017 3120 10069 3172
rect 10069 3120 10071 3172
rect 10015 3118 10071 3120
rect 10096 3172 10152 3174
rect 10096 3120 10098 3172
rect 10098 3120 10150 3172
rect 10150 3120 10152 3172
rect 10096 3118 10152 3120
rect 10177 3172 10233 3174
rect 10177 3120 10179 3172
rect 10179 3120 10231 3172
rect 10231 3120 10233 3172
rect 10177 3118 10233 3120
rect 10258 3172 10314 3174
rect 10258 3120 10260 3172
rect 10260 3120 10312 3172
rect 10312 3120 10314 3172
rect 10258 3118 10314 3120
rect 10339 3172 10395 3174
rect 10339 3120 10341 3172
rect 10341 3120 10393 3172
rect 10393 3120 10395 3172
rect 10339 3118 10395 3120
rect 10420 3172 10476 3174
rect 10420 3120 10422 3172
rect 10422 3120 10474 3172
rect 10474 3120 10476 3172
rect 10420 3118 10476 3120
rect 10502 3172 10558 3174
rect 10502 3120 10504 3172
rect 10504 3120 10556 3172
rect 10556 3120 10558 3172
rect 10502 3118 10558 3120
rect 10583 3172 10639 3174
rect 10583 3120 10585 3172
rect 10585 3120 10637 3172
rect 10637 3120 10639 3172
rect 10583 3118 10639 3120
rect 10664 3172 10720 3174
rect 10664 3120 10666 3172
rect 10666 3120 10718 3172
rect 10718 3120 10720 3172
rect 10664 3118 10720 3120
rect 10745 3172 10801 3174
rect 10745 3120 10747 3172
rect 10747 3120 10799 3172
rect 10799 3120 10801 3172
rect 10745 3118 10801 3120
rect 10826 3172 10882 3174
rect 10826 3120 10828 3172
rect 10828 3120 10880 3172
rect 10880 3120 10882 3172
rect 10826 3118 10882 3120
rect 10907 3172 10963 3174
rect 10907 3120 10909 3172
rect 10909 3120 10961 3172
rect 10961 3120 10963 3172
rect 10907 3118 10963 3120
rect 10988 3172 11044 3174
rect 10988 3120 10990 3172
rect 10990 3120 11042 3172
rect 11042 3120 11044 3172
rect 10988 3118 11044 3120
rect 11116 3172 11172 3174
rect 11116 3120 11118 3172
rect 11118 3120 11170 3172
rect 11170 3120 11172 3172
rect 11116 3118 11172 3120
rect 11197 3172 11253 3174
rect 11197 3120 11199 3172
rect 11199 3120 11251 3172
rect 11251 3120 11253 3172
rect 11197 3118 11253 3120
rect 11278 3172 11334 3174
rect 11278 3120 11280 3172
rect 11280 3120 11332 3172
rect 11332 3120 11334 3172
rect 11278 3118 11334 3120
rect 11359 3172 11415 3174
rect 11359 3120 11361 3172
rect 11361 3120 11413 3172
rect 11413 3120 11415 3172
rect 11359 3118 11415 3120
rect 11440 3172 11496 3174
rect 11440 3120 11442 3172
rect 11442 3120 11494 3172
rect 11494 3120 11496 3172
rect 11440 3118 11496 3120
rect 11521 3172 11577 3174
rect 11521 3120 11523 3172
rect 11523 3120 11575 3172
rect 11575 3120 11577 3172
rect 11521 3118 11577 3120
rect 11602 3172 11658 3174
rect 11602 3120 11604 3172
rect 11604 3120 11656 3172
rect 11656 3120 11658 3172
rect 11602 3118 11658 3120
rect 11684 3172 11740 3174
rect 11684 3120 11686 3172
rect 11686 3120 11738 3172
rect 11738 3120 11740 3172
rect 11684 3118 11740 3120
rect 11765 3172 11821 3174
rect 11765 3120 11767 3172
rect 11767 3120 11819 3172
rect 11819 3120 11821 3172
rect 11765 3118 11821 3120
rect 11846 3172 11902 3174
rect 11846 3120 11848 3172
rect 11848 3120 11900 3172
rect 11900 3120 11902 3172
rect 11846 3118 11902 3120
rect 11927 3172 11983 3174
rect 11927 3120 11929 3172
rect 11929 3120 11981 3172
rect 11981 3120 11983 3172
rect 11927 3118 11983 3120
rect 12008 3172 12064 3174
rect 12008 3120 12010 3172
rect 12010 3120 12062 3172
rect 12062 3120 12064 3172
rect 12008 3118 12064 3120
rect 12089 3172 12145 3174
rect 12089 3120 12091 3172
rect 12091 3120 12143 3172
rect 12143 3120 12145 3172
rect 12089 3118 12145 3120
rect 12170 3172 12226 3174
rect 12170 3120 12172 3172
rect 12172 3120 12224 3172
rect 12224 3120 12226 3172
rect 12170 3118 12226 3120
rect 12252 3172 12308 3174
rect 12252 3120 12254 3172
rect 12254 3120 12306 3172
rect 12306 3120 12308 3172
rect 12252 3118 12308 3120
rect 12333 3172 12389 3174
rect 12333 3120 12335 3172
rect 12335 3120 12387 3172
rect 12387 3120 12389 3172
rect 12333 3118 12389 3120
rect 12414 3172 12470 3174
rect 12414 3120 12416 3172
rect 12416 3120 12468 3172
rect 12468 3120 12470 3172
rect 12414 3118 12470 3120
rect 12495 3172 12551 3174
rect 12495 3120 12497 3172
rect 12497 3120 12549 3172
rect 12549 3120 12551 3172
rect 12495 3118 12551 3120
rect 12576 3172 12632 3174
rect 12576 3120 12578 3172
rect 12578 3120 12630 3172
rect 12630 3120 12632 3172
rect 12576 3118 12632 3120
rect 12657 3172 12713 3174
rect 12657 3120 12659 3172
rect 12659 3120 12711 3172
rect 12711 3120 12713 3172
rect 12657 3118 12713 3120
rect 12738 3172 12794 3174
rect 12738 3120 12740 3172
rect 12740 3120 12792 3172
rect 12792 3120 12794 3172
rect 12738 3118 12794 3120
rect 12820 3172 12876 3174
rect 12820 3120 12822 3172
rect 12822 3120 12874 3172
rect 12874 3120 12876 3172
rect 12820 3118 12876 3120
rect 12901 3172 12957 3174
rect 12901 3120 12903 3172
rect 12903 3120 12955 3172
rect 12955 3120 12957 3172
rect 12901 3118 12957 3120
rect 12982 3172 13038 3174
rect 12982 3120 12984 3172
rect 12984 3120 13036 3172
rect 13036 3120 13038 3172
rect 12982 3118 13038 3120
rect 13063 3172 13119 3174
rect 13063 3120 13065 3172
rect 13065 3120 13117 3172
rect 13117 3120 13119 3172
rect 13063 3118 13119 3120
rect 13144 3172 13200 3174
rect 13144 3120 13146 3172
rect 13146 3120 13198 3172
rect 13198 3120 13200 3172
rect 13144 3118 13200 3120
rect 13225 3172 13281 3174
rect 13225 3120 13227 3172
rect 13227 3120 13279 3172
rect 13279 3120 13281 3172
rect 13225 3118 13281 3120
rect 13306 3172 13362 3174
rect 13306 3120 13308 3172
rect 13308 3120 13360 3172
rect 13360 3120 13362 3172
rect 13306 3118 13362 3120
rect 13388 3172 13444 3174
rect 13388 3120 13390 3172
rect 13390 3120 13442 3172
rect 13442 3120 13444 3172
rect 13388 3118 13444 3120
rect 13469 3172 13525 3174
rect 13469 3120 13471 3172
rect 13471 3120 13523 3172
rect 13523 3120 13525 3172
rect 13469 3118 13525 3120
rect 13550 3172 13606 3174
rect 13550 3120 13552 3172
rect 13552 3120 13604 3172
rect 13604 3120 13606 3172
rect 13550 3118 13606 3120
rect 13631 3172 13687 3174
rect 13631 3120 13633 3172
rect 13633 3120 13685 3172
rect 13685 3120 13687 3172
rect 13631 3118 13687 3120
rect 13712 3172 13768 3174
rect 13712 3120 13714 3172
rect 13714 3120 13766 3172
rect 13766 3120 13768 3172
rect 13712 3118 13768 3120
rect 13793 3172 13849 3174
rect 13793 3120 13795 3172
rect 13795 3120 13847 3172
rect 13847 3120 13849 3172
rect 13793 3118 13849 3120
rect 13874 3172 13930 3174
rect 13874 3120 13876 3172
rect 13876 3120 13928 3172
rect 13928 3120 13930 3172
rect 13874 3118 13930 3120
rect 13956 3172 14012 3174
rect 13956 3120 13958 3172
rect 13958 3120 14010 3172
rect 14010 3120 14012 3172
rect 13956 3118 14012 3120
rect 14037 3172 14093 3174
rect 14037 3120 14039 3172
rect 14039 3120 14091 3172
rect 14091 3120 14093 3172
rect 14037 3118 14093 3120
rect 14118 3172 14174 3174
rect 14118 3120 14120 3172
rect 14120 3120 14172 3172
rect 14172 3120 14174 3172
rect 14118 3118 14174 3120
rect 14199 3172 14255 3174
rect 14199 3120 14201 3172
rect 14201 3120 14253 3172
rect 14253 3120 14255 3172
rect 14199 3118 14255 3120
rect 14280 3172 14336 3174
rect 14280 3120 14282 3172
rect 14282 3120 14334 3172
rect 14334 3120 14336 3172
rect 14280 3118 14336 3120
rect 14361 3172 14417 3174
rect 14361 3120 14363 3172
rect 14363 3120 14415 3172
rect 14415 3120 14417 3172
rect 14361 3118 14417 3120
rect 14442 3172 14498 3174
rect 14442 3120 14444 3172
rect 14444 3120 14496 3172
rect 14496 3120 14498 3172
rect 14442 3118 14498 3120
rect 14524 3172 14580 3174
rect 14524 3120 14526 3172
rect 14526 3120 14578 3172
rect 14578 3120 14580 3172
rect 14524 3118 14580 3120
rect 14605 3172 14661 3174
rect 14605 3120 14607 3172
rect 14607 3120 14659 3172
rect 14659 3120 14661 3172
rect 14605 3118 14661 3120
rect 14686 3172 14742 3174
rect 14686 3120 14688 3172
rect 14688 3120 14740 3172
rect 14740 3120 14742 3172
rect 14686 3118 14742 3120
rect 14767 3172 14823 3174
rect 14767 3120 14769 3172
rect 14769 3120 14821 3172
rect 14821 3120 14823 3172
rect 14767 3118 14823 3120
rect 14848 3172 14904 3174
rect 14848 3120 14850 3172
rect 14850 3120 14902 3172
rect 14902 3120 14904 3172
rect 14848 3118 14904 3120
rect 14929 3172 14985 3174
rect 14929 3120 14931 3172
rect 14931 3120 14983 3172
rect 14983 3120 14985 3172
rect 14929 3118 14985 3120
rect 15010 3172 15066 3174
rect 15010 3120 15012 3172
rect 15012 3120 15064 3172
rect 15064 3120 15066 3172
rect 15010 3118 15066 3120
rect 15092 3172 15148 3174
rect 15092 3120 15094 3172
rect 15094 3120 15146 3172
rect 15146 3120 15148 3172
rect 15092 3118 15148 3120
rect 15173 3172 15229 3174
rect 15173 3120 15175 3172
rect 15175 3120 15227 3172
rect 15227 3120 15229 3172
rect 15173 3118 15229 3120
rect 15254 3172 15310 3174
rect 15254 3120 15256 3172
rect 15256 3120 15308 3172
rect 15308 3120 15310 3172
rect 15254 3118 15310 3120
rect 15335 3172 15391 3174
rect 15335 3120 15337 3172
rect 15337 3120 15389 3172
rect 15389 3120 15391 3172
rect 15335 3118 15391 3120
rect 15416 3172 15472 3174
rect 15416 3120 15418 3172
rect 15418 3120 15470 3172
rect 15470 3120 15472 3172
rect 15416 3118 15472 3120
rect 15497 3172 15553 3174
rect 15497 3120 15499 3172
rect 15499 3120 15551 3172
rect 15551 3120 15553 3172
rect 15497 3118 15553 3120
rect 15578 3172 15634 3174
rect 15578 3120 15580 3172
rect 15580 3120 15632 3172
rect 15632 3120 15634 3172
rect 15578 3118 15634 3120
rect 15660 3172 15716 3174
rect 15660 3120 15662 3172
rect 15662 3120 15714 3172
rect 15714 3120 15716 3172
rect 15660 3118 15716 3120
rect 15741 3172 15797 3174
rect 15741 3120 15743 3172
rect 15743 3120 15795 3172
rect 15795 3120 15797 3172
rect 15741 3118 15797 3120
rect 15822 3172 15878 3174
rect 15822 3120 15824 3172
rect 15824 3120 15876 3172
rect 15876 3120 15878 3172
rect 15822 3118 15878 3120
rect 15903 3172 15959 3174
rect 15903 3120 15905 3172
rect 15905 3120 15957 3172
rect 15957 3120 15959 3172
rect 15903 3118 15959 3120
rect 15984 3172 16040 3174
rect 15984 3120 15986 3172
rect 15986 3120 16038 3172
rect 16038 3120 16040 3172
rect 15984 3118 16040 3120
rect 16065 3172 16121 3174
rect 16065 3120 16067 3172
rect 16067 3120 16119 3172
rect 16119 3120 16121 3172
rect 16065 3118 16121 3120
rect 16146 3172 16202 3174
rect 16146 3120 16148 3172
rect 16148 3120 16200 3172
rect 16200 3120 16202 3172
rect 16146 3118 16202 3120
rect 16228 3172 16284 3174
rect 16228 3120 16230 3172
rect 16230 3120 16282 3172
rect 16282 3120 16284 3172
rect 16228 3118 16284 3120
rect 16309 3172 16365 3174
rect 16309 3120 16311 3172
rect 16311 3120 16363 3172
rect 16363 3120 16365 3172
rect 16309 3118 16365 3120
rect 16390 3172 16446 3174
rect 16390 3120 16392 3172
rect 16392 3120 16444 3172
rect 16444 3120 16446 3172
rect 16390 3118 16446 3120
rect 16471 3172 16527 3174
rect 16471 3120 16473 3172
rect 16473 3120 16525 3172
rect 16525 3120 16527 3172
rect 16471 3118 16527 3120
rect 16552 3172 16608 3174
rect 16552 3120 16554 3172
rect 16554 3120 16606 3172
rect 16606 3120 16608 3172
rect 16552 3118 16608 3120
rect 16633 3172 16689 3174
rect 16633 3120 16635 3172
rect 16635 3120 16687 3172
rect 16687 3120 16689 3172
rect 16633 3118 16689 3120
rect 16714 3172 16770 3174
rect 16714 3120 16716 3172
rect 16716 3120 16768 3172
rect 16768 3120 16770 3172
rect 16714 3118 16770 3120
rect 16796 3172 16852 3174
rect 16796 3120 16798 3172
rect 16798 3120 16850 3172
rect 16850 3120 16852 3172
rect 16796 3118 16852 3120
rect 16877 3172 16933 3174
rect 16877 3120 16879 3172
rect 16879 3120 16931 3172
rect 16931 3120 16933 3172
rect 16877 3118 16933 3120
rect 16958 3172 17014 3174
rect 16958 3120 16960 3172
rect 16960 3120 17012 3172
rect 17012 3120 17014 3172
rect 16958 3118 17014 3120
rect 17039 3172 17095 3174
rect 17039 3120 17041 3172
rect 17041 3120 17093 3172
rect 17093 3120 17095 3172
rect 17039 3118 17095 3120
rect 17120 3172 17176 3174
rect 17120 3120 17122 3172
rect 17122 3120 17174 3172
rect 17174 3120 17176 3172
rect 17120 3118 17176 3120
rect 17201 3172 17257 3174
rect 17201 3120 17203 3172
rect 17203 3120 17255 3172
rect 17255 3120 17257 3172
rect 17201 3118 17257 3120
rect 17282 3172 17338 3174
rect 17282 3120 17284 3172
rect 17284 3120 17336 3172
rect 17336 3120 17338 3172
rect 17282 3118 17338 3120
rect 17364 3172 17420 3174
rect 17364 3120 17366 3172
rect 17366 3120 17418 3172
rect 17418 3120 17420 3172
rect 17364 3118 17420 3120
rect 17445 3172 17501 3174
rect 17445 3120 17447 3172
rect 17447 3120 17499 3172
rect 17499 3120 17501 3172
rect 17445 3118 17501 3120
rect 17526 3172 17582 3174
rect 17526 3120 17528 3172
rect 17528 3120 17580 3172
rect 17580 3120 17582 3172
rect 17526 3118 17582 3120
rect 17607 3172 17663 3174
rect 17607 3120 17609 3172
rect 17609 3120 17661 3172
rect 17661 3120 17663 3172
rect 17607 3118 17663 3120
rect 17688 3172 17744 3174
rect 17688 3120 17690 3172
rect 17690 3120 17742 3172
rect 17742 3120 17744 3172
rect 17688 3118 17744 3120
rect 17769 3172 17825 3174
rect 17769 3120 17771 3172
rect 17771 3120 17823 3172
rect 17823 3120 17825 3172
rect 17769 3118 17825 3120
rect 17850 3172 17906 3174
rect 17850 3120 17852 3172
rect 17852 3120 17904 3172
rect 17904 3120 17906 3172
rect 17850 3118 17906 3120
rect 17932 3172 17988 3174
rect 17932 3120 17934 3172
rect 17934 3120 17986 3172
rect 17986 3120 17988 3172
rect 17932 3118 17988 3120
rect 18013 3172 18069 3174
rect 18013 3120 18015 3172
rect 18015 3120 18067 3172
rect 18067 3120 18069 3172
rect 18013 3118 18069 3120
rect 18094 3172 18150 3174
rect 18094 3120 18096 3172
rect 18096 3120 18148 3172
rect 18148 3120 18150 3172
rect 18094 3118 18150 3120
rect 18175 3172 18231 3174
rect 18175 3120 18177 3172
rect 18177 3120 18229 3172
rect 18229 3120 18231 3172
rect 18175 3118 18231 3120
rect 18256 3172 18312 3174
rect 18256 3120 18258 3172
rect 18258 3120 18310 3172
rect 18310 3120 18312 3172
rect 18256 3118 18312 3120
rect 18337 3172 18393 3174
rect 18337 3120 18339 3172
rect 18339 3120 18391 3172
rect 18391 3120 18393 3172
rect 18337 3118 18393 3120
rect 18418 3172 18474 3174
rect 18418 3120 18420 3172
rect 18420 3120 18472 3172
rect 18472 3120 18474 3172
rect 18418 3118 18474 3120
rect 18500 3172 18556 3174
rect 18500 3120 18502 3172
rect 18502 3120 18554 3172
rect 18554 3120 18556 3172
rect 18500 3118 18556 3120
rect 18581 3172 18637 3174
rect 18581 3120 18583 3172
rect 18583 3120 18635 3172
rect 18635 3120 18637 3172
rect 18581 3118 18637 3120
rect 18662 3172 18718 3174
rect 18662 3120 18664 3172
rect 18664 3120 18716 3172
rect 18716 3120 18718 3172
rect 18662 3118 18718 3120
rect 18743 3172 18799 3174
rect 18743 3120 18745 3172
rect 18745 3120 18797 3172
rect 18797 3120 18799 3172
rect 18743 3118 18799 3120
rect 18824 3172 18880 3174
rect 18824 3120 18826 3172
rect 18826 3120 18878 3172
rect 18878 3120 18880 3172
rect 18824 3118 18880 3120
rect 18905 3172 18961 3174
rect 18905 3120 18907 3172
rect 18907 3120 18959 3172
rect 18959 3120 18961 3172
rect 18905 3118 18961 3120
rect 18986 3172 19042 3174
rect 18986 3120 18988 3172
rect 18988 3120 19040 3172
rect 19040 3120 19042 3172
rect 18986 3118 19042 3120
rect 19068 3172 19124 3174
rect 19068 3120 19070 3172
rect 19070 3120 19122 3172
rect 19122 3120 19124 3172
rect 19068 3118 19124 3120
rect 19149 3172 19205 3174
rect 19149 3120 19151 3172
rect 19151 3120 19203 3172
rect 19203 3120 19205 3172
rect 19149 3118 19205 3120
rect 19230 3172 19286 3174
rect 19230 3120 19232 3172
rect 19232 3120 19284 3172
rect 19284 3120 19286 3172
rect 19230 3118 19286 3120
rect 19311 3172 19367 3174
rect 19311 3120 19313 3172
rect 19313 3120 19365 3172
rect 19365 3120 19367 3172
rect 19311 3118 19367 3120
rect 19392 3172 19448 3174
rect 19392 3120 19394 3172
rect 19394 3120 19446 3172
rect 19446 3120 19448 3172
rect 19392 3118 19448 3120
rect 19473 3172 19529 3174
rect 19473 3120 19475 3172
rect 19475 3120 19527 3172
rect 19527 3120 19529 3172
rect 19473 3118 19529 3120
rect 19554 3172 19610 3174
rect 19554 3120 19556 3172
rect 19556 3120 19608 3172
rect 19608 3120 19610 3172
rect 19554 3118 19610 3120
rect 19636 3172 19692 3174
rect 19636 3120 19638 3172
rect 19638 3120 19690 3172
rect 19690 3120 19692 3172
rect 19636 3118 19692 3120
rect 19717 3172 19773 3174
rect 19717 3120 19719 3172
rect 19719 3120 19771 3172
rect 19771 3120 19773 3172
rect 19717 3118 19773 3120
rect 19798 3172 19854 3174
rect 19798 3120 19800 3172
rect 19800 3120 19852 3172
rect 19852 3120 19854 3172
rect 19798 3118 19854 3120
rect 19879 3172 19935 3174
rect 19879 3120 19881 3172
rect 19881 3120 19933 3172
rect 19933 3120 19935 3172
rect 19879 3118 19935 3120
rect 19960 3172 20016 3174
rect 19960 3120 19962 3172
rect 19962 3120 20014 3172
rect 20014 3120 20016 3172
rect 19960 3118 20016 3120
rect 20041 3172 20097 3174
rect 20041 3120 20043 3172
rect 20043 3120 20095 3172
rect 20095 3120 20097 3172
rect 20041 3118 20097 3120
rect 20122 3172 20178 3174
rect 20122 3120 20124 3172
rect 20124 3120 20176 3172
rect 20176 3120 20178 3172
rect 20122 3118 20178 3120
rect 20204 3172 20260 3174
rect 20204 3120 20206 3172
rect 20206 3120 20258 3172
rect 20258 3120 20260 3172
rect 20204 3118 20260 3120
rect 20285 3172 20341 3174
rect 20285 3120 20287 3172
rect 20287 3120 20339 3172
rect 20339 3120 20341 3172
rect 20285 3118 20341 3120
rect 20366 3172 20422 3174
rect 20366 3120 20368 3172
rect 20368 3120 20420 3172
rect 20420 3120 20422 3172
rect 20366 3118 20422 3120
rect 20447 3172 20503 3174
rect 20447 3120 20449 3172
rect 20449 3120 20501 3172
rect 20501 3120 20503 3172
rect 20447 3118 20503 3120
rect 20528 3172 20584 3174
rect 20528 3120 20530 3172
rect 20530 3120 20582 3172
rect 20582 3120 20584 3172
rect 20528 3118 20584 3120
rect 20609 3172 20665 3174
rect 20609 3120 20611 3172
rect 20611 3120 20663 3172
rect 20663 3120 20665 3172
rect 20609 3118 20665 3120
rect 20690 3172 20746 3174
rect 20690 3120 20692 3172
rect 20692 3120 20744 3172
rect 20744 3120 20746 3172
rect 20690 3118 20746 3120
rect 20772 3172 20828 3174
rect 20772 3120 20774 3172
rect 20774 3120 20826 3172
rect 20826 3120 20828 3172
rect 20772 3118 20828 3120
rect 20853 3172 20909 3174
rect 20853 3120 20855 3172
rect 20855 3120 20907 3172
rect 20907 3120 20909 3172
rect 20853 3118 20909 3120
rect 20934 3172 20990 3174
rect 20934 3120 20936 3172
rect 20936 3120 20988 3172
rect 20988 3120 20990 3172
rect 20934 3118 20990 3120
rect 21015 3172 21071 3174
rect 21015 3120 21017 3172
rect 21017 3120 21069 3172
rect 21069 3120 21071 3172
rect 21015 3118 21071 3120
rect 21096 3172 21152 3174
rect 21096 3120 21098 3172
rect 21098 3120 21150 3172
rect 21150 3120 21152 3172
rect 21096 3118 21152 3120
rect 21177 3172 21233 3174
rect 21177 3120 21179 3172
rect 21179 3120 21231 3172
rect 21231 3120 21233 3172
rect 21177 3118 21233 3120
rect 21258 3172 21314 3174
rect 21258 3120 21260 3172
rect 21260 3120 21312 3172
rect 21312 3120 21314 3172
rect 21258 3118 21314 3120
rect 21340 3172 21396 3174
rect 21340 3120 21342 3172
rect 21342 3120 21394 3172
rect 21394 3120 21396 3172
rect 21340 3118 21396 3120
rect 21421 3172 21477 3174
rect 21421 3120 21423 3172
rect 21423 3120 21475 3172
rect 21475 3120 21477 3172
rect 21421 3118 21477 3120
rect 21502 3172 21558 3174
rect 21502 3120 21504 3172
rect 21504 3120 21556 3172
rect 21556 3120 21558 3172
rect 21502 3118 21558 3120
rect 21583 3172 21639 3174
rect 21583 3120 21585 3172
rect 21585 3120 21637 3172
rect 21637 3120 21639 3172
rect 21583 3118 21639 3120
rect 21664 3172 21720 3174
rect 21664 3120 21666 3172
rect 21666 3120 21718 3172
rect 21718 3120 21720 3172
rect 21664 3118 21720 3120
rect 21745 3172 21801 3174
rect 21745 3120 21747 3172
rect 21747 3120 21799 3172
rect 21799 3120 21801 3172
rect 21745 3118 21801 3120
rect 21826 3172 21882 3174
rect 21826 3120 21828 3172
rect 21828 3120 21880 3172
rect 21880 3120 21882 3172
rect 21826 3118 21882 3120
rect 21908 3172 21964 3174
rect 21908 3120 21910 3172
rect 21910 3120 21962 3172
rect 21962 3120 21964 3172
rect 21908 3118 21964 3120
rect 21989 3172 22045 3174
rect 21989 3120 21991 3172
rect 21991 3120 22043 3172
rect 22043 3120 22045 3172
rect 21989 3118 22045 3120
rect 22070 3172 22126 3174
rect 22070 3120 22072 3172
rect 22072 3120 22124 3172
rect 22124 3120 22126 3172
rect 22070 3118 22126 3120
rect 22151 3172 22207 3174
rect 22151 3120 22153 3172
rect 22153 3120 22205 3172
rect 22205 3120 22207 3172
rect 22151 3118 22207 3120
rect 22232 3172 22288 3174
rect 22232 3120 22234 3172
rect 22234 3120 22286 3172
rect 22286 3120 22288 3172
rect 22232 3118 22288 3120
rect 22313 3172 22369 3174
rect 22313 3120 22315 3172
rect 22315 3120 22367 3172
rect 22367 3120 22369 3172
rect 22313 3118 22369 3120
rect 22394 3172 22450 3174
rect 22394 3120 22396 3172
rect 22396 3120 22448 3172
rect 22448 3120 22450 3172
rect 22394 3118 22450 3120
rect 22476 3172 22532 3174
rect 22476 3120 22478 3172
rect 22478 3120 22530 3172
rect 22530 3120 22532 3172
rect 22476 3118 22532 3120
rect 22557 3172 22613 3174
rect 22557 3120 22559 3172
rect 22559 3120 22611 3172
rect 22611 3120 22613 3172
rect 22557 3118 22613 3120
rect 22638 3172 22694 3174
rect 22638 3120 22640 3172
rect 22640 3120 22692 3172
rect 22692 3120 22694 3172
rect 22638 3118 22694 3120
rect 22719 3172 22775 3174
rect 22719 3120 22721 3172
rect 22721 3120 22773 3172
rect 22773 3120 22775 3172
rect 22719 3118 22775 3120
rect 22800 3172 22856 3174
rect 22800 3120 22802 3172
rect 22802 3120 22854 3172
rect 22854 3120 22856 3172
rect 22800 3118 22856 3120
rect 22881 3172 22937 3174
rect 22881 3120 22883 3172
rect 22883 3120 22935 3172
rect 22935 3120 22937 3172
rect 22881 3118 22937 3120
rect 22962 3172 23018 3174
rect 22962 3120 22964 3172
rect 22964 3120 23016 3172
rect 23016 3120 23018 3172
rect 22962 3118 23018 3120
rect 23044 3172 23100 3174
rect 23044 3120 23046 3172
rect 23046 3120 23098 3172
rect 23098 3120 23100 3172
rect 23044 3118 23100 3120
rect 23125 3172 23181 3174
rect 23125 3120 23127 3172
rect 23127 3120 23179 3172
rect 23179 3120 23181 3172
rect 23125 3118 23181 3120
rect 23206 3172 23262 3174
rect 23206 3120 23208 3172
rect 23208 3120 23260 3172
rect 23260 3120 23262 3172
rect 23206 3118 23262 3120
rect 23287 3172 23343 3174
rect 23287 3120 23289 3172
rect 23289 3120 23341 3172
rect 23341 3120 23343 3172
rect 23287 3118 23343 3120
rect 23368 3172 23424 3174
rect 23368 3120 23370 3172
rect 23370 3120 23422 3172
rect 23422 3120 23424 3172
rect 23368 3118 23424 3120
rect 23449 3172 23505 3174
rect 23449 3120 23451 3172
rect 23451 3120 23503 3172
rect 23503 3120 23505 3172
rect 23449 3118 23505 3120
rect 23530 3172 23586 3174
rect 23530 3120 23532 3172
rect 23532 3120 23584 3172
rect 23584 3120 23586 3172
rect 23530 3118 23586 3120
rect 23612 3172 23668 3174
rect 23612 3120 23614 3172
rect 23614 3120 23666 3172
rect 23666 3120 23668 3172
rect 23612 3118 23668 3120
rect 23693 3172 23749 3174
rect 23693 3120 23695 3172
rect 23695 3120 23747 3172
rect 23747 3120 23749 3172
rect 23693 3118 23749 3120
rect 23774 3172 23830 3174
rect 23774 3120 23776 3172
rect 23776 3120 23828 3172
rect 23828 3120 23830 3172
rect 23774 3118 23830 3120
rect 23855 3172 23911 3174
rect 23855 3120 23857 3172
rect 23857 3120 23909 3172
rect 23909 3120 23911 3172
rect 23855 3118 23911 3120
rect 23936 3172 23992 3174
rect 23936 3120 23938 3172
rect 23938 3120 23990 3172
rect 23990 3120 23992 3172
rect 23936 3118 23992 3120
rect 24017 3172 24073 3174
rect 24017 3120 24019 3172
rect 24019 3120 24071 3172
rect 24071 3120 24073 3172
rect 24017 3118 24073 3120
rect 24098 3172 24154 3174
rect 24098 3120 24100 3172
rect 24100 3120 24152 3172
rect 24152 3120 24154 3172
rect 24098 3118 24154 3120
rect 24180 3172 24236 3174
rect 24180 3120 24182 3172
rect 24182 3120 24234 3172
rect 24234 3120 24236 3172
rect 24180 3118 24236 3120
rect 24261 3172 24317 3174
rect 24261 3120 24263 3172
rect 24263 3120 24315 3172
rect 24315 3120 24317 3172
rect 24261 3118 24317 3120
rect 24342 3172 24398 3174
rect 24342 3120 24344 3172
rect 24344 3120 24396 3172
rect 24396 3120 24398 3172
rect 24342 3118 24398 3120
rect 24423 3172 24479 3174
rect 24423 3120 24425 3172
rect 24425 3120 24477 3172
rect 24477 3120 24479 3172
rect 24423 3118 24479 3120
rect 24504 3172 24560 3174
rect 24504 3120 24506 3172
rect 24506 3120 24558 3172
rect 24558 3120 24560 3172
rect 24504 3118 24560 3120
rect 24585 3172 24641 3174
rect 24585 3120 24587 3172
rect 24587 3120 24639 3172
rect 24639 3120 24641 3172
rect 24585 3118 24641 3120
rect 24666 3172 24722 3174
rect 24666 3120 24668 3172
rect 24668 3120 24720 3172
rect 24720 3120 24722 3172
rect 24666 3118 24722 3120
rect 3036 3068 3092 3070
rect 3036 3016 3038 3068
rect 3038 3016 3090 3068
rect 3090 3016 3092 3068
rect 3036 3014 3092 3016
rect 3118 3068 3174 3070
rect 3118 3016 3120 3068
rect 3120 3016 3172 3068
rect 3172 3016 3174 3068
rect 3118 3014 3174 3016
rect 3199 3068 3255 3070
rect 3199 3016 3201 3068
rect 3201 3016 3253 3068
rect 3253 3016 3255 3068
rect 3199 3014 3255 3016
rect 3280 3068 3336 3070
rect 3280 3016 3282 3068
rect 3282 3016 3334 3068
rect 3334 3016 3336 3068
rect 3280 3014 3336 3016
rect 3361 3068 3417 3070
rect 3361 3016 3363 3068
rect 3363 3016 3415 3068
rect 3415 3016 3417 3068
rect 3361 3014 3417 3016
rect 3442 3068 3498 3070
rect 3442 3016 3444 3068
rect 3444 3016 3496 3068
rect 3496 3016 3498 3068
rect 3442 3014 3498 3016
rect 3523 3068 3579 3070
rect 3523 3016 3525 3068
rect 3525 3016 3577 3068
rect 3577 3016 3579 3068
rect 3523 3014 3579 3016
rect 3604 3068 3660 3070
rect 3604 3016 3606 3068
rect 3606 3016 3658 3068
rect 3658 3016 3660 3068
rect 3604 3014 3660 3016
rect 3686 3068 3742 3070
rect 3686 3016 3688 3068
rect 3688 3016 3740 3068
rect 3740 3016 3742 3068
rect 3686 3014 3742 3016
rect 3767 3068 3823 3070
rect 3767 3016 3769 3068
rect 3769 3016 3821 3068
rect 3821 3016 3823 3068
rect 3767 3014 3823 3016
rect 3848 3068 3904 3070
rect 3848 3016 3850 3068
rect 3850 3016 3902 3068
rect 3902 3016 3904 3068
rect 3848 3014 3904 3016
rect 3929 3068 3985 3070
rect 3929 3016 3931 3068
rect 3931 3016 3983 3068
rect 3983 3016 3985 3068
rect 3929 3014 3985 3016
rect 4010 3068 4066 3070
rect 4010 3016 4012 3068
rect 4012 3016 4064 3068
rect 4064 3016 4066 3068
rect 4010 3014 4066 3016
rect 4091 3068 4147 3070
rect 4091 3016 4093 3068
rect 4093 3016 4145 3068
rect 4145 3016 4147 3068
rect 4091 3014 4147 3016
rect 4172 3068 4228 3070
rect 4172 3016 4174 3068
rect 4174 3016 4226 3068
rect 4226 3016 4228 3068
rect 4172 3014 4228 3016
rect 4254 3068 4310 3070
rect 4254 3016 4256 3068
rect 4256 3016 4308 3068
rect 4308 3016 4310 3068
rect 4254 3014 4310 3016
rect 4335 3068 4391 3070
rect 4335 3016 4337 3068
rect 4337 3016 4389 3068
rect 4389 3016 4391 3068
rect 4335 3014 4391 3016
rect 4416 3068 4472 3070
rect 4416 3016 4418 3068
rect 4418 3016 4470 3068
rect 4470 3016 4472 3068
rect 4416 3014 4472 3016
rect 4497 3068 4553 3070
rect 4497 3016 4499 3068
rect 4499 3016 4551 3068
rect 4551 3016 4553 3068
rect 4497 3014 4553 3016
rect 4578 3068 4634 3070
rect 4578 3016 4580 3068
rect 4580 3016 4632 3068
rect 4632 3016 4634 3068
rect 4578 3014 4634 3016
rect 4659 3068 4715 3070
rect 4659 3016 4661 3068
rect 4661 3016 4713 3068
rect 4713 3016 4715 3068
rect 4659 3014 4715 3016
rect 4740 3068 4796 3070
rect 4740 3016 4742 3068
rect 4742 3016 4794 3068
rect 4794 3016 4796 3068
rect 4740 3014 4796 3016
rect 4822 3068 4878 3070
rect 4822 3016 4824 3068
rect 4824 3016 4876 3068
rect 4876 3016 4878 3068
rect 4822 3014 4878 3016
rect 4903 3068 4959 3070
rect 4903 3016 4905 3068
rect 4905 3016 4957 3068
rect 4957 3016 4959 3068
rect 4903 3014 4959 3016
rect 4984 3068 5040 3070
rect 4984 3016 4986 3068
rect 4986 3016 5038 3068
rect 5038 3016 5040 3068
rect 4984 3014 5040 3016
rect 5065 3068 5121 3070
rect 5065 3016 5067 3068
rect 5067 3016 5119 3068
rect 5119 3016 5121 3068
rect 5065 3014 5121 3016
rect 5146 3068 5202 3070
rect 5146 3016 5148 3068
rect 5148 3016 5200 3068
rect 5200 3016 5202 3068
rect 5146 3014 5202 3016
rect 5227 3068 5283 3070
rect 5227 3016 5229 3068
rect 5229 3016 5281 3068
rect 5281 3016 5283 3068
rect 5227 3014 5283 3016
rect 5308 3068 5364 3070
rect 5308 3016 5310 3068
rect 5310 3016 5362 3068
rect 5362 3016 5364 3068
rect 5308 3014 5364 3016
rect 5390 3068 5446 3070
rect 5390 3016 5392 3068
rect 5392 3016 5444 3068
rect 5444 3016 5446 3068
rect 5390 3014 5446 3016
rect 5471 3068 5527 3070
rect 5471 3016 5473 3068
rect 5473 3016 5525 3068
rect 5525 3016 5527 3068
rect 5471 3014 5527 3016
rect 5552 3068 5608 3070
rect 5552 3016 5554 3068
rect 5554 3016 5606 3068
rect 5606 3016 5608 3068
rect 5552 3014 5608 3016
rect 5633 3068 5689 3070
rect 5633 3016 5635 3068
rect 5635 3016 5687 3068
rect 5687 3016 5689 3068
rect 5633 3014 5689 3016
rect 5714 3068 5770 3070
rect 5714 3016 5716 3068
rect 5716 3016 5768 3068
rect 5768 3016 5770 3068
rect 5714 3014 5770 3016
rect 5795 3068 5851 3070
rect 5795 3016 5797 3068
rect 5797 3016 5849 3068
rect 5849 3016 5851 3068
rect 5795 3014 5851 3016
rect 5876 3068 5932 3070
rect 5876 3016 5878 3068
rect 5878 3016 5930 3068
rect 5930 3016 5932 3068
rect 5876 3014 5932 3016
rect 5958 3068 6014 3070
rect 5958 3016 5960 3068
rect 5960 3016 6012 3068
rect 6012 3016 6014 3068
rect 5958 3014 6014 3016
rect 6039 3068 6095 3070
rect 6039 3016 6041 3068
rect 6041 3016 6093 3068
rect 6093 3016 6095 3068
rect 6039 3014 6095 3016
rect 6120 3068 6176 3070
rect 6120 3016 6122 3068
rect 6122 3016 6174 3068
rect 6174 3016 6176 3068
rect 6120 3014 6176 3016
rect 6201 3068 6257 3070
rect 6201 3016 6203 3068
rect 6203 3016 6255 3068
rect 6255 3016 6257 3068
rect 6201 3014 6257 3016
rect 6282 3068 6338 3070
rect 6282 3016 6284 3068
rect 6284 3016 6336 3068
rect 6336 3016 6338 3068
rect 6282 3014 6338 3016
rect 6363 3068 6419 3070
rect 6363 3016 6365 3068
rect 6365 3016 6417 3068
rect 6417 3016 6419 3068
rect 6363 3014 6419 3016
rect 6444 3068 6500 3070
rect 6444 3016 6446 3068
rect 6446 3016 6498 3068
rect 6498 3016 6500 3068
rect 6444 3014 6500 3016
rect 6526 3068 6582 3070
rect 6526 3016 6528 3068
rect 6528 3016 6580 3068
rect 6580 3016 6582 3068
rect 6526 3014 6582 3016
rect 6607 3068 6663 3070
rect 6607 3016 6609 3068
rect 6609 3016 6661 3068
rect 6661 3016 6663 3068
rect 6607 3014 6663 3016
rect 6688 3068 6744 3070
rect 6688 3016 6690 3068
rect 6690 3016 6742 3068
rect 6742 3016 6744 3068
rect 6688 3014 6744 3016
rect 6769 3068 6825 3070
rect 6769 3016 6771 3068
rect 6771 3016 6823 3068
rect 6823 3016 6825 3068
rect 6769 3014 6825 3016
rect 6850 3068 6906 3070
rect 6850 3016 6852 3068
rect 6852 3016 6904 3068
rect 6904 3016 6906 3068
rect 6850 3014 6906 3016
rect 6931 3068 6987 3070
rect 6931 3016 6933 3068
rect 6933 3016 6985 3068
rect 6985 3016 6987 3068
rect 6931 3014 6987 3016
rect 7012 3068 7068 3070
rect 7012 3016 7014 3068
rect 7014 3016 7066 3068
rect 7066 3016 7068 3068
rect 7012 3014 7068 3016
rect 7094 3068 7150 3070
rect 7094 3016 7096 3068
rect 7096 3016 7148 3068
rect 7148 3016 7150 3068
rect 7094 3014 7150 3016
rect 7175 3068 7231 3070
rect 7175 3016 7177 3068
rect 7177 3016 7229 3068
rect 7229 3016 7231 3068
rect 7175 3014 7231 3016
rect 7256 3068 7312 3070
rect 7256 3016 7258 3068
rect 7258 3016 7310 3068
rect 7310 3016 7312 3068
rect 7256 3014 7312 3016
rect 7337 3068 7393 3070
rect 7337 3016 7339 3068
rect 7339 3016 7391 3068
rect 7391 3016 7393 3068
rect 7337 3014 7393 3016
rect 7418 3068 7474 3070
rect 7418 3016 7420 3068
rect 7420 3016 7472 3068
rect 7472 3016 7474 3068
rect 7418 3014 7474 3016
rect 7499 3068 7555 3070
rect 7499 3016 7501 3068
rect 7501 3016 7553 3068
rect 7553 3016 7555 3068
rect 7499 3014 7555 3016
rect 7580 3068 7636 3070
rect 7580 3016 7582 3068
rect 7582 3016 7634 3068
rect 7634 3016 7636 3068
rect 7580 3014 7636 3016
rect 7662 3068 7718 3070
rect 7662 3016 7664 3068
rect 7664 3016 7716 3068
rect 7716 3016 7718 3068
rect 7662 3014 7718 3016
rect 7743 3068 7799 3070
rect 7743 3016 7745 3068
rect 7745 3016 7797 3068
rect 7797 3016 7799 3068
rect 7743 3014 7799 3016
rect 7824 3068 7880 3070
rect 7824 3016 7826 3068
rect 7826 3016 7878 3068
rect 7878 3016 7880 3068
rect 7824 3014 7880 3016
rect 7905 3068 7961 3070
rect 7905 3016 7907 3068
rect 7907 3016 7959 3068
rect 7959 3016 7961 3068
rect 7905 3014 7961 3016
rect 7986 3068 8042 3070
rect 7986 3016 7988 3068
rect 7988 3016 8040 3068
rect 8040 3016 8042 3068
rect 7986 3014 8042 3016
rect 8067 3068 8123 3070
rect 8067 3016 8069 3068
rect 8069 3016 8121 3068
rect 8121 3016 8123 3068
rect 8067 3014 8123 3016
rect 8148 3068 8204 3070
rect 8148 3016 8150 3068
rect 8150 3016 8202 3068
rect 8202 3016 8204 3068
rect 8148 3014 8204 3016
rect 8230 3068 8286 3070
rect 8230 3016 8232 3068
rect 8232 3016 8284 3068
rect 8284 3016 8286 3068
rect 8230 3014 8286 3016
rect 8311 3068 8367 3070
rect 8311 3016 8313 3068
rect 8313 3016 8365 3068
rect 8365 3016 8367 3068
rect 8311 3014 8367 3016
rect 8392 3068 8448 3070
rect 8392 3016 8394 3068
rect 8394 3016 8446 3068
rect 8446 3016 8448 3068
rect 8392 3014 8448 3016
rect 8473 3068 8529 3070
rect 8473 3016 8475 3068
rect 8475 3016 8527 3068
rect 8527 3016 8529 3068
rect 8473 3014 8529 3016
rect 8554 3068 8610 3070
rect 8554 3016 8556 3068
rect 8556 3016 8608 3068
rect 8608 3016 8610 3068
rect 8554 3014 8610 3016
rect 8635 3068 8691 3070
rect 8635 3016 8637 3068
rect 8637 3016 8689 3068
rect 8689 3016 8691 3068
rect 8635 3014 8691 3016
rect 8716 3068 8772 3070
rect 8716 3016 8718 3068
rect 8718 3016 8770 3068
rect 8770 3016 8772 3068
rect 8716 3014 8772 3016
rect 8798 3068 8854 3070
rect 8798 3016 8800 3068
rect 8800 3016 8852 3068
rect 8852 3016 8854 3068
rect 8798 3014 8854 3016
rect 8879 3068 8935 3070
rect 8879 3016 8881 3068
rect 8881 3016 8933 3068
rect 8933 3016 8935 3068
rect 8879 3014 8935 3016
rect 8960 3068 9016 3070
rect 8960 3016 8962 3068
rect 8962 3016 9014 3068
rect 9014 3016 9016 3068
rect 8960 3014 9016 3016
rect 9041 3068 9097 3070
rect 9041 3016 9043 3068
rect 9043 3016 9095 3068
rect 9095 3016 9097 3068
rect 9041 3014 9097 3016
rect 9122 3068 9178 3070
rect 9122 3016 9124 3068
rect 9124 3016 9176 3068
rect 9176 3016 9178 3068
rect 9122 3014 9178 3016
rect 9203 3068 9259 3070
rect 9203 3016 9205 3068
rect 9205 3016 9257 3068
rect 9257 3016 9259 3068
rect 9203 3014 9259 3016
rect 9284 3068 9340 3070
rect 9284 3016 9286 3068
rect 9286 3016 9338 3068
rect 9338 3016 9340 3068
rect 9284 3014 9340 3016
rect 9366 3068 9422 3070
rect 9366 3016 9368 3068
rect 9368 3016 9420 3068
rect 9420 3016 9422 3068
rect 9366 3014 9422 3016
rect 9447 3068 9503 3070
rect 9447 3016 9449 3068
rect 9449 3016 9501 3068
rect 9501 3016 9503 3068
rect 9447 3014 9503 3016
rect 9528 3068 9584 3070
rect 9528 3016 9530 3068
rect 9530 3016 9582 3068
rect 9582 3016 9584 3068
rect 9528 3014 9584 3016
rect 9609 3068 9665 3070
rect 9609 3016 9611 3068
rect 9611 3016 9663 3068
rect 9663 3016 9665 3068
rect 9609 3014 9665 3016
rect 9690 3068 9746 3070
rect 9690 3016 9692 3068
rect 9692 3016 9744 3068
rect 9744 3016 9746 3068
rect 9690 3014 9746 3016
rect 9771 3068 9827 3070
rect 9771 3016 9773 3068
rect 9773 3016 9825 3068
rect 9825 3016 9827 3068
rect 9771 3014 9827 3016
rect 9852 3068 9908 3070
rect 9852 3016 9854 3068
rect 9854 3016 9906 3068
rect 9906 3016 9908 3068
rect 9852 3014 9908 3016
rect 9934 3068 9990 3070
rect 9934 3016 9936 3068
rect 9936 3016 9988 3068
rect 9988 3016 9990 3068
rect 9934 3014 9990 3016
rect 10015 3068 10071 3070
rect 10015 3016 10017 3068
rect 10017 3016 10069 3068
rect 10069 3016 10071 3068
rect 10015 3014 10071 3016
rect 10096 3068 10152 3070
rect 10096 3016 10098 3068
rect 10098 3016 10150 3068
rect 10150 3016 10152 3068
rect 10096 3014 10152 3016
rect 10177 3068 10233 3070
rect 10177 3016 10179 3068
rect 10179 3016 10231 3068
rect 10231 3016 10233 3068
rect 10177 3014 10233 3016
rect 10258 3068 10314 3070
rect 10258 3016 10260 3068
rect 10260 3016 10312 3068
rect 10312 3016 10314 3068
rect 10258 3014 10314 3016
rect 10339 3068 10395 3070
rect 10339 3016 10341 3068
rect 10341 3016 10393 3068
rect 10393 3016 10395 3068
rect 10339 3014 10395 3016
rect 10420 3068 10476 3070
rect 10420 3016 10422 3068
rect 10422 3016 10474 3068
rect 10474 3016 10476 3068
rect 10420 3014 10476 3016
rect 10502 3068 10558 3070
rect 10502 3016 10504 3068
rect 10504 3016 10556 3068
rect 10556 3016 10558 3068
rect 10502 3014 10558 3016
rect 10583 3068 10639 3070
rect 10583 3016 10585 3068
rect 10585 3016 10637 3068
rect 10637 3016 10639 3068
rect 10583 3014 10639 3016
rect 10664 3068 10720 3070
rect 10664 3016 10666 3068
rect 10666 3016 10718 3068
rect 10718 3016 10720 3068
rect 10664 3014 10720 3016
rect 10745 3068 10801 3070
rect 10745 3016 10747 3068
rect 10747 3016 10799 3068
rect 10799 3016 10801 3068
rect 10745 3014 10801 3016
rect 10826 3068 10882 3070
rect 10826 3016 10828 3068
rect 10828 3016 10880 3068
rect 10880 3016 10882 3068
rect 10826 3014 10882 3016
rect 10907 3068 10963 3070
rect 10907 3016 10909 3068
rect 10909 3016 10961 3068
rect 10961 3016 10963 3068
rect 10907 3014 10963 3016
rect 10988 3068 11044 3070
rect 10988 3016 10990 3068
rect 10990 3016 11042 3068
rect 11042 3016 11044 3068
rect 10988 3014 11044 3016
rect 11116 3068 11172 3070
rect 11116 3016 11118 3068
rect 11118 3016 11170 3068
rect 11170 3016 11172 3068
rect 11116 3014 11172 3016
rect 11197 3068 11253 3070
rect 11197 3016 11199 3068
rect 11199 3016 11251 3068
rect 11251 3016 11253 3068
rect 11197 3014 11253 3016
rect 11278 3068 11334 3070
rect 11278 3016 11280 3068
rect 11280 3016 11332 3068
rect 11332 3016 11334 3068
rect 11278 3014 11334 3016
rect 11359 3068 11415 3070
rect 11359 3016 11361 3068
rect 11361 3016 11413 3068
rect 11413 3016 11415 3068
rect 11359 3014 11415 3016
rect 11440 3068 11496 3070
rect 11440 3016 11442 3068
rect 11442 3016 11494 3068
rect 11494 3016 11496 3068
rect 11440 3014 11496 3016
rect 11521 3068 11577 3070
rect 11521 3016 11523 3068
rect 11523 3016 11575 3068
rect 11575 3016 11577 3068
rect 11521 3014 11577 3016
rect 11602 3068 11658 3070
rect 11602 3016 11604 3068
rect 11604 3016 11656 3068
rect 11656 3016 11658 3068
rect 11602 3014 11658 3016
rect 11684 3068 11740 3070
rect 11684 3016 11686 3068
rect 11686 3016 11738 3068
rect 11738 3016 11740 3068
rect 11684 3014 11740 3016
rect 11765 3068 11821 3070
rect 11765 3016 11767 3068
rect 11767 3016 11819 3068
rect 11819 3016 11821 3068
rect 11765 3014 11821 3016
rect 11846 3068 11902 3070
rect 11846 3016 11848 3068
rect 11848 3016 11900 3068
rect 11900 3016 11902 3068
rect 11846 3014 11902 3016
rect 11927 3068 11983 3070
rect 11927 3016 11929 3068
rect 11929 3016 11981 3068
rect 11981 3016 11983 3068
rect 11927 3014 11983 3016
rect 12008 3068 12064 3070
rect 12008 3016 12010 3068
rect 12010 3016 12062 3068
rect 12062 3016 12064 3068
rect 12008 3014 12064 3016
rect 12089 3068 12145 3070
rect 12089 3016 12091 3068
rect 12091 3016 12143 3068
rect 12143 3016 12145 3068
rect 12089 3014 12145 3016
rect 12170 3068 12226 3070
rect 12170 3016 12172 3068
rect 12172 3016 12224 3068
rect 12224 3016 12226 3068
rect 12170 3014 12226 3016
rect 12252 3068 12308 3070
rect 12252 3016 12254 3068
rect 12254 3016 12306 3068
rect 12306 3016 12308 3068
rect 12252 3014 12308 3016
rect 12333 3068 12389 3070
rect 12333 3016 12335 3068
rect 12335 3016 12387 3068
rect 12387 3016 12389 3068
rect 12333 3014 12389 3016
rect 12414 3068 12470 3070
rect 12414 3016 12416 3068
rect 12416 3016 12468 3068
rect 12468 3016 12470 3068
rect 12414 3014 12470 3016
rect 12495 3068 12551 3070
rect 12495 3016 12497 3068
rect 12497 3016 12549 3068
rect 12549 3016 12551 3068
rect 12495 3014 12551 3016
rect 12576 3068 12632 3070
rect 12576 3016 12578 3068
rect 12578 3016 12630 3068
rect 12630 3016 12632 3068
rect 12576 3014 12632 3016
rect 12657 3068 12713 3070
rect 12657 3016 12659 3068
rect 12659 3016 12711 3068
rect 12711 3016 12713 3068
rect 12657 3014 12713 3016
rect 12738 3068 12794 3070
rect 12738 3016 12740 3068
rect 12740 3016 12792 3068
rect 12792 3016 12794 3068
rect 12738 3014 12794 3016
rect 12820 3068 12876 3070
rect 12820 3016 12822 3068
rect 12822 3016 12874 3068
rect 12874 3016 12876 3068
rect 12820 3014 12876 3016
rect 12901 3068 12957 3070
rect 12901 3016 12903 3068
rect 12903 3016 12955 3068
rect 12955 3016 12957 3068
rect 12901 3014 12957 3016
rect 12982 3068 13038 3070
rect 12982 3016 12984 3068
rect 12984 3016 13036 3068
rect 13036 3016 13038 3068
rect 12982 3014 13038 3016
rect 13063 3068 13119 3070
rect 13063 3016 13065 3068
rect 13065 3016 13117 3068
rect 13117 3016 13119 3068
rect 13063 3014 13119 3016
rect 13144 3068 13200 3070
rect 13144 3016 13146 3068
rect 13146 3016 13198 3068
rect 13198 3016 13200 3068
rect 13144 3014 13200 3016
rect 13225 3068 13281 3070
rect 13225 3016 13227 3068
rect 13227 3016 13279 3068
rect 13279 3016 13281 3068
rect 13225 3014 13281 3016
rect 13306 3068 13362 3070
rect 13306 3016 13308 3068
rect 13308 3016 13360 3068
rect 13360 3016 13362 3068
rect 13306 3014 13362 3016
rect 13388 3068 13444 3070
rect 13388 3016 13390 3068
rect 13390 3016 13442 3068
rect 13442 3016 13444 3068
rect 13388 3014 13444 3016
rect 13469 3068 13525 3070
rect 13469 3016 13471 3068
rect 13471 3016 13523 3068
rect 13523 3016 13525 3068
rect 13469 3014 13525 3016
rect 13550 3068 13606 3070
rect 13550 3016 13552 3068
rect 13552 3016 13604 3068
rect 13604 3016 13606 3068
rect 13550 3014 13606 3016
rect 13631 3068 13687 3070
rect 13631 3016 13633 3068
rect 13633 3016 13685 3068
rect 13685 3016 13687 3068
rect 13631 3014 13687 3016
rect 13712 3068 13768 3070
rect 13712 3016 13714 3068
rect 13714 3016 13766 3068
rect 13766 3016 13768 3068
rect 13712 3014 13768 3016
rect 13793 3068 13849 3070
rect 13793 3016 13795 3068
rect 13795 3016 13847 3068
rect 13847 3016 13849 3068
rect 13793 3014 13849 3016
rect 13874 3068 13930 3070
rect 13874 3016 13876 3068
rect 13876 3016 13928 3068
rect 13928 3016 13930 3068
rect 13874 3014 13930 3016
rect 13956 3068 14012 3070
rect 13956 3016 13958 3068
rect 13958 3016 14010 3068
rect 14010 3016 14012 3068
rect 13956 3014 14012 3016
rect 14037 3068 14093 3070
rect 14037 3016 14039 3068
rect 14039 3016 14091 3068
rect 14091 3016 14093 3068
rect 14037 3014 14093 3016
rect 14118 3068 14174 3070
rect 14118 3016 14120 3068
rect 14120 3016 14172 3068
rect 14172 3016 14174 3068
rect 14118 3014 14174 3016
rect 14199 3068 14255 3070
rect 14199 3016 14201 3068
rect 14201 3016 14253 3068
rect 14253 3016 14255 3068
rect 14199 3014 14255 3016
rect 14280 3068 14336 3070
rect 14280 3016 14282 3068
rect 14282 3016 14334 3068
rect 14334 3016 14336 3068
rect 14280 3014 14336 3016
rect 14361 3068 14417 3070
rect 14361 3016 14363 3068
rect 14363 3016 14415 3068
rect 14415 3016 14417 3068
rect 14361 3014 14417 3016
rect 14442 3068 14498 3070
rect 14442 3016 14444 3068
rect 14444 3016 14496 3068
rect 14496 3016 14498 3068
rect 14442 3014 14498 3016
rect 14524 3068 14580 3070
rect 14524 3016 14526 3068
rect 14526 3016 14578 3068
rect 14578 3016 14580 3068
rect 14524 3014 14580 3016
rect 14605 3068 14661 3070
rect 14605 3016 14607 3068
rect 14607 3016 14659 3068
rect 14659 3016 14661 3068
rect 14605 3014 14661 3016
rect 14686 3068 14742 3070
rect 14686 3016 14688 3068
rect 14688 3016 14740 3068
rect 14740 3016 14742 3068
rect 14686 3014 14742 3016
rect 14767 3068 14823 3070
rect 14767 3016 14769 3068
rect 14769 3016 14821 3068
rect 14821 3016 14823 3068
rect 14767 3014 14823 3016
rect 14848 3068 14904 3070
rect 14848 3016 14850 3068
rect 14850 3016 14902 3068
rect 14902 3016 14904 3068
rect 14848 3014 14904 3016
rect 14929 3068 14985 3070
rect 14929 3016 14931 3068
rect 14931 3016 14983 3068
rect 14983 3016 14985 3068
rect 14929 3014 14985 3016
rect 15010 3068 15066 3070
rect 15010 3016 15012 3068
rect 15012 3016 15064 3068
rect 15064 3016 15066 3068
rect 15010 3014 15066 3016
rect 15092 3068 15148 3070
rect 15092 3016 15094 3068
rect 15094 3016 15146 3068
rect 15146 3016 15148 3068
rect 15092 3014 15148 3016
rect 15173 3068 15229 3070
rect 15173 3016 15175 3068
rect 15175 3016 15227 3068
rect 15227 3016 15229 3068
rect 15173 3014 15229 3016
rect 15254 3068 15310 3070
rect 15254 3016 15256 3068
rect 15256 3016 15308 3068
rect 15308 3016 15310 3068
rect 15254 3014 15310 3016
rect 15335 3068 15391 3070
rect 15335 3016 15337 3068
rect 15337 3016 15389 3068
rect 15389 3016 15391 3068
rect 15335 3014 15391 3016
rect 15416 3068 15472 3070
rect 15416 3016 15418 3068
rect 15418 3016 15470 3068
rect 15470 3016 15472 3068
rect 15416 3014 15472 3016
rect 15497 3068 15553 3070
rect 15497 3016 15499 3068
rect 15499 3016 15551 3068
rect 15551 3016 15553 3068
rect 15497 3014 15553 3016
rect 15578 3068 15634 3070
rect 15578 3016 15580 3068
rect 15580 3016 15632 3068
rect 15632 3016 15634 3068
rect 15578 3014 15634 3016
rect 15660 3068 15716 3070
rect 15660 3016 15662 3068
rect 15662 3016 15714 3068
rect 15714 3016 15716 3068
rect 15660 3014 15716 3016
rect 15741 3068 15797 3070
rect 15741 3016 15743 3068
rect 15743 3016 15795 3068
rect 15795 3016 15797 3068
rect 15741 3014 15797 3016
rect 15822 3068 15878 3070
rect 15822 3016 15824 3068
rect 15824 3016 15876 3068
rect 15876 3016 15878 3068
rect 15822 3014 15878 3016
rect 15903 3068 15959 3070
rect 15903 3016 15905 3068
rect 15905 3016 15957 3068
rect 15957 3016 15959 3068
rect 15903 3014 15959 3016
rect 15984 3068 16040 3070
rect 15984 3016 15986 3068
rect 15986 3016 16038 3068
rect 16038 3016 16040 3068
rect 15984 3014 16040 3016
rect 16065 3068 16121 3070
rect 16065 3016 16067 3068
rect 16067 3016 16119 3068
rect 16119 3016 16121 3068
rect 16065 3014 16121 3016
rect 16146 3068 16202 3070
rect 16146 3016 16148 3068
rect 16148 3016 16200 3068
rect 16200 3016 16202 3068
rect 16146 3014 16202 3016
rect 16228 3068 16284 3070
rect 16228 3016 16230 3068
rect 16230 3016 16282 3068
rect 16282 3016 16284 3068
rect 16228 3014 16284 3016
rect 16309 3068 16365 3070
rect 16309 3016 16311 3068
rect 16311 3016 16363 3068
rect 16363 3016 16365 3068
rect 16309 3014 16365 3016
rect 16390 3068 16446 3070
rect 16390 3016 16392 3068
rect 16392 3016 16444 3068
rect 16444 3016 16446 3068
rect 16390 3014 16446 3016
rect 16471 3068 16527 3070
rect 16471 3016 16473 3068
rect 16473 3016 16525 3068
rect 16525 3016 16527 3068
rect 16471 3014 16527 3016
rect 16552 3068 16608 3070
rect 16552 3016 16554 3068
rect 16554 3016 16606 3068
rect 16606 3016 16608 3068
rect 16552 3014 16608 3016
rect 16633 3068 16689 3070
rect 16633 3016 16635 3068
rect 16635 3016 16687 3068
rect 16687 3016 16689 3068
rect 16633 3014 16689 3016
rect 16714 3068 16770 3070
rect 16714 3016 16716 3068
rect 16716 3016 16768 3068
rect 16768 3016 16770 3068
rect 16714 3014 16770 3016
rect 16796 3068 16852 3070
rect 16796 3016 16798 3068
rect 16798 3016 16850 3068
rect 16850 3016 16852 3068
rect 16796 3014 16852 3016
rect 16877 3068 16933 3070
rect 16877 3016 16879 3068
rect 16879 3016 16931 3068
rect 16931 3016 16933 3068
rect 16877 3014 16933 3016
rect 16958 3068 17014 3070
rect 16958 3016 16960 3068
rect 16960 3016 17012 3068
rect 17012 3016 17014 3068
rect 16958 3014 17014 3016
rect 17039 3068 17095 3070
rect 17039 3016 17041 3068
rect 17041 3016 17093 3068
rect 17093 3016 17095 3068
rect 17039 3014 17095 3016
rect 17120 3068 17176 3070
rect 17120 3016 17122 3068
rect 17122 3016 17174 3068
rect 17174 3016 17176 3068
rect 17120 3014 17176 3016
rect 17201 3068 17257 3070
rect 17201 3016 17203 3068
rect 17203 3016 17255 3068
rect 17255 3016 17257 3068
rect 17201 3014 17257 3016
rect 17282 3068 17338 3070
rect 17282 3016 17284 3068
rect 17284 3016 17336 3068
rect 17336 3016 17338 3068
rect 17282 3014 17338 3016
rect 17364 3068 17420 3070
rect 17364 3016 17366 3068
rect 17366 3016 17418 3068
rect 17418 3016 17420 3068
rect 17364 3014 17420 3016
rect 17445 3068 17501 3070
rect 17445 3016 17447 3068
rect 17447 3016 17499 3068
rect 17499 3016 17501 3068
rect 17445 3014 17501 3016
rect 17526 3068 17582 3070
rect 17526 3016 17528 3068
rect 17528 3016 17580 3068
rect 17580 3016 17582 3068
rect 17526 3014 17582 3016
rect 17607 3068 17663 3070
rect 17607 3016 17609 3068
rect 17609 3016 17661 3068
rect 17661 3016 17663 3068
rect 17607 3014 17663 3016
rect 17688 3068 17744 3070
rect 17688 3016 17690 3068
rect 17690 3016 17742 3068
rect 17742 3016 17744 3068
rect 17688 3014 17744 3016
rect 17769 3068 17825 3070
rect 17769 3016 17771 3068
rect 17771 3016 17823 3068
rect 17823 3016 17825 3068
rect 17769 3014 17825 3016
rect 17850 3068 17906 3070
rect 17850 3016 17852 3068
rect 17852 3016 17904 3068
rect 17904 3016 17906 3068
rect 17850 3014 17906 3016
rect 17932 3068 17988 3070
rect 17932 3016 17934 3068
rect 17934 3016 17986 3068
rect 17986 3016 17988 3068
rect 17932 3014 17988 3016
rect 18013 3068 18069 3070
rect 18013 3016 18015 3068
rect 18015 3016 18067 3068
rect 18067 3016 18069 3068
rect 18013 3014 18069 3016
rect 18094 3068 18150 3070
rect 18094 3016 18096 3068
rect 18096 3016 18148 3068
rect 18148 3016 18150 3068
rect 18094 3014 18150 3016
rect 18175 3068 18231 3070
rect 18175 3016 18177 3068
rect 18177 3016 18229 3068
rect 18229 3016 18231 3068
rect 18175 3014 18231 3016
rect 18256 3068 18312 3070
rect 18256 3016 18258 3068
rect 18258 3016 18310 3068
rect 18310 3016 18312 3068
rect 18256 3014 18312 3016
rect 18337 3068 18393 3070
rect 18337 3016 18339 3068
rect 18339 3016 18391 3068
rect 18391 3016 18393 3068
rect 18337 3014 18393 3016
rect 18418 3068 18474 3070
rect 18418 3016 18420 3068
rect 18420 3016 18472 3068
rect 18472 3016 18474 3068
rect 18418 3014 18474 3016
rect 18500 3068 18556 3070
rect 18500 3016 18502 3068
rect 18502 3016 18554 3068
rect 18554 3016 18556 3068
rect 18500 3014 18556 3016
rect 18581 3068 18637 3070
rect 18581 3016 18583 3068
rect 18583 3016 18635 3068
rect 18635 3016 18637 3068
rect 18581 3014 18637 3016
rect 18662 3068 18718 3070
rect 18662 3016 18664 3068
rect 18664 3016 18716 3068
rect 18716 3016 18718 3068
rect 18662 3014 18718 3016
rect 18743 3068 18799 3070
rect 18743 3016 18745 3068
rect 18745 3016 18797 3068
rect 18797 3016 18799 3068
rect 18743 3014 18799 3016
rect 18824 3068 18880 3070
rect 18824 3016 18826 3068
rect 18826 3016 18878 3068
rect 18878 3016 18880 3068
rect 18824 3014 18880 3016
rect 18905 3068 18961 3070
rect 18905 3016 18907 3068
rect 18907 3016 18959 3068
rect 18959 3016 18961 3068
rect 18905 3014 18961 3016
rect 18986 3068 19042 3070
rect 18986 3016 18988 3068
rect 18988 3016 19040 3068
rect 19040 3016 19042 3068
rect 18986 3014 19042 3016
rect 19068 3068 19124 3070
rect 19068 3016 19070 3068
rect 19070 3016 19122 3068
rect 19122 3016 19124 3068
rect 19068 3014 19124 3016
rect 19149 3068 19205 3070
rect 19149 3016 19151 3068
rect 19151 3016 19203 3068
rect 19203 3016 19205 3068
rect 19149 3014 19205 3016
rect 19230 3068 19286 3070
rect 19230 3016 19232 3068
rect 19232 3016 19284 3068
rect 19284 3016 19286 3068
rect 19230 3014 19286 3016
rect 19311 3068 19367 3070
rect 19311 3016 19313 3068
rect 19313 3016 19365 3068
rect 19365 3016 19367 3068
rect 19311 3014 19367 3016
rect 19392 3068 19448 3070
rect 19392 3016 19394 3068
rect 19394 3016 19446 3068
rect 19446 3016 19448 3068
rect 19392 3014 19448 3016
rect 19473 3068 19529 3070
rect 19473 3016 19475 3068
rect 19475 3016 19527 3068
rect 19527 3016 19529 3068
rect 19473 3014 19529 3016
rect 19554 3068 19610 3070
rect 19554 3016 19556 3068
rect 19556 3016 19608 3068
rect 19608 3016 19610 3068
rect 19554 3014 19610 3016
rect 19636 3068 19692 3070
rect 19636 3016 19638 3068
rect 19638 3016 19690 3068
rect 19690 3016 19692 3068
rect 19636 3014 19692 3016
rect 19717 3068 19773 3070
rect 19717 3016 19719 3068
rect 19719 3016 19771 3068
rect 19771 3016 19773 3068
rect 19717 3014 19773 3016
rect 19798 3068 19854 3070
rect 19798 3016 19800 3068
rect 19800 3016 19852 3068
rect 19852 3016 19854 3068
rect 19798 3014 19854 3016
rect 19879 3068 19935 3070
rect 19879 3016 19881 3068
rect 19881 3016 19933 3068
rect 19933 3016 19935 3068
rect 19879 3014 19935 3016
rect 19960 3068 20016 3070
rect 19960 3016 19962 3068
rect 19962 3016 20014 3068
rect 20014 3016 20016 3068
rect 19960 3014 20016 3016
rect 20041 3068 20097 3070
rect 20041 3016 20043 3068
rect 20043 3016 20095 3068
rect 20095 3016 20097 3068
rect 20041 3014 20097 3016
rect 20122 3068 20178 3070
rect 20122 3016 20124 3068
rect 20124 3016 20176 3068
rect 20176 3016 20178 3068
rect 20122 3014 20178 3016
rect 20204 3068 20260 3070
rect 20204 3016 20206 3068
rect 20206 3016 20258 3068
rect 20258 3016 20260 3068
rect 20204 3014 20260 3016
rect 20285 3068 20341 3070
rect 20285 3016 20287 3068
rect 20287 3016 20339 3068
rect 20339 3016 20341 3068
rect 20285 3014 20341 3016
rect 20366 3068 20422 3070
rect 20366 3016 20368 3068
rect 20368 3016 20420 3068
rect 20420 3016 20422 3068
rect 20366 3014 20422 3016
rect 20447 3068 20503 3070
rect 20447 3016 20449 3068
rect 20449 3016 20501 3068
rect 20501 3016 20503 3068
rect 20447 3014 20503 3016
rect 20528 3068 20584 3070
rect 20528 3016 20530 3068
rect 20530 3016 20582 3068
rect 20582 3016 20584 3068
rect 20528 3014 20584 3016
rect 20609 3068 20665 3070
rect 20609 3016 20611 3068
rect 20611 3016 20663 3068
rect 20663 3016 20665 3068
rect 20609 3014 20665 3016
rect 20690 3068 20746 3070
rect 20690 3016 20692 3068
rect 20692 3016 20744 3068
rect 20744 3016 20746 3068
rect 20690 3014 20746 3016
rect 20772 3068 20828 3070
rect 20772 3016 20774 3068
rect 20774 3016 20826 3068
rect 20826 3016 20828 3068
rect 20772 3014 20828 3016
rect 20853 3068 20909 3070
rect 20853 3016 20855 3068
rect 20855 3016 20907 3068
rect 20907 3016 20909 3068
rect 20853 3014 20909 3016
rect 20934 3068 20990 3070
rect 20934 3016 20936 3068
rect 20936 3016 20988 3068
rect 20988 3016 20990 3068
rect 20934 3014 20990 3016
rect 21015 3068 21071 3070
rect 21015 3016 21017 3068
rect 21017 3016 21069 3068
rect 21069 3016 21071 3068
rect 21015 3014 21071 3016
rect 21096 3068 21152 3070
rect 21096 3016 21098 3068
rect 21098 3016 21150 3068
rect 21150 3016 21152 3068
rect 21096 3014 21152 3016
rect 21177 3068 21233 3070
rect 21177 3016 21179 3068
rect 21179 3016 21231 3068
rect 21231 3016 21233 3068
rect 21177 3014 21233 3016
rect 21258 3068 21314 3070
rect 21258 3016 21260 3068
rect 21260 3016 21312 3068
rect 21312 3016 21314 3068
rect 21258 3014 21314 3016
rect 21340 3068 21396 3070
rect 21340 3016 21342 3068
rect 21342 3016 21394 3068
rect 21394 3016 21396 3068
rect 21340 3014 21396 3016
rect 21421 3068 21477 3070
rect 21421 3016 21423 3068
rect 21423 3016 21475 3068
rect 21475 3016 21477 3068
rect 21421 3014 21477 3016
rect 21502 3068 21558 3070
rect 21502 3016 21504 3068
rect 21504 3016 21556 3068
rect 21556 3016 21558 3068
rect 21502 3014 21558 3016
rect 21583 3068 21639 3070
rect 21583 3016 21585 3068
rect 21585 3016 21637 3068
rect 21637 3016 21639 3068
rect 21583 3014 21639 3016
rect 21664 3068 21720 3070
rect 21664 3016 21666 3068
rect 21666 3016 21718 3068
rect 21718 3016 21720 3068
rect 21664 3014 21720 3016
rect 21745 3068 21801 3070
rect 21745 3016 21747 3068
rect 21747 3016 21799 3068
rect 21799 3016 21801 3068
rect 21745 3014 21801 3016
rect 21826 3068 21882 3070
rect 21826 3016 21828 3068
rect 21828 3016 21880 3068
rect 21880 3016 21882 3068
rect 21826 3014 21882 3016
rect 21908 3068 21964 3070
rect 21908 3016 21910 3068
rect 21910 3016 21962 3068
rect 21962 3016 21964 3068
rect 21908 3014 21964 3016
rect 21989 3068 22045 3070
rect 21989 3016 21991 3068
rect 21991 3016 22043 3068
rect 22043 3016 22045 3068
rect 21989 3014 22045 3016
rect 22070 3068 22126 3070
rect 22070 3016 22072 3068
rect 22072 3016 22124 3068
rect 22124 3016 22126 3068
rect 22070 3014 22126 3016
rect 22151 3068 22207 3070
rect 22151 3016 22153 3068
rect 22153 3016 22205 3068
rect 22205 3016 22207 3068
rect 22151 3014 22207 3016
rect 22232 3068 22288 3070
rect 22232 3016 22234 3068
rect 22234 3016 22286 3068
rect 22286 3016 22288 3068
rect 22232 3014 22288 3016
rect 22313 3068 22369 3070
rect 22313 3016 22315 3068
rect 22315 3016 22367 3068
rect 22367 3016 22369 3068
rect 22313 3014 22369 3016
rect 22394 3068 22450 3070
rect 22394 3016 22396 3068
rect 22396 3016 22448 3068
rect 22448 3016 22450 3068
rect 22394 3014 22450 3016
rect 22476 3068 22532 3070
rect 22476 3016 22478 3068
rect 22478 3016 22530 3068
rect 22530 3016 22532 3068
rect 22476 3014 22532 3016
rect 22557 3068 22613 3070
rect 22557 3016 22559 3068
rect 22559 3016 22611 3068
rect 22611 3016 22613 3068
rect 22557 3014 22613 3016
rect 22638 3068 22694 3070
rect 22638 3016 22640 3068
rect 22640 3016 22692 3068
rect 22692 3016 22694 3068
rect 22638 3014 22694 3016
rect 22719 3068 22775 3070
rect 22719 3016 22721 3068
rect 22721 3016 22773 3068
rect 22773 3016 22775 3068
rect 22719 3014 22775 3016
rect 22800 3068 22856 3070
rect 22800 3016 22802 3068
rect 22802 3016 22854 3068
rect 22854 3016 22856 3068
rect 22800 3014 22856 3016
rect 22881 3068 22937 3070
rect 22881 3016 22883 3068
rect 22883 3016 22935 3068
rect 22935 3016 22937 3068
rect 22881 3014 22937 3016
rect 22962 3068 23018 3070
rect 22962 3016 22964 3068
rect 22964 3016 23016 3068
rect 23016 3016 23018 3068
rect 22962 3014 23018 3016
rect 23044 3068 23100 3070
rect 23044 3016 23046 3068
rect 23046 3016 23098 3068
rect 23098 3016 23100 3068
rect 23044 3014 23100 3016
rect 23125 3068 23181 3070
rect 23125 3016 23127 3068
rect 23127 3016 23179 3068
rect 23179 3016 23181 3068
rect 23125 3014 23181 3016
rect 23206 3068 23262 3070
rect 23206 3016 23208 3068
rect 23208 3016 23260 3068
rect 23260 3016 23262 3068
rect 23206 3014 23262 3016
rect 23287 3068 23343 3070
rect 23287 3016 23289 3068
rect 23289 3016 23341 3068
rect 23341 3016 23343 3068
rect 23287 3014 23343 3016
rect 23368 3068 23424 3070
rect 23368 3016 23370 3068
rect 23370 3016 23422 3068
rect 23422 3016 23424 3068
rect 23368 3014 23424 3016
rect 23449 3068 23505 3070
rect 23449 3016 23451 3068
rect 23451 3016 23503 3068
rect 23503 3016 23505 3068
rect 23449 3014 23505 3016
rect 23530 3068 23586 3070
rect 23530 3016 23532 3068
rect 23532 3016 23584 3068
rect 23584 3016 23586 3068
rect 23530 3014 23586 3016
rect 23612 3068 23668 3070
rect 23612 3016 23614 3068
rect 23614 3016 23666 3068
rect 23666 3016 23668 3068
rect 23612 3014 23668 3016
rect 23693 3068 23749 3070
rect 23693 3016 23695 3068
rect 23695 3016 23747 3068
rect 23747 3016 23749 3068
rect 23693 3014 23749 3016
rect 23774 3068 23830 3070
rect 23774 3016 23776 3068
rect 23776 3016 23828 3068
rect 23828 3016 23830 3068
rect 23774 3014 23830 3016
rect 23855 3068 23911 3070
rect 23855 3016 23857 3068
rect 23857 3016 23909 3068
rect 23909 3016 23911 3068
rect 23855 3014 23911 3016
rect 23936 3068 23992 3070
rect 23936 3016 23938 3068
rect 23938 3016 23990 3068
rect 23990 3016 23992 3068
rect 23936 3014 23992 3016
rect 24017 3068 24073 3070
rect 24017 3016 24019 3068
rect 24019 3016 24071 3068
rect 24071 3016 24073 3068
rect 24017 3014 24073 3016
rect 24098 3068 24154 3070
rect 24098 3016 24100 3068
rect 24100 3016 24152 3068
rect 24152 3016 24154 3068
rect 24098 3014 24154 3016
rect 24180 3068 24236 3070
rect 24180 3016 24182 3068
rect 24182 3016 24234 3068
rect 24234 3016 24236 3068
rect 24180 3014 24236 3016
rect 24261 3068 24317 3070
rect 24261 3016 24263 3068
rect 24263 3016 24315 3068
rect 24315 3016 24317 3068
rect 24261 3014 24317 3016
rect 24342 3068 24398 3070
rect 24342 3016 24344 3068
rect 24344 3016 24396 3068
rect 24396 3016 24398 3068
rect 24342 3014 24398 3016
rect 24423 3068 24479 3070
rect 24423 3016 24425 3068
rect 24425 3016 24477 3068
rect 24477 3016 24479 3068
rect 24423 3014 24479 3016
rect 24504 3068 24560 3070
rect 24504 3016 24506 3068
rect 24506 3016 24558 3068
rect 24558 3016 24560 3068
rect 24504 3014 24560 3016
rect 24585 3068 24641 3070
rect 24585 3016 24587 3068
rect 24587 3016 24639 3068
rect 24639 3016 24641 3068
rect 24585 3014 24641 3016
rect 24666 3068 24722 3070
rect 24666 3016 24668 3068
rect 24668 3016 24720 3068
rect 24720 3016 24722 3068
rect 24666 3014 24722 3016
rect 3036 2964 3092 2966
rect 3036 2912 3038 2964
rect 3038 2912 3090 2964
rect 3090 2912 3092 2964
rect 3036 2910 3092 2912
rect 3118 2964 3174 2966
rect 3118 2912 3120 2964
rect 3120 2912 3172 2964
rect 3172 2912 3174 2964
rect 3118 2910 3174 2912
rect 3199 2964 3255 2966
rect 3199 2912 3201 2964
rect 3201 2912 3253 2964
rect 3253 2912 3255 2964
rect 3199 2910 3255 2912
rect 3280 2964 3336 2966
rect 3280 2912 3282 2964
rect 3282 2912 3334 2964
rect 3334 2912 3336 2964
rect 3280 2910 3336 2912
rect 3361 2964 3417 2966
rect 3361 2912 3363 2964
rect 3363 2912 3415 2964
rect 3415 2912 3417 2964
rect 3361 2910 3417 2912
rect 3442 2964 3498 2966
rect 3442 2912 3444 2964
rect 3444 2912 3496 2964
rect 3496 2912 3498 2964
rect 3442 2910 3498 2912
rect 3523 2964 3579 2966
rect 3523 2912 3525 2964
rect 3525 2912 3577 2964
rect 3577 2912 3579 2964
rect 3523 2910 3579 2912
rect 3604 2964 3660 2966
rect 3604 2912 3606 2964
rect 3606 2912 3658 2964
rect 3658 2912 3660 2964
rect 3604 2910 3660 2912
rect 3686 2964 3742 2966
rect 3686 2912 3688 2964
rect 3688 2912 3740 2964
rect 3740 2912 3742 2964
rect 3686 2910 3742 2912
rect 3767 2964 3823 2966
rect 3767 2912 3769 2964
rect 3769 2912 3821 2964
rect 3821 2912 3823 2964
rect 3767 2910 3823 2912
rect 3848 2964 3904 2966
rect 3848 2912 3850 2964
rect 3850 2912 3902 2964
rect 3902 2912 3904 2964
rect 3848 2910 3904 2912
rect 3929 2964 3985 2966
rect 3929 2912 3931 2964
rect 3931 2912 3983 2964
rect 3983 2912 3985 2964
rect 3929 2910 3985 2912
rect 4010 2964 4066 2966
rect 4010 2912 4012 2964
rect 4012 2912 4064 2964
rect 4064 2912 4066 2964
rect 4010 2910 4066 2912
rect 4091 2964 4147 2966
rect 4091 2912 4093 2964
rect 4093 2912 4145 2964
rect 4145 2912 4147 2964
rect 4091 2910 4147 2912
rect 4172 2964 4228 2966
rect 4172 2912 4174 2964
rect 4174 2912 4226 2964
rect 4226 2912 4228 2964
rect 4172 2910 4228 2912
rect 4254 2964 4310 2966
rect 4254 2912 4256 2964
rect 4256 2912 4308 2964
rect 4308 2912 4310 2964
rect 4254 2910 4310 2912
rect 4335 2964 4391 2966
rect 4335 2912 4337 2964
rect 4337 2912 4389 2964
rect 4389 2912 4391 2964
rect 4335 2910 4391 2912
rect 4416 2964 4472 2966
rect 4416 2912 4418 2964
rect 4418 2912 4470 2964
rect 4470 2912 4472 2964
rect 4416 2910 4472 2912
rect 4497 2964 4553 2966
rect 4497 2912 4499 2964
rect 4499 2912 4551 2964
rect 4551 2912 4553 2964
rect 4497 2910 4553 2912
rect 4578 2964 4634 2966
rect 4578 2912 4580 2964
rect 4580 2912 4632 2964
rect 4632 2912 4634 2964
rect 4578 2910 4634 2912
rect 4659 2964 4715 2966
rect 4659 2912 4661 2964
rect 4661 2912 4713 2964
rect 4713 2912 4715 2964
rect 4659 2910 4715 2912
rect 4740 2964 4796 2966
rect 4740 2912 4742 2964
rect 4742 2912 4794 2964
rect 4794 2912 4796 2964
rect 4740 2910 4796 2912
rect 4822 2964 4878 2966
rect 4822 2912 4824 2964
rect 4824 2912 4876 2964
rect 4876 2912 4878 2964
rect 4822 2910 4878 2912
rect 4903 2964 4959 2966
rect 4903 2912 4905 2964
rect 4905 2912 4957 2964
rect 4957 2912 4959 2964
rect 4903 2910 4959 2912
rect 4984 2964 5040 2966
rect 4984 2912 4986 2964
rect 4986 2912 5038 2964
rect 5038 2912 5040 2964
rect 4984 2910 5040 2912
rect 5065 2964 5121 2966
rect 5065 2912 5067 2964
rect 5067 2912 5119 2964
rect 5119 2912 5121 2964
rect 5065 2910 5121 2912
rect 5146 2964 5202 2966
rect 5146 2912 5148 2964
rect 5148 2912 5200 2964
rect 5200 2912 5202 2964
rect 5146 2910 5202 2912
rect 5227 2964 5283 2966
rect 5227 2912 5229 2964
rect 5229 2912 5281 2964
rect 5281 2912 5283 2964
rect 5227 2910 5283 2912
rect 5308 2964 5364 2966
rect 5308 2912 5310 2964
rect 5310 2912 5362 2964
rect 5362 2912 5364 2964
rect 5308 2910 5364 2912
rect 5390 2964 5446 2966
rect 5390 2912 5392 2964
rect 5392 2912 5444 2964
rect 5444 2912 5446 2964
rect 5390 2910 5446 2912
rect 5471 2964 5527 2966
rect 5471 2912 5473 2964
rect 5473 2912 5525 2964
rect 5525 2912 5527 2964
rect 5471 2910 5527 2912
rect 5552 2964 5608 2966
rect 5552 2912 5554 2964
rect 5554 2912 5606 2964
rect 5606 2912 5608 2964
rect 5552 2910 5608 2912
rect 5633 2964 5689 2966
rect 5633 2912 5635 2964
rect 5635 2912 5687 2964
rect 5687 2912 5689 2964
rect 5633 2910 5689 2912
rect 5714 2964 5770 2966
rect 5714 2912 5716 2964
rect 5716 2912 5768 2964
rect 5768 2912 5770 2964
rect 5714 2910 5770 2912
rect 5795 2964 5851 2966
rect 5795 2912 5797 2964
rect 5797 2912 5849 2964
rect 5849 2912 5851 2964
rect 5795 2910 5851 2912
rect 5876 2964 5932 2966
rect 5876 2912 5878 2964
rect 5878 2912 5930 2964
rect 5930 2912 5932 2964
rect 5876 2910 5932 2912
rect 5958 2964 6014 2966
rect 5958 2912 5960 2964
rect 5960 2912 6012 2964
rect 6012 2912 6014 2964
rect 5958 2910 6014 2912
rect 6039 2964 6095 2966
rect 6039 2912 6041 2964
rect 6041 2912 6093 2964
rect 6093 2912 6095 2964
rect 6039 2910 6095 2912
rect 6120 2964 6176 2966
rect 6120 2912 6122 2964
rect 6122 2912 6174 2964
rect 6174 2912 6176 2964
rect 6120 2910 6176 2912
rect 6201 2964 6257 2966
rect 6201 2912 6203 2964
rect 6203 2912 6255 2964
rect 6255 2912 6257 2964
rect 6201 2910 6257 2912
rect 6282 2964 6338 2966
rect 6282 2912 6284 2964
rect 6284 2912 6336 2964
rect 6336 2912 6338 2964
rect 6282 2910 6338 2912
rect 6363 2964 6419 2966
rect 6363 2912 6365 2964
rect 6365 2912 6417 2964
rect 6417 2912 6419 2964
rect 6363 2910 6419 2912
rect 6444 2964 6500 2966
rect 6444 2912 6446 2964
rect 6446 2912 6498 2964
rect 6498 2912 6500 2964
rect 6444 2910 6500 2912
rect 6526 2964 6582 2966
rect 6526 2912 6528 2964
rect 6528 2912 6580 2964
rect 6580 2912 6582 2964
rect 6526 2910 6582 2912
rect 6607 2964 6663 2966
rect 6607 2912 6609 2964
rect 6609 2912 6661 2964
rect 6661 2912 6663 2964
rect 6607 2910 6663 2912
rect 6688 2964 6744 2966
rect 6688 2912 6690 2964
rect 6690 2912 6742 2964
rect 6742 2912 6744 2964
rect 6688 2910 6744 2912
rect 6769 2964 6825 2966
rect 6769 2912 6771 2964
rect 6771 2912 6823 2964
rect 6823 2912 6825 2964
rect 6769 2910 6825 2912
rect 6850 2964 6906 2966
rect 6850 2912 6852 2964
rect 6852 2912 6904 2964
rect 6904 2912 6906 2964
rect 6850 2910 6906 2912
rect 6931 2964 6987 2966
rect 6931 2912 6933 2964
rect 6933 2912 6985 2964
rect 6985 2912 6987 2964
rect 6931 2910 6987 2912
rect 7012 2964 7068 2966
rect 7012 2912 7014 2964
rect 7014 2912 7066 2964
rect 7066 2912 7068 2964
rect 7012 2910 7068 2912
rect 7094 2964 7150 2966
rect 7094 2912 7096 2964
rect 7096 2912 7148 2964
rect 7148 2912 7150 2964
rect 7094 2910 7150 2912
rect 7175 2964 7231 2966
rect 7175 2912 7177 2964
rect 7177 2912 7229 2964
rect 7229 2912 7231 2964
rect 7175 2910 7231 2912
rect 7256 2964 7312 2966
rect 7256 2912 7258 2964
rect 7258 2912 7310 2964
rect 7310 2912 7312 2964
rect 7256 2910 7312 2912
rect 7337 2964 7393 2966
rect 7337 2912 7339 2964
rect 7339 2912 7391 2964
rect 7391 2912 7393 2964
rect 7337 2910 7393 2912
rect 7418 2964 7474 2966
rect 7418 2912 7420 2964
rect 7420 2912 7472 2964
rect 7472 2912 7474 2964
rect 7418 2910 7474 2912
rect 7499 2964 7555 2966
rect 7499 2912 7501 2964
rect 7501 2912 7553 2964
rect 7553 2912 7555 2964
rect 7499 2910 7555 2912
rect 7580 2964 7636 2966
rect 7580 2912 7582 2964
rect 7582 2912 7634 2964
rect 7634 2912 7636 2964
rect 7580 2910 7636 2912
rect 7662 2964 7718 2966
rect 7662 2912 7664 2964
rect 7664 2912 7716 2964
rect 7716 2912 7718 2964
rect 7662 2910 7718 2912
rect 7743 2964 7799 2966
rect 7743 2912 7745 2964
rect 7745 2912 7797 2964
rect 7797 2912 7799 2964
rect 7743 2910 7799 2912
rect 7824 2964 7880 2966
rect 7824 2912 7826 2964
rect 7826 2912 7878 2964
rect 7878 2912 7880 2964
rect 7824 2910 7880 2912
rect 7905 2964 7961 2966
rect 7905 2912 7907 2964
rect 7907 2912 7959 2964
rect 7959 2912 7961 2964
rect 7905 2910 7961 2912
rect 7986 2964 8042 2966
rect 7986 2912 7988 2964
rect 7988 2912 8040 2964
rect 8040 2912 8042 2964
rect 7986 2910 8042 2912
rect 8067 2964 8123 2966
rect 8067 2912 8069 2964
rect 8069 2912 8121 2964
rect 8121 2912 8123 2964
rect 8067 2910 8123 2912
rect 8148 2964 8204 2966
rect 8148 2912 8150 2964
rect 8150 2912 8202 2964
rect 8202 2912 8204 2964
rect 8148 2910 8204 2912
rect 8230 2964 8286 2966
rect 8230 2912 8232 2964
rect 8232 2912 8284 2964
rect 8284 2912 8286 2964
rect 8230 2910 8286 2912
rect 8311 2964 8367 2966
rect 8311 2912 8313 2964
rect 8313 2912 8365 2964
rect 8365 2912 8367 2964
rect 8311 2910 8367 2912
rect 8392 2964 8448 2966
rect 8392 2912 8394 2964
rect 8394 2912 8446 2964
rect 8446 2912 8448 2964
rect 8392 2910 8448 2912
rect 8473 2964 8529 2966
rect 8473 2912 8475 2964
rect 8475 2912 8527 2964
rect 8527 2912 8529 2964
rect 8473 2910 8529 2912
rect 8554 2964 8610 2966
rect 8554 2912 8556 2964
rect 8556 2912 8608 2964
rect 8608 2912 8610 2964
rect 8554 2910 8610 2912
rect 8635 2964 8691 2966
rect 8635 2912 8637 2964
rect 8637 2912 8689 2964
rect 8689 2912 8691 2964
rect 8635 2910 8691 2912
rect 8716 2964 8772 2966
rect 8716 2912 8718 2964
rect 8718 2912 8770 2964
rect 8770 2912 8772 2964
rect 8716 2910 8772 2912
rect 8798 2964 8854 2966
rect 8798 2912 8800 2964
rect 8800 2912 8852 2964
rect 8852 2912 8854 2964
rect 8798 2910 8854 2912
rect 8879 2964 8935 2966
rect 8879 2912 8881 2964
rect 8881 2912 8933 2964
rect 8933 2912 8935 2964
rect 8879 2910 8935 2912
rect 8960 2964 9016 2966
rect 8960 2912 8962 2964
rect 8962 2912 9014 2964
rect 9014 2912 9016 2964
rect 8960 2910 9016 2912
rect 9041 2964 9097 2966
rect 9041 2912 9043 2964
rect 9043 2912 9095 2964
rect 9095 2912 9097 2964
rect 9041 2910 9097 2912
rect 9122 2964 9178 2966
rect 9122 2912 9124 2964
rect 9124 2912 9176 2964
rect 9176 2912 9178 2964
rect 9122 2910 9178 2912
rect 9203 2964 9259 2966
rect 9203 2912 9205 2964
rect 9205 2912 9257 2964
rect 9257 2912 9259 2964
rect 9203 2910 9259 2912
rect 9284 2964 9340 2966
rect 9284 2912 9286 2964
rect 9286 2912 9338 2964
rect 9338 2912 9340 2964
rect 9284 2910 9340 2912
rect 9366 2964 9422 2966
rect 9366 2912 9368 2964
rect 9368 2912 9420 2964
rect 9420 2912 9422 2964
rect 9366 2910 9422 2912
rect 9447 2964 9503 2966
rect 9447 2912 9449 2964
rect 9449 2912 9501 2964
rect 9501 2912 9503 2964
rect 9447 2910 9503 2912
rect 9528 2964 9584 2966
rect 9528 2912 9530 2964
rect 9530 2912 9582 2964
rect 9582 2912 9584 2964
rect 9528 2910 9584 2912
rect 9609 2964 9665 2966
rect 9609 2912 9611 2964
rect 9611 2912 9663 2964
rect 9663 2912 9665 2964
rect 9609 2910 9665 2912
rect 9690 2964 9746 2966
rect 9690 2912 9692 2964
rect 9692 2912 9744 2964
rect 9744 2912 9746 2964
rect 9690 2910 9746 2912
rect 9771 2964 9827 2966
rect 9771 2912 9773 2964
rect 9773 2912 9825 2964
rect 9825 2912 9827 2964
rect 9771 2910 9827 2912
rect 9852 2964 9908 2966
rect 9852 2912 9854 2964
rect 9854 2912 9906 2964
rect 9906 2912 9908 2964
rect 9852 2910 9908 2912
rect 9934 2964 9990 2966
rect 9934 2912 9936 2964
rect 9936 2912 9988 2964
rect 9988 2912 9990 2964
rect 9934 2910 9990 2912
rect 10015 2964 10071 2966
rect 10015 2912 10017 2964
rect 10017 2912 10069 2964
rect 10069 2912 10071 2964
rect 10015 2910 10071 2912
rect 10096 2964 10152 2966
rect 10096 2912 10098 2964
rect 10098 2912 10150 2964
rect 10150 2912 10152 2964
rect 10096 2910 10152 2912
rect 10177 2964 10233 2966
rect 10177 2912 10179 2964
rect 10179 2912 10231 2964
rect 10231 2912 10233 2964
rect 10177 2910 10233 2912
rect 10258 2964 10314 2966
rect 10258 2912 10260 2964
rect 10260 2912 10312 2964
rect 10312 2912 10314 2964
rect 10258 2910 10314 2912
rect 10339 2964 10395 2966
rect 10339 2912 10341 2964
rect 10341 2912 10393 2964
rect 10393 2912 10395 2964
rect 10339 2910 10395 2912
rect 10420 2964 10476 2966
rect 10420 2912 10422 2964
rect 10422 2912 10474 2964
rect 10474 2912 10476 2964
rect 10420 2910 10476 2912
rect 10502 2964 10558 2966
rect 10502 2912 10504 2964
rect 10504 2912 10556 2964
rect 10556 2912 10558 2964
rect 10502 2910 10558 2912
rect 10583 2964 10639 2966
rect 10583 2912 10585 2964
rect 10585 2912 10637 2964
rect 10637 2912 10639 2964
rect 10583 2910 10639 2912
rect 10664 2964 10720 2966
rect 10664 2912 10666 2964
rect 10666 2912 10718 2964
rect 10718 2912 10720 2964
rect 10664 2910 10720 2912
rect 10745 2964 10801 2966
rect 10745 2912 10747 2964
rect 10747 2912 10799 2964
rect 10799 2912 10801 2964
rect 10745 2910 10801 2912
rect 10826 2964 10882 2966
rect 10826 2912 10828 2964
rect 10828 2912 10880 2964
rect 10880 2912 10882 2964
rect 10826 2910 10882 2912
rect 10907 2964 10963 2966
rect 10907 2912 10909 2964
rect 10909 2912 10961 2964
rect 10961 2912 10963 2964
rect 10907 2910 10963 2912
rect 10988 2964 11044 2966
rect 10988 2912 10990 2964
rect 10990 2912 11042 2964
rect 11042 2912 11044 2964
rect 10988 2910 11044 2912
rect 11116 2964 11172 2966
rect 11116 2912 11118 2964
rect 11118 2912 11170 2964
rect 11170 2912 11172 2964
rect 11116 2910 11172 2912
rect 11197 2964 11253 2966
rect 11197 2912 11199 2964
rect 11199 2912 11251 2964
rect 11251 2912 11253 2964
rect 11197 2910 11253 2912
rect 11278 2964 11334 2966
rect 11278 2912 11280 2964
rect 11280 2912 11332 2964
rect 11332 2912 11334 2964
rect 11278 2910 11334 2912
rect 11359 2964 11415 2966
rect 11359 2912 11361 2964
rect 11361 2912 11413 2964
rect 11413 2912 11415 2964
rect 11359 2910 11415 2912
rect 11440 2964 11496 2966
rect 11440 2912 11442 2964
rect 11442 2912 11494 2964
rect 11494 2912 11496 2964
rect 11440 2910 11496 2912
rect 11521 2964 11577 2966
rect 11521 2912 11523 2964
rect 11523 2912 11575 2964
rect 11575 2912 11577 2964
rect 11521 2910 11577 2912
rect 11602 2964 11658 2966
rect 11602 2912 11604 2964
rect 11604 2912 11656 2964
rect 11656 2912 11658 2964
rect 11602 2910 11658 2912
rect 11684 2964 11740 2966
rect 11684 2912 11686 2964
rect 11686 2912 11738 2964
rect 11738 2912 11740 2964
rect 11684 2910 11740 2912
rect 11765 2964 11821 2966
rect 11765 2912 11767 2964
rect 11767 2912 11819 2964
rect 11819 2912 11821 2964
rect 11765 2910 11821 2912
rect 11846 2964 11902 2966
rect 11846 2912 11848 2964
rect 11848 2912 11900 2964
rect 11900 2912 11902 2964
rect 11846 2910 11902 2912
rect 11927 2964 11983 2966
rect 11927 2912 11929 2964
rect 11929 2912 11981 2964
rect 11981 2912 11983 2964
rect 11927 2910 11983 2912
rect 12008 2964 12064 2966
rect 12008 2912 12010 2964
rect 12010 2912 12062 2964
rect 12062 2912 12064 2964
rect 12008 2910 12064 2912
rect 12089 2964 12145 2966
rect 12089 2912 12091 2964
rect 12091 2912 12143 2964
rect 12143 2912 12145 2964
rect 12089 2910 12145 2912
rect 12170 2964 12226 2966
rect 12170 2912 12172 2964
rect 12172 2912 12224 2964
rect 12224 2912 12226 2964
rect 12170 2910 12226 2912
rect 12252 2964 12308 2966
rect 12252 2912 12254 2964
rect 12254 2912 12306 2964
rect 12306 2912 12308 2964
rect 12252 2910 12308 2912
rect 12333 2964 12389 2966
rect 12333 2912 12335 2964
rect 12335 2912 12387 2964
rect 12387 2912 12389 2964
rect 12333 2910 12389 2912
rect 12414 2964 12470 2966
rect 12414 2912 12416 2964
rect 12416 2912 12468 2964
rect 12468 2912 12470 2964
rect 12414 2910 12470 2912
rect 12495 2964 12551 2966
rect 12495 2912 12497 2964
rect 12497 2912 12549 2964
rect 12549 2912 12551 2964
rect 12495 2910 12551 2912
rect 12576 2964 12632 2966
rect 12576 2912 12578 2964
rect 12578 2912 12630 2964
rect 12630 2912 12632 2964
rect 12576 2910 12632 2912
rect 12657 2964 12713 2966
rect 12657 2912 12659 2964
rect 12659 2912 12711 2964
rect 12711 2912 12713 2964
rect 12657 2910 12713 2912
rect 12738 2964 12794 2966
rect 12738 2912 12740 2964
rect 12740 2912 12792 2964
rect 12792 2912 12794 2964
rect 12738 2910 12794 2912
rect 12820 2964 12876 2966
rect 12820 2912 12822 2964
rect 12822 2912 12874 2964
rect 12874 2912 12876 2964
rect 12820 2910 12876 2912
rect 12901 2964 12957 2966
rect 12901 2912 12903 2964
rect 12903 2912 12955 2964
rect 12955 2912 12957 2964
rect 12901 2910 12957 2912
rect 12982 2964 13038 2966
rect 12982 2912 12984 2964
rect 12984 2912 13036 2964
rect 13036 2912 13038 2964
rect 12982 2910 13038 2912
rect 13063 2964 13119 2966
rect 13063 2912 13065 2964
rect 13065 2912 13117 2964
rect 13117 2912 13119 2964
rect 13063 2910 13119 2912
rect 13144 2964 13200 2966
rect 13144 2912 13146 2964
rect 13146 2912 13198 2964
rect 13198 2912 13200 2964
rect 13144 2910 13200 2912
rect 13225 2964 13281 2966
rect 13225 2912 13227 2964
rect 13227 2912 13279 2964
rect 13279 2912 13281 2964
rect 13225 2910 13281 2912
rect 13306 2964 13362 2966
rect 13306 2912 13308 2964
rect 13308 2912 13360 2964
rect 13360 2912 13362 2964
rect 13306 2910 13362 2912
rect 13388 2964 13444 2966
rect 13388 2912 13390 2964
rect 13390 2912 13442 2964
rect 13442 2912 13444 2964
rect 13388 2910 13444 2912
rect 13469 2964 13525 2966
rect 13469 2912 13471 2964
rect 13471 2912 13523 2964
rect 13523 2912 13525 2964
rect 13469 2910 13525 2912
rect 13550 2964 13606 2966
rect 13550 2912 13552 2964
rect 13552 2912 13604 2964
rect 13604 2912 13606 2964
rect 13550 2910 13606 2912
rect 13631 2964 13687 2966
rect 13631 2912 13633 2964
rect 13633 2912 13685 2964
rect 13685 2912 13687 2964
rect 13631 2910 13687 2912
rect 13712 2964 13768 2966
rect 13712 2912 13714 2964
rect 13714 2912 13766 2964
rect 13766 2912 13768 2964
rect 13712 2910 13768 2912
rect 13793 2964 13849 2966
rect 13793 2912 13795 2964
rect 13795 2912 13847 2964
rect 13847 2912 13849 2964
rect 13793 2910 13849 2912
rect 13874 2964 13930 2966
rect 13874 2912 13876 2964
rect 13876 2912 13928 2964
rect 13928 2912 13930 2964
rect 13874 2910 13930 2912
rect 13956 2964 14012 2966
rect 13956 2912 13958 2964
rect 13958 2912 14010 2964
rect 14010 2912 14012 2964
rect 13956 2910 14012 2912
rect 14037 2964 14093 2966
rect 14037 2912 14039 2964
rect 14039 2912 14091 2964
rect 14091 2912 14093 2964
rect 14037 2910 14093 2912
rect 14118 2964 14174 2966
rect 14118 2912 14120 2964
rect 14120 2912 14172 2964
rect 14172 2912 14174 2964
rect 14118 2910 14174 2912
rect 14199 2964 14255 2966
rect 14199 2912 14201 2964
rect 14201 2912 14253 2964
rect 14253 2912 14255 2964
rect 14199 2910 14255 2912
rect 14280 2964 14336 2966
rect 14280 2912 14282 2964
rect 14282 2912 14334 2964
rect 14334 2912 14336 2964
rect 14280 2910 14336 2912
rect 14361 2964 14417 2966
rect 14361 2912 14363 2964
rect 14363 2912 14415 2964
rect 14415 2912 14417 2964
rect 14361 2910 14417 2912
rect 14442 2964 14498 2966
rect 14442 2912 14444 2964
rect 14444 2912 14496 2964
rect 14496 2912 14498 2964
rect 14442 2910 14498 2912
rect 14524 2964 14580 2966
rect 14524 2912 14526 2964
rect 14526 2912 14578 2964
rect 14578 2912 14580 2964
rect 14524 2910 14580 2912
rect 14605 2964 14661 2966
rect 14605 2912 14607 2964
rect 14607 2912 14659 2964
rect 14659 2912 14661 2964
rect 14605 2910 14661 2912
rect 14686 2964 14742 2966
rect 14686 2912 14688 2964
rect 14688 2912 14740 2964
rect 14740 2912 14742 2964
rect 14686 2910 14742 2912
rect 14767 2964 14823 2966
rect 14767 2912 14769 2964
rect 14769 2912 14821 2964
rect 14821 2912 14823 2964
rect 14767 2910 14823 2912
rect 14848 2964 14904 2966
rect 14848 2912 14850 2964
rect 14850 2912 14902 2964
rect 14902 2912 14904 2964
rect 14848 2910 14904 2912
rect 14929 2964 14985 2966
rect 14929 2912 14931 2964
rect 14931 2912 14983 2964
rect 14983 2912 14985 2964
rect 14929 2910 14985 2912
rect 15010 2964 15066 2966
rect 15010 2912 15012 2964
rect 15012 2912 15064 2964
rect 15064 2912 15066 2964
rect 15010 2910 15066 2912
rect 15092 2964 15148 2966
rect 15092 2912 15094 2964
rect 15094 2912 15146 2964
rect 15146 2912 15148 2964
rect 15092 2910 15148 2912
rect 15173 2964 15229 2966
rect 15173 2912 15175 2964
rect 15175 2912 15227 2964
rect 15227 2912 15229 2964
rect 15173 2910 15229 2912
rect 15254 2964 15310 2966
rect 15254 2912 15256 2964
rect 15256 2912 15308 2964
rect 15308 2912 15310 2964
rect 15254 2910 15310 2912
rect 15335 2964 15391 2966
rect 15335 2912 15337 2964
rect 15337 2912 15389 2964
rect 15389 2912 15391 2964
rect 15335 2910 15391 2912
rect 15416 2964 15472 2966
rect 15416 2912 15418 2964
rect 15418 2912 15470 2964
rect 15470 2912 15472 2964
rect 15416 2910 15472 2912
rect 15497 2964 15553 2966
rect 15497 2912 15499 2964
rect 15499 2912 15551 2964
rect 15551 2912 15553 2964
rect 15497 2910 15553 2912
rect 15578 2964 15634 2966
rect 15578 2912 15580 2964
rect 15580 2912 15632 2964
rect 15632 2912 15634 2964
rect 15578 2910 15634 2912
rect 15660 2964 15716 2966
rect 15660 2912 15662 2964
rect 15662 2912 15714 2964
rect 15714 2912 15716 2964
rect 15660 2910 15716 2912
rect 15741 2964 15797 2966
rect 15741 2912 15743 2964
rect 15743 2912 15795 2964
rect 15795 2912 15797 2964
rect 15741 2910 15797 2912
rect 15822 2964 15878 2966
rect 15822 2912 15824 2964
rect 15824 2912 15876 2964
rect 15876 2912 15878 2964
rect 15822 2910 15878 2912
rect 15903 2964 15959 2966
rect 15903 2912 15905 2964
rect 15905 2912 15957 2964
rect 15957 2912 15959 2964
rect 15903 2910 15959 2912
rect 15984 2964 16040 2966
rect 15984 2912 15986 2964
rect 15986 2912 16038 2964
rect 16038 2912 16040 2964
rect 15984 2910 16040 2912
rect 16065 2964 16121 2966
rect 16065 2912 16067 2964
rect 16067 2912 16119 2964
rect 16119 2912 16121 2964
rect 16065 2910 16121 2912
rect 16146 2964 16202 2966
rect 16146 2912 16148 2964
rect 16148 2912 16200 2964
rect 16200 2912 16202 2964
rect 16146 2910 16202 2912
rect 16228 2964 16284 2966
rect 16228 2912 16230 2964
rect 16230 2912 16282 2964
rect 16282 2912 16284 2964
rect 16228 2910 16284 2912
rect 16309 2964 16365 2966
rect 16309 2912 16311 2964
rect 16311 2912 16363 2964
rect 16363 2912 16365 2964
rect 16309 2910 16365 2912
rect 16390 2964 16446 2966
rect 16390 2912 16392 2964
rect 16392 2912 16444 2964
rect 16444 2912 16446 2964
rect 16390 2910 16446 2912
rect 16471 2964 16527 2966
rect 16471 2912 16473 2964
rect 16473 2912 16525 2964
rect 16525 2912 16527 2964
rect 16471 2910 16527 2912
rect 16552 2964 16608 2966
rect 16552 2912 16554 2964
rect 16554 2912 16606 2964
rect 16606 2912 16608 2964
rect 16552 2910 16608 2912
rect 16633 2964 16689 2966
rect 16633 2912 16635 2964
rect 16635 2912 16687 2964
rect 16687 2912 16689 2964
rect 16633 2910 16689 2912
rect 16714 2964 16770 2966
rect 16714 2912 16716 2964
rect 16716 2912 16768 2964
rect 16768 2912 16770 2964
rect 16714 2910 16770 2912
rect 16796 2964 16852 2966
rect 16796 2912 16798 2964
rect 16798 2912 16850 2964
rect 16850 2912 16852 2964
rect 16796 2910 16852 2912
rect 16877 2964 16933 2966
rect 16877 2912 16879 2964
rect 16879 2912 16931 2964
rect 16931 2912 16933 2964
rect 16877 2910 16933 2912
rect 16958 2964 17014 2966
rect 16958 2912 16960 2964
rect 16960 2912 17012 2964
rect 17012 2912 17014 2964
rect 16958 2910 17014 2912
rect 17039 2964 17095 2966
rect 17039 2912 17041 2964
rect 17041 2912 17093 2964
rect 17093 2912 17095 2964
rect 17039 2910 17095 2912
rect 17120 2964 17176 2966
rect 17120 2912 17122 2964
rect 17122 2912 17174 2964
rect 17174 2912 17176 2964
rect 17120 2910 17176 2912
rect 17201 2964 17257 2966
rect 17201 2912 17203 2964
rect 17203 2912 17255 2964
rect 17255 2912 17257 2964
rect 17201 2910 17257 2912
rect 17282 2964 17338 2966
rect 17282 2912 17284 2964
rect 17284 2912 17336 2964
rect 17336 2912 17338 2964
rect 17282 2910 17338 2912
rect 17364 2964 17420 2966
rect 17364 2912 17366 2964
rect 17366 2912 17418 2964
rect 17418 2912 17420 2964
rect 17364 2910 17420 2912
rect 17445 2964 17501 2966
rect 17445 2912 17447 2964
rect 17447 2912 17499 2964
rect 17499 2912 17501 2964
rect 17445 2910 17501 2912
rect 17526 2964 17582 2966
rect 17526 2912 17528 2964
rect 17528 2912 17580 2964
rect 17580 2912 17582 2964
rect 17526 2910 17582 2912
rect 17607 2964 17663 2966
rect 17607 2912 17609 2964
rect 17609 2912 17661 2964
rect 17661 2912 17663 2964
rect 17607 2910 17663 2912
rect 17688 2964 17744 2966
rect 17688 2912 17690 2964
rect 17690 2912 17742 2964
rect 17742 2912 17744 2964
rect 17688 2910 17744 2912
rect 17769 2964 17825 2966
rect 17769 2912 17771 2964
rect 17771 2912 17823 2964
rect 17823 2912 17825 2964
rect 17769 2910 17825 2912
rect 17850 2964 17906 2966
rect 17850 2912 17852 2964
rect 17852 2912 17904 2964
rect 17904 2912 17906 2964
rect 17850 2910 17906 2912
rect 17932 2964 17988 2966
rect 17932 2912 17934 2964
rect 17934 2912 17986 2964
rect 17986 2912 17988 2964
rect 17932 2910 17988 2912
rect 18013 2964 18069 2966
rect 18013 2912 18015 2964
rect 18015 2912 18067 2964
rect 18067 2912 18069 2964
rect 18013 2910 18069 2912
rect 18094 2964 18150 2966
rect 18094 2912 18096 2964
rect 18096 2912 18148 2964
rect 18148 2912 18150 2964
rect 18094 2910 18150 2912
rect 18175 2964 18231 2966
rect 18175 2912 18177 2964
rect 18177 2912 18229 2964
rect 18229 2912 18231 2964
rect 18175 2910 18231 2912
rect 18256 2964 18312 2966
rect 18256 2912 18258 2964
rect 18258 2912 18310 2964
rect 18310 2912 18312 2964
rect 18256 2910 18312 2912
rect 18337 2964 18393 2966
rect 18337 2912 18339 2964
rect 18339 2912 18391 2964
rect 18391 2912 18393 2964
rect 18337 2910 18393 2912
rect 18418 2964 18474 2966
rect 18418 2912 18420 2964
rect 18420 2912 18472 2964
rect 18472 2912 18474 2964
rect 18418 2910 18474 2912
rect 18500 2964 18556 2966
rect 18500 2912 18502 2964
rect 18502 2912 18554 2964
rect 18554 2912 18556 2964
rect 18500 2910 18556 2912
rect 18581 2964 18637 2966
rect 18581 2912 18583 2964
rect 18583 2912 18635 2964
rect 18635 2912 18637 2964
rect 18581 2910 18637 2912
rect 18662 2964 18718 2966
rect 18662 2912 18664 2964
rect 18664 2912 18716 2964
rect 18716 2912 18718 2964
rect 18662 2910 18718 2912
rect 18743 2964 18799 2966
rect 18743 2912 18745 2964
rect 18745 2912 18797 2964
rect 18797 2912 18799 2964
rect 18743 2910 18799 2912
rect 18824 2964 18880 2966
rect 18824 2912 18826 2964
rect 18826 2912 18878 2964
rect 18878 2912 18880 2964
rect 18824 2910 18880 2912
rect 18905 2964 18961 2966
rect 18905 2912 18907 2964
rect 18907 2912 18959 2964
rect 18959 2912 18961 2964
rect 18905 2910 18961 2912
rect 18986 2964 19042 2966
rect 18986 2912 18988 2964
rect 18988 2912 19040 2964
rect 19040 2912 19042 2964
rect 18986 2910 19042 2912
rect 19068 2964 19124 2966
rect 19068 2912 19070 2964
rect 19070 2912 19122 2964
rect 19122 2912 19124 2964
rect 19068 2910 19124 2912
rect 19149 2964 19205 2966
rect 19149 2912 19151 2964
rect 19151 2912 19203 2964
rect 19203 2912 19205 2964
rect 19149 2910 19205 2912
rect 19230 2964 19286 2966
rect 19230 2912 19232 2964
rect 19232 2912 19284 2964
rect 19284 2912 19286 2964
rect 19230 2910 19286 2912
rect 19311 2964 19367 2966
rect 19311 2912 19313 2964
rect 19313 2912 19365 2964
rect 19365 2912 19367 2964
rect 19311 2910 19367 2912
rect 19392 2964 19448 2966
rect 19392 2912 19394 2964
rect 19394 2912 19446 2964
rect 19446 2912 19448 2964
rect 19392 2910 19448 2912
rect 19473 2964 19529 2966
rect 19473 2912 19475 2964
rect 19475 2912 19527 2964
rect 19527 2912 19529 2964
rect 19473 2910 19529 2912
rect 19554 2964 19610 2966
rect 19554 2912 19556 2964
rect 19556 2912 19608 2964
rect 19608 2912 19610 2964
rect 19554 2910 19610 2912
rect 19636 2964 19692 2966
rect 19636 2912 19638 2964
rect 19638 2912 19690 2964
rect 19690 2912 19692 2964
rect 19636 2910 19692 2912
rect 19717 2964 19773 2966
rect 19717 2912 19719 2964
rect 19719 2912 19771 2964
rect 19771 2912 19773 2964
rect 19717 2910 19773 2912
rect 19798 2964 19854 2966
rect 19798 2912 19800 2964
rect 19800 2912 19852 2964
rect 19852 2912 19854 2964
rect 19798 2910 19854 2912
rect 19879 2964 19935 2966
rect 19879 2912 19881 2964
rect 19881 2912 19933 2964
rect 19933 2912 19935 2964
rect 19879 2910 19935 2912
rect 19960 2964 20016 2966
rect 19960 2912 19962 2964
rect 19962 2912 20014 2964
rect 20014 2912 20016 2964
rect 19960 2910 20016 2912
rect 20041 2964 20097 2966
rect 20041 2912 20043 2964
rect 20043 2912 20095 2964
rect 20095 2912 20097 2964
rect 20041 2910 20097 2912
rect 20122 2964 20178 2966
rect 20122 2912 20124 2964
rect 20124 2912 20176 2964
rect 20176 2912 20178 2964
rect 20122 2910 20178 2912
rect 20204 2964 20260 2966
rect 20204 2912 20206 2964
rect 20206 2912 20258 2964
rect 20258 2912 20260 2964
rect 20204 2910 20260 2912
rect 20285 2964 20341 2966
rect 20285 2912 20287 2964
rect 20287 2912 20339 2964
rect 20339 2912 20341 2964
rect 20285 2910 20341 2912
rect 20366 2964 20422 2966
rect 20366 2912 20368 2964
rect 20368 2912 20420 2964
rect 20420 2912 20422 2964
rect 20366 2910 20422 2912
rect 20447 2964 20503 2966
rect 20447 2912 20449 2964
rect 20449 2912 20501 2964
rect 20501 2912 20503 2964
rect 20447 2910 20503 2912
rect 20528 2964 20584 2966
rect 20528 2912 20530 2964
rect 20530 2912 20582 2964
rect 20582 2912 20584 2964
rect 20528 2910 20584 2912
rect 20609 2964 20665 2966
rect 20609 2912 20611 2964
rect 20611 2912 20663 2964
rect 20663 2912 20665 2964
rect 20609 2910 20665 2912
rect 20690 2964 20746 2966
rect 20690 2912 20692 2964
rect 20692 2912 20744 2964
rect 20744 2912 20746 2964
rect 20690 2910 20746 2912
rect 20772 2964 20828 2966
rect 20772 2912 20774 2964
rect 20774 2912 20826 2964
rect 20826 2912 20828 2964
rect 20772 2910 20828 2912
rect 20853 2964 20909 2966
rect 20853 2912 20855 2964
rect 20855 2912 20907 2964
rect 20907 2912 20909 2964
rect 20853 2910 20909 2912
rect 20934 2964 20990 2966
rect 20934 2912 20936 2964
rect 20936 2912 20988 2964
rect 20988 2912 20990 2964
rect 20934 2910 20990 2912
rect 21015 2964 21071 2966
rect 21015 2912 21017 2964
rect 21017 2912 21069 2964
rect 21069 2912 21071 2964
rect 21015 2910 21071 2912
rect 21096 2964 21152 2966
rect 21096 2912 21098 2964
rect 21098 2912 21150 2964
rect 21150 2912 21152 2964
rect 21096 2910 21152 2912
rect 21177 2964 21233 2966
rect 21177 2912 21179 2964
rect 21179 2912 21231 2964
rect 21231 2912 21233 2964
rect 21177 2910 21233 2912
rect 21258 2964 21314 2966
rect 21258 2912 21260 2964
rect 21260 2912 21312 2964
rect 21312 2912 21314 2964
rect 21258 2910 21314 2912
rect 21340 2964 21396 2966
rect 21340 2912 21342 2964
rect 21342 2912 21394 2964
rect 21394 2912 21396 2964
rect 21340 2910 21396 2912
rect 21421 2964 21477 2966
rect 21421 2912 21423 2964
rect 21423 2912 21475 2964
rect 21475 2912 21477 2964
rect 21421 2910 21477 2912
rect 21502 2964 21558 2966
rect 21502 2912 21504 2964
rect 21504 2912 21556 2964
rect 21556 2912 21558 2964
rect 21502 2910 21558 2912
rect 21583 2964 21639 2966
rect 21583 2912 21585 2964
rect 21585 2912 21637 2964
rect 21637 2912 21639 2964
rect 21583 2910 21639 2912
rect 21664 2964 21720 2966
rect 21664 2912 21666 2964
rect 21666 2912 21718 2964
rect 21718 2912 21720 2964
rect 21664 2910 21720 2912
rect 21745 2964 21801 2966
rect 21745 2912 21747 2964
rect 21747 2912 21799 2964
rect 21799 2912 21801 2964
rect 21745 2910 21801 2912
rect 21826 2964 21882 2966
rect 21826 2912 21828 2964
rect 21828 2912 21880 2964
rect 21880 2912 21882 2964
rect 21826 2910 21882 2912
rect 21908 2964 21964 2966
rect 21908 2912 21910 2964
rect 21910 2912 21962 2964
rect 21962 2912 21964 2964
rect 21908 2910 21964 2912
rect 21989 2964 22045 2966
rect 21989 2912 21991 2964
rect 21991 2912 22043 2964
rect 22043 2912 22045 2964
rect 21989 2910 22045 2912
rect 22070 2964 22126 2966
rect 22070 2912 22072 2964
rect 22072 2912 22124 2964
rect 22124 2912 22126 2964
rect 22070 2910 22126 2912
rect 22151 2964 22207 2966
rect 22151 2912 22153 2964
rect 22153 2912 22205 2964
rect 22205 2912 22207 2964
rect 22151 2910 22207 2912
rect 22232 2964 22288 2966
rect 22232 2912 22234 2964
rect 22234 2912 22286 2964
rect 22286 2912 22288 2964
rect 22232 2910 22288 2912
rect 22313 2964 22369 2966
rect 22313 2912 22315 2964
rect 22315 2912 22367 2964
rect 22367 2912 22369 2964
rect 22313 2910 22369 2912
rect 22394 2964 22450 2966
rect 22394 2912 22396 2964
rect 22396 2912 22448 2964
rect 22448 2912 22450 2964
rect 22394 2910 22450 2912
rect 22476 2964 22532 2966
rect 22476 2912 22478 2964
rect 22478 2912 22530 2964
rect 22530 2912 22532 2964
rect 22476 2910 22532 2912
rect 22557 2964 22613 2966
rect 22557 2912 22559 2964
rect 22559 2912 22611 2964
rect 22611 2912 22613 2964
rect 22557 2910 22613 2912
rect 22638 2964 22694 2966
rect 22638 2912 22640 2964
rect 22640 2912 22692 2964
rect 22692 2912 22694 2964
rect 22638 2910 22694 2912
rect 22719 2964 22775 2966
rect 22719 2912 22721 2964
rect 22721 2912 22773 2964
rect 22773 2912 22775 2964
rect 22719 2910 22775 2912
rect 22800 2964 22856 2966
rect 22800 2912 22802 2964
rect 22802 2912 22854 2964
rect 22854 2912 22856 2964
rect 22800 2910 22856 2912
rect 22881 2964 22937 2966
rect 22881 2912 22883 2964
rect 22883 2912 22935 2964
rect 22935 2912 22937 2964
rect 22881 2910 22937 2912
rect 22962 2964 23018 2966
rect 22962 2912 22964 2964
rect 22964 2912 23016 2964
rect 23016 2912 23018 2964
rect 22962 2910 23018 2912
rect 23044 2964 23100 2966
rect 23044 2912 23046 2964
rect 23046 2912 23098 2964
rect 23098 2912 23100 2964
rect 23044 2910 23100 2912
rect 23125 2964 23181 2966
rect 23125 2912 23127 2964
rect 23127 2912 23179 2964
rect 23179 2912 23181 2964
rect 23125 2910 23181 2912
rect 23206 2964 23262 2966
rect 23206 2912 23208 2964
rect 23208 2912 23260 2964
rect 23260 2912 23262 2964
rect 23206 2910 23262 2912
rect 23287 2964 23343 2966
rect 23287 2912 23289 2964
rect 23289 2912 23341 2964
rect 23341 2912 23343 2964
rect 23287 2910 23343 2912
rect 23368 2964 23424 2966
rect 23368 2912 23370 2964
rect 23370 2912 23422 2964
rect 23422 2912 23424 2964
rect 23368 2910 23424 2912
rect 23449 2964 23505 2966
rect 23449 2912 23451 2964
rect 23451 2912 23503 2964
rect 23503 2912 23505 2964
rect 23449 2910 23505 2912
rect 23530 2964 23586 2966
rect 23530 2912 23532 2964
rect 23532 2912 23584 2964
rect 23584 2912 23586 2964
rect 23530 2910 23586 2912
rect 23612 2964 23668 2966
rect 23612 2912 23614 2964
rect 23614 2912 23666 2964
rect 23666 2912 23668 2964
rect 23612 2910 23668 2912
rect 23693 2964 23749 2966
rect 23693 2912 23695 2964
rect 23695 2912 23747 2964
rect 23747 2912 23749 2964
rect 23693 2910 23749 2912
rect 23774 2964 23830 2966
rect 23774 2912 23776 2964
rect 23776 2912 23828 2964
rect 23828 2912 23830 2964
rect 23774 2910 23830 2912
rect 23855 2964 23911 2966
rect 23855 2912 23857 2964
rect 23857 2912 23909 2964
rect 23909 2912 23911 2964
rect 23855 2910 23911 2912
rect 23936 2964 23992 2966
rect 23936 2912 23938 2964
rect 23938 2912 23990 2964
rect 23990 2912 23992 2964
rect 23936 2910 23992 2912
rect 24017 2964 24073 2966
rect 24017 2912 24019 2964
rect 24019 2912 24071 2964
rect 24071 2912 24073 2964
rect 24017 2910 24073 2912
rect 24098 2964 24154 2966
rect 24098 2912 24100 2964
rect 24100 2912 24152 2964
rect 24152 2912 24154 2964
rect 24098 2910 24154 2912
rect 24180 2964 24236 2966
rect 24180 2912 24182 2964
rect 24182 2912 24234 2964
rect 24234 2912 24236 2964
rect 24180 2910 24236 2912
rect 24261 2964 24317 2966
rect 24261 2912 24263 2964
rect 24263 2912 24315 2964
rect 24315 2912 24317 2964
rect 24261 2910 24317 2912
rect 24342 2964 24398 2966
rect 24342 2912 24344 2964
rect 24344 2912 24396 2964
rect 24396 2912 24398 2964
rect 24342 2910 24398 2912
rect 24423 2964 24479 2966
rect 24423 2912 24425 2964
rect 24425 2912 24477 2964
rect 24477 2912 24479 2964
rect 24423 2910 24479 2912
rect 24504 2964 24560 2966
rect 24504 2912 24506 2964
rect 24506 2912 24558 2964
rect 24558 2912 24560 2964
rect 24504 2910 24560 2912
rect 24585 2964 24641 2966
rect 24585 2912 24587 2964
rect 24587 2912 24639 2964
rect 24639 2912 24641 2964
rect 24585 2910 24641 2912
rect 24666 2964 24722 2966
rect 24666 2912 24668 2964
rect 24668 2912 24720 2964
rect 24720 2912 24722 2964
rect 24666 2910 24722 2912
rect 6915 2107 6917 2667
rect 6917 2107 6969 2667
rect 6969 2107 6971 2667
rect 7151 2107 7153 2667
rect 7153 2107 7205 2667
rect 7205 2107 7207 2667
rect 7387 2107 7389 2667
rect 7389 2107 7441 2667
rect 7441 2107 7443 2667
rect 7623 2107 7625 2667
rect 7625 2107 7677 2667
rect 7677 2107 7679 2667
rect 7859 2107 7861 2667
rect 7861 2107 7913 2667
rect 7913 2107 7915 2667
rect 8095 2107 8097 2667
rect 8097 2107 8149 2667
rect 8149 2107 8151 2667
rect 8331 2107 8333 2667
rect 8333 2107 8385 2667
rect 8385 2107 8387 2667
rect 8567 2107 8569 2667
rect 8569 2107 8621 2667
rect 8621 2107 8623 2667
rect 8913 2107 8915 2667
rect 8915 2107 8967 2667
rect 8967 2107 8969 2667
rect 9149 2107 9151 2667
rect 9151 2107 9203 2667
rect 9203 2107 9205 2667
rect 9385 2107 9387 2667
rect 9387 2107 9439 2667
rect 9439 2107 9441 2667
rect 9621 2107 9623 2667
rect 9623 2107 9675 2667
rect 9675 2107 9677 2667
rect 9857 2107 9859 2667
rect 9859 2107 9911 2667
rect 9911 2107 9913 2667
rect 10093 2107 10095 2667
rect 10095 2107 10147 2667
rect 10147 2107 10149 2667
rect 10329 2107 10331 2667
rect 10331 2107 10383 2667
rect 10383 2107 10385 2667
rect 10565 2107 10567 2667
rect 10567 2107 10619 2667
rect 10619 2107 10621 2667
rect 12607 2106 12609 2666
rect 12609 2106 12661 2666
rect 12661 2106 12663 2666
rect 12843 2106 12845 2666
rect 12845 2106 12897 2666
rect 12897 2106 12899 2666
rect 13079 2106 13081 2666
rect 13081 2106 13133 2666
rect 13133 2106 13135 2666
rect 13315 2106 13317 2666
rect 13317 2106 13369 2666
rect 13369 2106 13371 2666
rect 13551 2106 13553 2666
rect 13553 2106 13605 2666
rect 13605 2106 13607 2666
rect 13787 2106 13789 2666
rect 13789 2106 13841 2666
rect 13841 2106 13843 2666
rect 14023 2106 14025 2666
rect 14025 2106 14077 2666
rect 14077 2106 14079 2666
rect 14259 2106 14261 2666
rect 14261 2106 14313 2666
rect 14313 2106 14315 2666
rect 14495 2106 14497 2666
rect 14497 2106 14549 2666
rect 14549 2106 14551 2666
rect 14731 2106 14733 2666
rect 14733 2106 14785 2666
rect 14785 2106 14787 2666
rect 14967 2106 14969 2666
rect 14969 2106 15021 2666
rect 15021 2106 15023 2666
rect 15203 2106 15205 2666
rect 15205 2106 15257 2666
rect 15257 2106 15259 2666
rect 15439 2106 15441 2666
rect 15441 2106 15493 2666
rect 15493 2106 15495 2666
rect 16730 2106 16732 2666
rect 16732 2106 16784 2666
rect 16784 2106 16786 2666
rect 16966 2106 16968 2666
rect 16968 2106 17020 2666
rect 17020 2106 17022 2666
rect 17202 2106 17204 2666
rect 17204 2106 17256 2666
rect 17256 2106 17258 2666
rect 17438 2106 17440 2666
rect 17440 2106 17492 2666
rect 17492 2106 17494 2666
rect 17674 2106 17676 2666
rect 17676 2106 17728 2666
rect 17728 2106 17730 2666
rect 17910 2106 17912 2666
rect 17912 2106 17964 2666
rect 17964 2106 17966 2666
rect 18146 2106 18148 2666
rect 18148 2106 18200 2666
rect 18200 2106 18202 2666
rect 18382 2106 18384 2666
rect 18384 2106 18436 2666
rect 18436 2106 18438 2666
rect 18618 2106 18620 2666
rect 18620 2106 18672 2666
rect 18672 2106 18674 2666
rect 18854 2106 18856 2666
rect 18856 2106 18908 2666
rect 18908 2106 18910 2666
rect 19090 2106 19092 2666
rect 19092 2106 19144 2666
rect 19144 2106 19146 2666
rect 19326 2106 19328 2666
rect 19328 2106 19380 2666
rect 19380 2106 19382 2666
rect 19562 2106 19564 2666
rect 19564 2106 19616 2666
rect 19616 2106 19618 2666
rect 20853 2106 20855 2666
rect 20855 2106 20907 2666
rect 20907 2106 20909 2666
rect 21089 2106 21091 2666
rect 21091 2106 21143 2666
rect 21143 2106 21145 2666
rect 21325 2106 21327 2666
rect 21327 2106 21379 2666
rect 21379 2106 21381 2666
rect 21561 2106 21563 2666
rect 21563 2106 21615 2666
rect 21615 2106 21617 2666
rect 21797 2106 21799 2666
rect 21799 2106 21851 2666
rect 21851 2106 21853 2666
rect 22033 2106 22035 2666
rect 22035 2106 22087 2666
rect 22087 2106 22089 2666
rect 22269 2106 22271 2666
rect 22271 2106 22323 2666
rect 22323 2106 22325 2666
rect 22505 2106 22507 2666
rect 22507 2106 22559 2666
rect 22559 2106 22561 2666
rect 22741 2106 22743 2666
rect 22743 2106 22795 2666
rect 22795 2106 22797 2666
rect 22977 2106 22979 2666
rect 22979 2106 23031 2666
rect 23031 2106 23033 2666
rect 23213 2106 23215 2666
rect 23215 2106 23267 2666
rect 23267 2106 23269 2666
rect 23449 2106 23451 2666
rect 23451 2106 23503 2666
rect 23503 2106 23505 2666
rect 23685 2106 23687 2666
rect 23687 2106 23739 2666
rect 23739 2106 23741 2666
rect 4775 1569 4831 1593
rect 4775 1537 4801 1569
rect 4801 1537 4831 1569
rect 4856 1537 4912 1593
rect 4937 1537 4993 1593
rect 5018 1569 5074 1593
rect 5018 1537 5037 1569
rect 5037 1537 5074 1569
rect 5099 1537 5155 1593
rect 5180 1537 5236 1593
rect 5261 1569 5317 1593
rect 5261 1537 5273 1569
rect 5273 1537 5317 1569
rect 5363 1537 5419 1593
rect 5444 1537 5500 1593
rect 5525 1569 5581 1593
rect 5525 1537 5561 1569
rect 5561 1537 5581 1569
rect 5606 1537 5662 1593
rect 5687 1537 5743 1593
rect 5768 1569 5824 1593
rect 5768 1537 5797 1569
rect 5797 1537 5824 1569
rect 5849 1537 5905 1593
rect 5951 1569 6007 1593
rect 6032 1569 6088 1593
rect 5951 1537 5981 1569
rect 5981 1537 6007 1569
rect 6032 1537 6033 1569
rect 6033 1537 6088 1569
rect 6113 1537 6169 1593
rect 6194 1569 6250 1593
rect 6194 1537 6217 1569
rect 6217 1537 6250 1569
rect 6275 1537 6331 1593
rect 6356 1537 6412 1593
rect 6437 1569 6493 1593
rect 6437 1537 6453 1569
rect 6453 1537 6493 1569
rect 6517 1537 6573 1593
rect 6598 1537 6654 1593
rect 6679 1569 6735 1593
rect 6679 1537 6689 1569
rect 6689 1537 6735 1569
rect 6760 1537 6816 1593
rect 6841 1537 6897 1593
rect 6922 1569 6978 1593
rect 6922 1537 6925 1569
rect 6925 1537 6977 1569
rect 6977 1537 6978 1569
rect 7003 1537 7059 1593
rect 7090 1537 7146 1593
rect 7171 1569 7227 1593
rect 7171 1537 7213 1569
rect 7213 1537 7227 1569
rect 7252 1537 7308 1593
rect 7333 1537 7389 1593
rect 7414 1569 7470 1593
rect 7414 1537 7449 1569
rect 7449 1537 7470 1569
rect 7495 1537 7551 1593
rect 7576 1537 7632 1593
rect 7656 1569 7712 1593
rect 7656 1537 7685 1569
rect 7685 1537 7712 1569
rect 7737 1537 7793 1593
rect 7818 1569 7874 1593
rect 7899 1569 7955 1593
rect 7818 1537 7869 1569
rect 7869 1537 7874 1569
rect 7899 1537 7921 1569
rect 7921 1537 7955 1569
rect 7980 1537 8036 1593
rect 8061 1569 8117 1593
rect 8142 1569 8198 1593
rect 8061 1537 8105 1569
rect 8105 1537 8117 1569
rect 8142 1537 8157 1569
rect 8157 1537 8198 1569
rect 8222 1537 8278 1593
rect 8303 1569 8359 1593
rect 8384 1569 8440 1593
rect 8303 1537 8341 1569
rect 8341 1537 8359 1569
rect 8384 1537 8393 1569
rect 8393 1537 8440 1569
rect 8465 1537 8521 1593
rect 8546 1569 8602 1593
rect 8627 1569 8683 1593
rect 8546 1537 8577 1569
rect 8577 1537 8602 1569
rect 8627 1537 8629 1569
rect 8629 1537 8683 1569
rect 8708 1537 8764 1593
rect 8788 1569 8844 1593
rect 8788 1537 8813 1569
rect 8813 1537 8844 1569
rect 8869 1537 8925 1593
rect 8950 1537 9006 1593
rect 9031 1569 9087 1593
rect 9031 1537 9049 1569
rect 9049 1537 9087 1569
rect 9112 1537 9168 1593
rect 9193 1537 9249 1593
rect 9274 1569 9330 1593
rect 9274 1537 9285 1569
rect 9285 1537 9330 1569
rect 9357 1537 9413 1593
rect 9438 1537 9494 1593
rect 9519 1569 9575 1593
rect 9519 1537 9521 1569
rect 9521 1537 9573 1569
rect 9573 1537 9575 1569
rect 9600 1537 9656 1593
rect 9681 1537 9737 1593
rect 9762 1569 9818 1593
rect 9762 1537 9809 1569
rect 9809 1537 9818 1569
rect 9843 1537 9899 1593
rect 9923 1537 9979 1593
rect 10004 1569 10060 1593
rect 10004 1537 10045 1569
rect 10045 1537 10060 1569
rect 10085 1537 10141 1593
rect 10166 1537 10222 1593
rect 10247 1569 10303 1593
rect 10247 1537 10281 1569
rect 10281 1537 10303 1569
rect 10328 1537 10384 1593
rect 10409 1537 10465 1593
rect 10489 1569 10545 1593
rect 10489 1537 10517 1569
rect 10517 1537 10545 1569
rect 10570 1537 10626 1593
rect 10651 1569 10707 1593
rect 10732 1569 10788 1593
rect 10651 1537 10701 1569
rect 10701 1537 10707 1569
rect 10732 1537 10753 1569
rect 10753 1537 10788 1569
rect 10813 1537 10869 1593
rect 10894 1537 10950 1593
rect 10975 1537 11031 1593
rect 11055 1537 11111 1593
rect 11136 1537 11192 1593
rect 11217 1537 11273 1593
rect 11298 1537 11354 1593
rect 11379 1537 11435 1593
rect 11460 1537 11516 1593
rect 11541 1537 11597 1593
rect 4775 1433 4801 1489
rect 4801 1433 4831 1489
rect 4856 1433 4912 1489
rect 4937 1433 4993 1489
rect 5018 1433 5037 1489
rect 5037 1433 5074 1489
rect 5099 1433 5155 1489
rect 5180 1433 5236 1489
rect 5261 1433 5273 1489
rect 5273 1433 5317 1489
rect 5363 1433 5419 1489
rect 5444 1433 5500 1489
rect 5525 1433 5561 1489
rect 5561 1433 5581 1489
rect 5606 1433 5662 1489
rect 5687 1433 5743 1489
rect 5768 1433 5797 1489
rect 5797 1433 5824 1489
rect 5849 1433 5905 1489
rect 5951 1433 5981 1489
rect 5981 1433 6007 1489
rect 6032 1433 6033 1489
rect 6033 1433 6088 1489
rect 6113 1433 6169 1489
rect 6194 1433 6217 1489
rect 6217 1433 6250 1489
rect 6275 1433 6331 1489
rect 6356 1433 6412 1489
rect 6437 1433 6453 1489
rect 6453 1433 6493 1489
rect 6517 1433 6573 1489
rect 6598 1433 6654 1489
rect 6679 1433 6689 1489
rect 6689 1433 6735 1489
rect 6760 1433 6816 1489
rect 6841 1433 6897 1489
rect 6922 1433 6925 1489
rect 6925 1433 6977 1489
rect 6977 1433 6978 1489
rect 7003 1433 7059 1489
rect 7090 1433 7146 1489
rect 7171 1433 7213 1489
rect 7213 1433 7227 1489
rect 7252 1433 7308 1489
rect 7333 1433 7389 1489
rect 7414 1433 7449 1489
rect 7449 1433 7470 1489
rect 7495 1433 7551 1489
rect 7576 1433 7632 1489
rect 7656 1433 7685 1489
rect 7685 1433 7712 1489
rect 7737 1433 7793 1489
rect 7818 1433 7869 1489
rect 7869 1433 7874 1489
rect 7899 1433 7921 1489
rect 7921 1433 7955 1489
rect 7980 1433 8036 1489
rect 8061 1433 8105 1489
rect 8105 1433 8117 1489
rect 8142 1433 8157 1489
rect 8157 1433 8198 1489
rect 8222 1433 8278 1489
rect 8303 1433 8341 1489
rect 8341 1433 8359 1489
rect 8384 1433 8393 1489
rect 8393 1433 8440 1489
rect 8465 1433 8521 1489
rect 8546 1433 8577 1489
rect 8577 1433 8602 1489
rect 8627 1433 8629 1489
rect 8629 1433 8683 1489
rect 8708 1433 8764 1489
rect 8788 1433 8813 1489
rect 8813 1433 8844 1489
rect 8869 1433 8925 1489
rect 8950 1433 9006 1489
rect 9031 1433 9049 1489
rect 9049 1433 9087 1489
rect 9112 1433 9168 1489
rect 9193 1433 9249 1489
rect 9274 1433 9285 1489
rect 9285 1433 9330 1489
rect 9357 1433 9413 1489
rect 9438 1433 9494 1489
rect 9519 1433 9521 1489
rect 9521 1433 9573 1489
rect 9573 1433 9575 1489
rect 9600 1433 9656 1489
rect 9681 1433 9737 1489
rect 9762 1433 9809 1489
rect 9809 1433 9818 1489
rect 9843 1433 9899 1489
rect 9923 1433 9979 1489
rect 10004 1433 10045 1489
rect 10045 1433 10060 1489
rect 10085 1433 10141 1489
rect 10166 1433 10222 1489
rect 10247 1433 10281 1489
rect 10281 1433 10303 1489
rect 10328 1433 10384 1489
rect 10409 1433 10465 1489
rect 10489 1433 10517 1489
rect 10517 1433 10545 1489
rect 10570 1433 10626 1489
rect 10651 1433 10701 1489
rect 10701 1433 10707 1489
rect 10732 1433 10753 1489
rect 10753 1433 10788 1489
rect 10813 1433 10869 1489
rect 10894 1433 10950 1489
rect 10975 1433 11031 1489
rect 11055 1433 11111 1489
rect 11136 1433 11192 1489
rect 11217 1433 11273 1489
rect 11298 1433 11354 1489
rect 11379 1433 11435 1489
rect 11460 1433 11516 1489
rect 11541 1433 11597 1489
rect 4775 1329 4801 1385
rect 4801 1329 4831 1385
rect 4856 1329 4912 1385
rect 4937 1329 4993 1385
rect 5018 1329 5037 1385
rect 5037 1329 5074 1385
rect 5099 1329 5155 1385
rect 5180 1329 5236 1385
rect 5261 1329 5273 1385
rect 5273 1329 5317 1385
rect 5363 1329 5419 1385
rect 5444 1329 5500 1385
rect 5525 1329 5561 1385
rect 5561 1329 5581 1385
rect 5606 1329 5662 1385
rect 5687 1329 5743 1385
rect 5768 1329 5797 1385
rect 5797 1329 5824 1385
rect 5849 1329 5905 1385
rect 5951 1329 5981 1385
rect 5981 1329 6007 1385
rect 6032 1329 6033 1385
rect 6033 1329 6088 1385
rect 6113 1329 6169 1385
rect 6194 1329 6217 1385
rect 6217 1329 6250 1385
rect 6275 1329 6331 1385
rect 6356 1329 6412 1385
rect 6437 1329 6453 1385
rect 6453 1329 6493 1385
rect 6517 1329 6573 1385
rect 6598 1329 6654 1385
rect 6679 1329 6689 1385
rect 6689 1329 6735 1385
rect 6760 1329 6816 1385
rect 6841 1329 6897 1385
rect 6922 1329 6925 1385
rect 6925 1329 6977 1385
rect 6977 1329 6978 1385
rect 7003 1329 7059 1385
rect 7090 1329 7146 1385
rect 7171 1329 7213 1385
rect 7213 1329 7227 1385
rect 7252 1329 7308 1385
rect 7333 1329 7389 1385
rect 7414 1329 7449 1385
rect 7449 1329 7470 1385
rect 7495 1329 7551 1385
rect 7576 1329 7632 1385
rect 7656 1329 7685 1385
rect 7685 1329 7712 1385
rect 7737 1329 7793 1385
rect 7818 1329 7869 1385
rect 7869 1329 7874 1385
rect 7899 1329 7921 1385
rect 7921 1329 7955 1385
rect 7980 1329 8036 1385
rect 8061 1329 8105 1385
rect 8105 1329 8117 1385
rect 8142 1329 8157 1385
rect 8157 1329 8198 1385
rect 8222 1329 8278 1385
rect 8303 1329 8341 1385
rect 8341 1329 8359 1385
rect 8384 1329 8393 1385
rect 8393 1329 8440 1385
rect 8465 1329 8521 1385
rect 8546 1329 8577 1385
rect 8577 1329 8602 1385
rect 8627 1329 8629 1385
rect 8629 1329 8683 1385
rect 8708 1329 8764 1385
rect 8788 1329 8813 1385
rect 8813 1329 8844 1385
rect 8869 1329 8925 1385
rect 8950 1329 9006 1385
rect 9031 1329 9049 1385
rect 9049 1329 9087 1385
rect 9112 1329 9168 1385
rect 9193 1329 9249 1385
rect 9274 1329 9285 1385
rect 9285 1329 9330 1385
rect 9357 1329 9413 1385
rect 9438 1329 9494 1385
rect 9519 1329 9521 1385
rect 9521 1329 9573 1385
rect 9573 1329 9575 1385
rect 9600 1329 9656 1385
rect 9681 1329 9737 1385
rect 9762 1329 9809 1385
rect 9809 1329 9818 1385
rect 9843 1329 9899 1385
rect 9923 1329 9979 1385
rect 10004 1329 10045 1385
rect 10045 1329 10060 1385
rect 10085 1329 10141 1385
rect 10166 1329 10222 1385
rect 10247 1329 10281 1385
rect 10281 1329 10303 1385
rect 10328 1329 10384 1385
rect 10409 1329 10465 1385
rect 10489 1329 10517 1385
rect 10517 1329 10545 1385
rect 10570 1329 10626 1385
rect 10651 1329 10701 1385
rect 10701 1329 10707 1385
rect 10732 1329 10753 1385
rect 10753 1329 10788 1385
rect 10813 1329 10869 1385
rect 10894 1329 10950 1385
rect 10975 1329 11031 1385
rect 11055 1329 11111 1385
rect 11136 1329 11192 1385
rect 11217 1329 11273 1385
rect 11298 1329 11354 1385
rect 11379 1329 11435 1385
rect 11460 1329 11516 1385
rect 11541 1329 11597 1385
rect 4915 610 4917 1170
rect 4917 610 4969 1170
rect 4969 610 4971 1170
rect 5151 610 5153 1170
rect 5153 610 5205 1170
rect 5205 610 5207 1170
rect 5387 610 5389 1170
rect 5389 610 5441 1170
rect 5441 610 5443 1170
rect 5623 610 5625 1170
rect 5625 610 5677 1170
rect 5677 610 5679 1170
rect 5859 610 5861 1170
rect 5861 610 5913 1170
rect 5913 610 5915 1170
rect 6095 610 6097 1170
rect 6097 610 6149 1170
rect 6149 610 6151 1170
rect 6331 610 6333 1170
rect 6333 610 6385 1170
rect 6385 610 6387 1170
rect 6567 610 6569 1170
rect 6569 610 6621 1170
rect 6621 610 6623 1170
rect 6803 610 6805 1170
rect 6805 610 6857 1170
rect 6857 610 6859 1170
rect 7039 610 7041 1170
rect 7041 610 7093 1170
rect 7093 610 7095 1170
rect 7275 610 7277 1170
rect 7277 610 7329 1170
rect 7329 610 7331 1170
rect 7511 610 7513 1170
rect 7513 610 7565 1170
rect 7565 610 7567 1170
rect 7747 610 7749 1170
rect 7749 610 7801 1170
rect 7801 610 7803 1170
rect 7983 610 7985 1170
rect 7985 610 8037 1170
rect 8037 610 8039 1170
rect 8219 610 8221 1170
rect 8221 610 8273 1170
rect 8273 610 8275 1170
rect 8455 610 8457 1170
rect 8457 610 8509 1170
rect 8509 610 8511 1170
rect 8691 610 8693 1170
rect 8693 610 8745 1170
rect 8745 610 8747 1170
rect 8927 610 8929 1170
rect 8929 610 8981 1170
rect 8981 610 8983 1170
rect 9163 610 9165 1170
rect 9165 610 9217 1170
rect 9217 610 9219 1170
rect 9399 610 9401 1170
rect 9401 610 9453 1170
rect 9453 610 9455 1170
rect 9635 610 9637 1170
rect 9637 610 9689 1170
rect 9689 610 9691 1170
rect 9871 610 9873 1170
rect 9873 610 9925 1170
rect 9925 610 9927 1170
rect 10107 610 10109 1170
rect 10109 610 10161 1170
rect 10161 610 10163 1170
rect 10343 610 10345 1170
rect 10345 610 10397 1170
rect 10397 610 10399 1170
rect 10579 610 10581 1170
rect 10581 610 10633 1170
rect 10633 610 10635 1170
rect 4915 -226 4917 334
rect 4917 -226 4969 334
rect 4969 -226 4971 334
rect 5151 -226 5153 334
rect 5153 -226 5205 334
rect 5205 -226 5207 334
rect 5387 -226 5389 334
rect 5389 -226 5441 334
rect 5441 -226 5443 334
rect 5623 -226 5625 334
rect 5625 -226 5677 334
rect 5677 -226 5679 334
rect 5859 -226 5861 334
rect 5861 -226 5913 334
rect 5913 -226 5915 334
rect 6095 -226 6097 334
rect 6097 -226 6149 334
rect 6149 -226 6151 334
rect 6331 -226 6333 334
rect 6333 -226 6385 334
rect 6385 -226 6387 334
rect 6567 -226 6569 334
rect 6569 -226 6621 334
rect 6621 -226 6623 334
rect 6803 -226 6805 334
rect 6805 -226 6857 334
rect 6857 -226 6859 334
rect 7039 -226 7041 334
rect 7041 -226 7093 334
rect 7093 -226 7095 334
rect 7275 -226 7277 334
rect 7277 -226 7329 334
rect 7329 -226 7331 334
rect 7511 -226 7513 334
rect 7513 -226 7565 334
rect 7565 -226 7567 334
rect 7747 -226 7749 334
rect 7749 -226 7801 334
rect 7801 -226 7803 334
rect 7983 -226 7985 334
rect 7985 -226 8037 334
rect 8037 -226 8039 334
rect 8219 -226 8221 334
rect 8221 -226 8273 334
rect 8273 -226 8275 334
rect 8455 -226 8457 334
rect 8457 -226 8509 334
rect 8509 -226 8511 334
rect 8691 -226 8693 334
rect 8693 -226 8745 334
rect 8745 -226 8747 334
rect 8927 -226 8929 334
rect 8929 -226 8981 334
rect 8981 -226 8983 334
rect 9163 -226 9165 334
rect 9165 -226 9217 334
rect 9217 -226 9219 334
rect 9399 -226 9401 334
rect 9401 -226 9453 334
rect 9453 -226 9455 334
rect 9635 -226 9637 334
rect 9637 -226 9689 334
rect 9689 -226 9691 334
rect 9871 -226 9873 334
rect 9873 -226 9925 334
rect 9925 -226 9927 334
rect 10107 -226 10109 334
rect 10109 -226 10161 334
rect 10161 -226 10163 334
rect 10343 -226 10345 334
rect 10345 -226 10397 334
rect 10397 -226 10399 334
rect 10579 -226 10581 334
rect 10581 -226 10633 334
rect 10633 -226 10635 334
rect 12607 1270 12609 1830
rect 12609 1270 12661 1830
rect 12661 1270 12663 1830
rect 12843 1270 12845 1830
rect 12845 1270 12897 1830
rect 12897 1270 12899 1830
rect 13079 1270 13081 1830
rect 13081 1270 13133 1830
rect 13133 1270 13135 1830
rect 13315 1270 13317 1830
rect 13317 1270 13369 1830
rect 13369 1270 13371 1830
rect 13551 1270 13553 1830
rect 13553 1270 13605 1830
rect 13605 1270 13607 1830
rect 13787 1270 13789 1830
rect 13789 1270 13841 1830
rect 13841 1270 13843 1830
rect 14023 1270 14025 1830
rect 14025 1270 14077 1830
rect 14077 1270 14079 1830
rect 14259 1270 14261 1830
rect 14261 1270 14313 1830
rect 14313 1270 14315 1830
rect 14495 1270 14497 1830
rect 14497 1270 14549 1830
rect 14549 1270 14551 1830
rect 14731 1270 14733 1830
rect 14733 1270 14785 1830
rect 14785 1270 14787 1830
rect 14967 1270 14969 1830
rect 14969 1270 15021 1830
rect 15021 1270 15023 1830
rect 15203 1270 15205 1830
rect 15205 1270 15257 1830
rect 15257 1270 15259 1830
rect 15439 1270 15441 1830
rect 15441 1270 15493 1830
rect 15493 1270 15495 1830
rect 16730 1270 16732 1830
rect 16732 1270 16784 1830
rect 16784 1270 16786 1830
rect 16966 1270 16968 1830
rect 16968 1270 17020 1830
rect 17020 1270 17022 1830
rect 17202 1270 17204 1830
rect 17204 1270 17256 1830
rect 17256 1270 17258 1830
rect 17438 1270 17440 1830
rect 17440 1270 17492 1830
rect 17492 1270 17494 1830
rect 17674 1270 17676 1830
rect 17676 1270 17728 1830
rect 17728 1270 17730 1830
rect 17910 1270 17912 1830
rect 17912 1270 17964 1830
rect 17964 1270 17966 1830
rect 18146 1270 18148 1830
rect 18148 1270 18200 1830
rect 18200 1270 18202 1830
rect 18382 1270 18384 1830
rect 18384 1270 18436 1830
rect 18436 1270 18438 1830
rect 18618 1270 18620 1830
rect 18620 1270 18672 1830
rect 18672 1270 18674 1830
rect 18854 1270 18856 1830
rect 18856 1270 18908 1830
rect 18908 1270 18910 1830
rect 19090 1270 19092 1830
rect 19092 1270 19144 1830
rect 19144 1270 19146 1830
rect 19326 1270 19328 1830
rect 19328 1270 19380 1830
rect 19380 1270 19382 1830
rect 19562 1270 19564 1830
rect 19564 1270 19616 1830
rect 19616 1270 19618 1830
rect 20853 1270 20855 1830
rect 20855 1270 20907 1830
rect 20907 1270 20909 1830
rect 21089 1270 21091 1830
rect 21091 1270 21143 1830
rect 21143 1270 21145 1830
rect 21325 1270 21327 1830
rect 21327 1270 21379 1830
rect 21379 1270 21381 1830
rect 21561 1270 21563 1830
rect 21563 1270 21615 1830
rect 21615 1270 21617 1830
rect 21797 1270 21799 1830
rect 21799 1270 21851 1830
rect 21851 1270 21853 1830
rect 22033 1270 22035 1830
rect 22035 1270 22087 1830
rect 22087 1270 22089 1830
rect 22269 1270 22271 1830
rect 22271 1270 22323 1830
rect 22323 1270 22325 1830
rect 22505 1270 22507 1830
rect 22507 1270 22559 1830
rect 22559 1270 22561 1830
rect 22741 1270 22743 1830
rect 22743 1270 22795 1830
rect 22795 1270 22797 1830
rect 22977 1270 22979 1830
rect 22979 1270 23031 1830
rect 23031 1270 23033 1830
rect 23213 1270 23215 1830
rect 23215 1270 23267 1830
rect 23267 1270 23269 1830
rect 23449 1270 23451 1830
rect 23451 1270 23503 1830
rect 23503 1270 23505 1830
rect 23685 1270 23687 1830
rect 23687 1270 23739 1830
rect 23739 1270 23741 1830
rect 4915 -1440 4917 -880
rect 4917 -1440 4969 -880
rect 4969 -1440 4971 -880
rect 5151 -1440 5153 -880
rect 5153 -1440 5205 -880
rect 5205 -1440 5207 -880
rect 5387 -1440 5389 -880
rect 5389 -1440 5441 -880
rect 5441 -1440 5443 -880
rect 5623 -1440 5625 -880
rect 5625 -1440 5677 -880
rect 5677 -1440 5679 -880
rect 5859 -1440 5861 -880
rect 5861 -1440 5913 -880
rect 5913 -1440 5915 -880
rect 6095 -1440 6097 -880
rect 6097 -1440 6149 -880
rect 6149 -1440 6151 -880
rect 6331 -1440 6333 -880
rect 6333 -1440 6385 -880
rect 6385 -1440 6387 -880
rect 6567 -1440 6569 -880
rect 6569 -1440 6621 -880
rect 6621 -1440 6623 -880
rect 6803 -1440 6805 -880
rect 6805 -1440 6857 -880
rect 6857 -1440 6859 -880
rect 7039 -1440 7041 -880
rect 7041 -1440 7093 -880
rect 7093 -1440 7095 -880
rect 7275 -1440 7277 -880
rect 7277 -1440 7329 -880
rect 7329 -1440 7331 -880
rect 7511 -1440 7513 -880
rect 7513 -1440 7565 -880
rect 7565 -1440 7567 -880
rect 7747 -1440 7749 -880
rect 7749 -1440 7801 -880
rect 7801 -1440 7803 -880
rect 7983 -1440 7985 -880
rect 7985 -1440 8037 -880
rect 8037 -1440 8039 -880
rect 8219 -1440 8221 -880
rect 8221 -1440 8273 -880
rect 8273 -1440 8275 -880
rect 8455 -1440 8457 -880
rect 8457 -1440 8509 -880
rect 8509 -1440 8511 -880
rect 8691 -1440 8693 -880
rect 8693 -1440 8745 -880
rect 8745 -1440 8747 -880
rect 8927 -1440 8929 -880
rect 8929 -1440 8981 -880
rect 8981 -1440 8983 -880
rect 9163 -1440 9165 -880
rect 9165 -1440 9217 -880
rect 9217 -1440 9219 -880
rect 9399 -1440 9401 -880
rect 9401 -1440 9453 -880
rect 9453 -1440 9455 -880
rect 9635 -1440 9637 -880
rect 9637 -1440 9689 -880
rect 9689 -1440 9691 -880
rect 9871 -1440 9873 -880
rect 9873 -1440 9925 -880
rect 9925 -1440 9927 -880
rect 10107 -1440 10109 -880
rect 10109 -1440 10161 -880
rect 10161 -1440 10163 -880
rect 10343 -1440 10345 -880
rect 10345 -1440 10397 -880
rect 10397 -1440 10399 -880
rect 10579 -1440 10581 -880
rect 10581 -1440 10633 -880
rect 10633 -1440 10635 -880
rect 4915 -2276 4917 -1716
rect 4917 -2276 4969 -1716
rect 4969 -2276 4971 -1716
rect 5151 -2276 5153 -1716
rect 5153 -2276 5205 -1716
rect 5205 -2276 5207 -1716
rect 5387 -2276 5389 -1716
rect 5389 -2276 5441 -1716
rect 5441 -2276 5443 -1716
rect 5623 -2276 5625 -1716
rect 5625 -2276 5677 -1716
rect 5677 -2276 5679 -1716
rect 5859 -2276 5861 -1716
rect 5861 -2276 5913 -1716
rect 5913 -2276 5915 -1716
rect 6095 -2276 6097 -1716
rect 6097 -2276 6149 -1716
rect 6149 -2276 6151 -1716
rect 6331 -2276 6333 -1716
rect 6333 -2276 6385 -1716
rect 6385 -2276 6387 -1716
rect 6567 -2276 6569 -1716
rect 6569 -2276 6621 -1716
rect 6621 -2276 6623 -1716
rect 6803 -2276 6805 -1716
rect 6805 -2276 6857 -1716
rect 6857 -2276 6859 -1716
rect 7039 -2276 7041 -1716
rect 7041 -2276 7093 -1716
rect 7093 -2276 7095 -1716
rect 7275 -2276 7277 -1716
rect 7277 -2276 7329 -1716
rect 7329 -2276 7331 -1716
rect 7511 -2276 7513 -1716
rect 7513 -2276 7565 -1716
rect 7565 -2276 7567 -1716
rect 7747 -2276 7749 -1716
rect 7749 -2276 7801 -1716
rect 7801 -2276 7803 -1716
rect 7983 -2276 7985 -1716
rect 7985 -2276 8037 -1716
rect 8037 -2276 8039 -1716
rect 8219 -2276 8221 -1716
rect 8221 -2276 8273 -1716
rect 8273 -2276 8275 -1716
rect 8455 -2276 8457 -1716
rect 8457 -2276 8509 -1716
rect 8509 -2276 8511 -1716
rect 8691 -2276 8693 -1716
rect 8693 -2276 8745 -1716
rect 8745 -2276 8747 -1716
rect 8927 -2276 8929 -1716
rect 8929 -2276 8981 -1716
rect 8981 -2276 8983 -1716
rect 9163 -2276 9165 -1716
rect 9165 -2276 9217 -1716
rect 9217 -2276 9219 -1716
rect 9399 -2276 9401 -1716
rect 9401 -2276 9453 -1716
rect 9453 -2276 9455 -1716
rect 9635 -2276 9637 -1716
rect 9637 -2276 9689 -1716
rect 9689 -2276 9691 -1716
rect 9871 -2276 9873 -1716
rect 9873 -2276 9925 -1716
rect 9925 -2276 9927 -1716
rect 10107 -2276 10109 -1716
rect 10109 -2276 10161 -1716
rect 10161 -2276 10163 -1716
rect 10343 -2276 10345 -1716
rect 10345 -2276 10397 -1716
rect 10397 -2276 10399 -1716
rect 10579 -2276 10581 -1716
rect 10581 -2276 10633 -1716
rect 10633 -2276 10635 -1716
rect 4919 -3490 4921 -2930
rect 4921 -3490 4973 -2930
rect 4973 -3490 4975 -2930
rect 5155 -3490 5157 -2930
rect 5157 -3490 5209 -2930
rect 5209 -3490 5211 -2930
rect 5391 -3490 5393 -2930
rect 5393 -3490 5445 -2930
rect 5445 -3490 5447 -2930
rect 5627 -3490 5629 -2930
rect 5629 -3490 5681 -2930
rect 5681 -3490 5683 -2930
rect 5863 -3490 5865 -2930
rect 5865 -3490 5917 -2930
rect 5917 -3490 5919 -2930
rect 6099 -3490 6101 -2930
rect 6101 -3490 6153 -2930
rect 6153 -3490 6155 -2930
rect 6335 -3490 6337 -2930
rect 6337 -3490 6389 -2930
rect 6389 -3490 6391 -2930
rect 6571 -3490 6573 -2930
rect 6573 -3490 6625 -2930
rect 6625 -3490 6627 -2930
rect 6807 -3490 6809 -2930
rect 6809 -3490 6861 -2930
rect 6861 -3490 6863 -2930
rect 7043 -3490 7045 -2930
rect 7045 -3490 7097 -2930
rect 7097 -3490 7099 -2930
rect 7279 -3490 7281 -2930
rect 7281 -3490 7333 -2930
rect 7333 -3490 7335 -2930
rect 7515 -3490 7517 -2930
rect 7517 -3490 7569 -2930
rect 7569 -3490 7571 -2930
rect 7751 -3490 7753 -2930
rect 7753 -3490 7805 -2930
rect 7805 -3490 7807 -2930
rect 7987 -3490 7989 -2930
rect 7989 -3490 8041 -2930
rect 8041 -3490 8043 -2930
rect 8223 -3490 8225 -2930
rect 8225 -3490 8277 -2930
rect 8277 -3490 8279 -2930
rect 8459 -3490 8461 -2930
rect 8461 -3490 8513 -2930
rect 8513 -3490 8515 -2930
rect 8695 -3490 8697 -2930
rect 8697 -3490 8749 -2930
rect 8749 -3490 8751 -2930
rect 8931 -3490 8933 -2930
rect 8933 -3490 8985 -2930
rect 8985 -3490 8987 -2930
rect 9167 -3490 9169 -2930
rect 9169 -3490 9221 -2930
rect 9221 -3490 9223 -2930
rect 9403 -3490 9405 -2930
rect 9405 -3490 9457 -2930
rect 9457 -3490 9459 -2930
rect 9639 -3490 9641 -2930
rect 9641 -3490 9693 -2930
rect 9693 -3490 9695 -2930
rect 9875 -3490 9877 -2930
rect 9877 -3490 9929 -2930
rect 9929 -3490 9931 -2930
rect 10111 -3490 10113 -2930
rect 10113 -3490 10165 -2930
rect 10165 -3490 10167 -2930
rect 10347 -3490 10349 -2930
rect 10349 -3490 10401 -2930
rect 10401 -3490 10403 -2930
rect 10583 -3490 10585 -2930
rect 10585 -3490 10637 -2930
rect 10637 -3490 10639 -2930
rect 4919 -4326 4921 -3766
rect 4921 -4326 4973 -3766
rect 4973 -4326 4975 -3766
rect 5155 -4326 5157 -3766
rect 5157 -4326 5209 -3766
rect 5209 -4326 5211 -3766
rect 5391 -4326 5393 -3766
rect 5393 -4326 5445 -3766
rect 5445 -4326 5447 -3766
rect 5627 -4326 5629 -3766
rect 5629 -4326 5681 -3766
rect 5681 -4326 5683 -3766
rect 5863 -4326 5865 -3766
rect 5865 -4326 5917 -3766
rect 5917 -4326 5919 -3766
rect 6099 -4326 6101 -3766
rect 6101 -4326 6153 -3766
rect 6153 -4326 6155 -3766
rect 6335 -4326 6337 -3766
rect 6337 -4326 6389 -3766
rect 6389 -4326 6391 -3766
rect 6571 -4326 6573 -3766
rect 6573 -4326 6625 -3766
rect 6625 -4326 6627 -3766
rect 6807 -4326 6809 -3766
rect 6809 -4326 6861 -3766
rect 6861 -4326 6863 -3766
rect 7043 -4326 7045 -3766
rect 7045 -4326 7097 -3766
rect 7097 -4326 7099 -3766
rect 7279 -4326 7281 -3766
rect 7281 -4326 7333 -3766
rect 7333 -4326 7335 -3766
rect 7515 -4326 7517 -3766
rect 7517 -4326 7569 -3766
rect 7569 -4326 7571 -3766
rect 7751 -4326 7753 -3766
rect 7753 -4326 7805 -3766
rect 7805 -4326 7807 -3766
rect 7987 -4326 7989 -3766
rect 7989 -4326 8041 -3766
rect 8041 -4326 8043 -3766
rect 8223 -4326 8225 -3766
rect 8225 -4326 8277 -3766
rect 8277 -4326 8279 -3766
rect 8459 -4326 8461 -3766
rect 8461 -4326 8513 -3766
rect 8513 -4326 8515 -3766
rect 8695 -4326 8697 -3766
rect 8697 -4326 8749 -3766
rect 8749 -4326 8751 -3766
rect 8931 -4326 8933 -3766
rect 8933 -4326 8985 -3766
rect 8985 -4326 8987 -3766
rect 9167 -4326 9169 -3766
rect 9169 -4326 9221 -3766
rect 9221 -4326 9223 -3766
rect 9403 -4326 9405 -3766
rect 9405 -4326 9457 -3766
rect 9457 -4326 9459 -3766
rect 9639 -4326 9641 -3766
rect 9641 -4326 9693 -3766
rect 9693 -4326 9695 -3766
rect 9875 -4326 9877 -3766
rect 9877 -4326 9929 -3766
rect 9929 -4326 9931 -3766
rect 10111 -4326 10113 -3766
rect 10113 -4326 10165 -3766
rect 10165 -4326 10167 -3766
rect 10347 -4326 10349 -3766
rect 10349 -4326 10401 -3766
rect 10401 -4326 10403 -3766
rect 10583 -4326 10585 -3766
rect 10585 -4326 10637 -3766
rect 10637 -4326 10639 -3766
rect 4919 -5540 4921 -4980
rect 4921 -5540 4973 -4980
rect 4973 -5540 4975 -4980
rect 5155 -5540 5157 -4980
rect 5157 -5540 5209 -4980
rect 5209 -5540 5211 -4980
rect 5391 -5540 5393 -4980
rect 5393 -5540 5445 -4980
rect 5445 -5540 5447 -4980
rect 5627 -5540 5629 -4980
rect 5629 -5540 5681 -4980
rect 5681 -5540 5683 -4980
rect 5863 -5540 5865 -4980
rect 5865 -5540 5917 -4980
rect 5917 -5540 5919 -4980
rect 6099 -5540 6101 -4980
rect 6101 -5540 6153 -4980
rect 6153 -5540 6155 -4980
rect 6335 -5540 6337 -4980
rect 6337 -5540 6389 -4980
rect 6389 -5540 6391 -4980
rect 6571 -5540 6573 -4980
rect 6573 -5540 6625 -4980
rect 6625 -5540 6627 -4980
rect 6807 -5540 6809 -4980
rect 6809 -5540 6861 -4980
rect 6861 -5540 6863 -4980
rect 7043 -5540 7045 -4980
rect 7045 -5540 7097 -4980
rect 7097 -5540 7099 -4980
rect 7279 -5540 7281 -4980
rect 7281 -5540 7333 -4980
rect 7333 -5540 7335 -4980
rect 7515 -5540 7517 -4980
rect 7517 -5540 7569 -4980
rect 7569 -5540 7571 -4980
rect 7751 -5540 7753 -4980
rect 7753 -5540 7805 -4980
rect 7805 -5540 7807 -4980
rect 7987 -5540 7989 -4980
rect 7989 -5540 8041 -4980
rect 8041 -5540 8043 -4980
rect 8223 -5540 8225 -4980
rect 8225 -5540 8277 -4980
rect 8277 -5540 8279 -4980
rect 8459 -5540 8461 -4980
rect 8461 -5540 8513 -4980
rect 8513 -5540 8515 -4980
rect 8695 -5540 8697 -4980
rect 8697 -5540 8749 -4980
rect 8749 -5540 8751 -4980
rect 8931 -5540 8933 -4980
rect 8933 -5540 8985 -4980
rect 8985 -5540 8987 -4980
rect 9167 -5540 9169 -4980
rect 9169 -5540 9221 -4980
rect 9221 -5540 9223 -4980
rect 9403 -5540 9405 -4980
rect 9405 -5540 9457 -4980
rect 9457 -5540 9459 -4980
rect 9639 -5540 9641 -4980
rect 9641 -5540 9693 -4980
rect 9693 -5540 9695 -4980
rect 9875 -5540 9877 -4980
rect 9877 -5540 9929 -4980
rect 9929 -5540 9931 -4980
rect 10111 -5540 10113 -4980
rect 10113 -5540 10165 -4980
rect 10165 -5540 10167 -4980
rect 10347 -5540 10349 -4980
rect 10349 -5540 10401 -4980
rect 10401 -5540 10403 -4980
rect 10583 -5540 10585 -4980
rect 10585 -5540 10637 -4980
rect 10637 -5540 10639 -4980
rect 4919 -6376 4921 -5816
rect 4921 -6376 4973 -5816
rect 4973 -6376 4975 -5816
rect 5155 -6376 5157 -5816
rect 5157 -6376 5209 -5816
rect 5209 -6376 5211 -5816
rect 5391 -6376 5393 -5816
rect 5393 -6376 5445 -5816
rect 5445 -6376 5447 -5816
rect 5627 -6376 5629 -5816
rect 5629 -6376 5681 -5816
rect 5681 -6376 5683 -5816
rect 5863 -6376 5865 -5816
rect 5865 -6376 5917 -5816
rect 5917 -6376 5919 -5816
rect 6099 -6376 6101 -5816
rect 6101 -6376 6153 -5816
rect 6153 -6376 6155 -5816
rect 6335 -6376 6337 -5816
rect 6337 -6376 6389 -5816
rect 6389 -6376 6391 -5816
rect 6571 -6376 6573 -5816
rect 6573 -6376 6625 -5816
rect 6625 -6376 6627 -5816
rect 6807 -6376 6809 -5816
rect 6809 -6376 6861 -5816
rect 6861 -6376 6863 -5816
rect 7043 -6376 7045 -5816
rect 7045 -6376 7097 -5816
rect 7097 -6376 7099 -5816
rect 7279 -6376 7281 -5816
rect 7281 -6376 7333 -5816
rect 7333 -6376 7335 -5816
rect 7515 -6376 7517 -5816
rect 7517 -6376 7569 -5816
rect 7569 -6376 7571 -5816
rect 7751 -6376 7753 -5816
rect 7753 -6376 7805 -5816
rect 7805 -6376 7807 -5816
rect 7987 -6376 7989 -5816
rect 7989 -6376 8041 -5816
rect 8041 -6376 8043 -5816
rect 8223 -6376 8225 -5816
rect 8225 -6376 8277 -5816
rect 8277 -6376 8279 -5816
rect 8459 -6376 8461 -5816
rect 8461 -6376 8513 -5816
rect 8513 -6376 8515 -5816
rect 8695 -6376 8697 -5816
rect 8697 -6376 8749 -5816
rect 8749 -6376 8751 -5816
rect 8931 -6376 8933 -5816
rect 8933 -6376 8985 -5816
rect 8985 -6376 8987 -5816
rect 9167 -6376 9169 -5816
rect 9169 -6376 9221 -5816
rect 9221 -6376 9223 -5816
rect 9403 -6376 9405 -5816
rect 9405 -6376 9457 -5816
rect 9457 -6376 9459 -5816
rect 9639 -6376 9641 -5816
rect 9641 -6376 9693 -5816
rect 9693 -6376 9695 -5816
rect 9875 -6376 9877 -5816
rect 9877 -6376 9929 -5816
rect 9929 -6376 9931 -5816
rect 10111 -6376 10113 -5816
rect 10113 -6376 10165 -5816
rect 10165 -6376 10167 -5816
rect 10347 -6376 10349 -5816
rect 10349 -6376 10401 -5816
rect 10401 -6376 10403 -5816
rect 10583 -6376 10585 -5816
rect 10585 -6376 10637 -5816
rect 10637 -6376 10639 -5816
rect 11066 -6700 11122 -6698
rect 11066 -6752 11068 -6700
rect 11068 -6752 11120 -6700
rect 11120 -6752 11122 -6700
rect 11066 -6754 11122 -6752
rect 11147 -6700 11203 -6698
rect 11147 -6752 11149 -6700
rect 11149 -6752 11201 -6700
rect 11201 -6752 11203 -6700
rect 11147 -6754 11203 -6752
rect 11228 -6700 11284 -6698
rect 11228 -6752 11230 -6700
rect 11230 -6752 11282 -6700
rect 11282 -6752 11284 -6700
rect 11228 -6754 11284 -6752
rect 11309 -6700 11365 -6698
rect 11309 -6752 11311 -6700
rect 11311 -6752 11363 -6700
rect 11363 -6752 11365 -6700
rect 11309 -6754 11365 -6752
rect 11390 -6700 11446 -6698
rect 11390 -6752 11392 -6700
rect 11392 -6752 11444 -6700
rect 11444 -6752 11446 -6700
rect 11390 -6754 11446 -6752
rect 11471 -6700 11527 -6698
rect 11471 -6752 11473 -6700
rect 11473 -6752 11525 -6700
rect 11525 -6752 11527 -6700
rect 11471 -6754 11527 -6752
rect 11552 -6700 11608 -6698
rect 11552 -6752 11554 -6700
rect 11554 -6752 11606 -6700
rect 11606 -6752 11608 -6700
rect 11552 -6754 11608 -6752
rect 11066 -6804 11122 -6802
rect 11066 -6856 11068 -6804
rect 11068 -6856 11120 -6804
rect 11120 -6856 11122 -6804
rect 11066 -6858 11122 -6856
rect 11147 -6804 11203 -6802
rect 11147 -6856 11149 -6804
rect 11149 -6856 11201 -6804
rect 11201 -6856 11203 -6804
rect 11147 -6858 11203 -6856
rect 11228 -6804 11284 -6802
rect 11228 -6856 11230 -6804
rect 11230 -6856 11282 -6804
rect 11282 -6856 11284 -6804
rect 11228 -6858 11284 -6856
rect 11309 -6804 11365 -6802
rect 11309 -6856 11311 -6804
rect 11311 -6856 11363 -6804
rect 11363 -6856 11365 -6804
rect 11309 -6858 11365 -6856
rect 11390 -6804 11446 -6802
rect 11390 -6856 11392 -6804
rect 11392 -6856 11444 -6804
rect 11444 -6856 11446 -6804
rect 11390 -6858 11446 -6856
rect 11471 -6804 11527 -6802
rect 11471 -6856 11473 -6804
rect 11473 -6856 11525 -6804
rect 11525 -6856 11527 -6804
rect 11471 -6858 11527 -6856
rect 11552 -6804 11608 -6802
rect 11552 -6856 11554 -6804
rect 11554 -6856 11606 -6804
rect 11606 -6856 11608 -6804
rect 11552 -6858 11608 -6856
rect 11066 -6908 11122 -6906
rect 11066 -6960 11068 -6908
rect 11068 -6960 11120 -6908
rect 11120 -6960 11122 -6908
rect 11066 -6962 11122 -6960
rect 11147 -6908 11203 -6906
rect 11147 -6960 11149 -6908
rect 11149 -6960 11201 -6908
rect 11201 -6960 11203 -6908
rect 11147 -6962 11203 -6960
rect 11228 -6908 11284 -6906
rect 11228 -6960 11230 -6908
rect 11230 -6960 11282 -6908
rect 11282 -6960 11284 -6908
rect 11228 -6962 11284 -6960
rect 11309 -6908 11365 -6906
rect 11309 -6960 11311 -6908
rect 11311 -6960 11363 -6908
rect 11363 -6960 11365 -6908
rect 11309 -6962 11365 -6960
rect 11390 -6908 11446 -6906
rect 11390 -6960 11392 -6908
rect 11392 -6960 11444 -6908
rect 11444 -6960 11446 -6908
rect 11390 -6962 11446 -6960
rect 11471 -6908 11527 -6906
rect 11471 -6960 11473 -6908
rect 11473 -6960 11525 -6908
rect 11525 -6960 11527 -6908
rect 11471 -6962 11527 -6960
rect 11552 -6908 11608 -6906
rect 11552 -6960 11554 -6908
rect 11554 -6960 11606 -6908
rect 11606 -6960 11608 -6908
rect 11552 -6962 11608 -6960
rect 4092 -7063 4148 -7061
rect 4092 -7115 4094 -7063
rect 4094 -7115 4146 -7063
rect 4146 -7115 4148 -7063
rect 4092 -7117 4148 -7115
rect 4173 -7063 4229 -7061
rect 4173 -7115 4175 -7063
rect 4175 -7115 4227 -7063
rect 4227 -7115 4229 -7063
rect 4173 -7117 4229 -7115
rect 4254 -7063 4310 -7061
rect 4254 -7115 4256 -7063
rect 4256 -7115 4308 -7063
rect 4308 -7115 4310 -7063
rect 4254 -7117 4310 -7115
rect 4335 -7063 4391 -7061
rect 4335 -7115 4337 -7063
rect 4337 -7115 4389 -7063
rect 4389 -7115 4391 -7063
rect 4335 -7117 4391 -7115
rect 4416 -7063 4472 -7061
rect 4416 -7115 4418 -7063
rect 4418 -7115 4470 -7063
rect 4470 -7115 4472 -7063
rect 4416 -7117 4472 -7115
rect 4497 -7063 4553 -7061
rect 4497 -7115 4499 -7063
rect 4499 -7115 4551 -7063
rect 4551 -7115 4553 -7063
rect 4497 -7117 4553 -7115
rect 4578 -7063 4634 -7061
rect 4578 -7115 4580 -7063
rect 4580 -7115 4632 -7063
rect 4632 -7115 4634 -7063
rect 4578 -7117 4634 -7115
rect 4660 -7063 4716 -7061
rect 4660 -7115 4662 -7063
rect 4662 -7115 4714 -7063
rect 4714 -7115 4716 -7063
rect 4660 -7117 4716 -7115
rect 4741 -7063 4797 -7061
rect 4741 -7115 4743 -7063
rect 4743 -7115 4795 -7063
rect 4795 -7115 4797 -7063
rect 4741 -7117 4797 -7115
rect 4822 -7063 4878 -7061
rect 4822 -7115 4824 -7063
rect 4824 -7115 4876 -7063
rect 4876 -7115 4878 -7063
rect 4822 -7117 4878 -7115
rect 4903 -7063 4959 -7061
rect 4903 -7115 4905 -7063
rect 4905 -7115 4957 -7063
rect 4957 -7115 4959 -7063
rect 4903 -7117 4959 -7115
rect 4984 -7063 5040 -7061
rect 4984 -7115 4986 -7063
rect 4986 -7115 5038 -7063
rect 5038 -7115 5040 -7063
rect 4984 -7117 5040 -7115
rect 5065 -7063 5121 -7061
rect 5065 -7115 5067 -7063
rect 5067 -7115 5119 -7063
rect 5119 -7115 5121 -7063
rect 5065 -7117 5121 -7115
rect 5146 -7063 5202 -7061
rect 5146 -7115 5148 -7063
rect 5148 -7115 5200 -7063
rect 5200 -7115 5202 -7063
rect 5146 -7117 5202 -7115
rect 5228 -7063 5284 -7061
rect 5228 -7115 5230 -7063
rect 5230 -7115 5282 -7063
rect 5282 -7115 5284 -7063
rect 5228 -7117 5284 -7115
rect 5309 -7063 5365 -7061
rect 5309 -7115 5311 -7063
rect 5311 -7115 5363 -7063
rect 5363 -7115 5365 -7063
rect 5309 -7117 5365 -7115
rect 5390 -7063 5446 -7061
rect 5390 -7115 5392 -7063
rect 5392 -7115 5444 -7063
rect 5444 -7115 5446 -7063
rect 5390 -7117 5446 -7115
rect 4092 -7167 4148 -7165
rect 4092 -7219 4094 -7167
rect 4094 -7219 4146 -7167
rect 4146 -7219 4148 -7167
rect 4092 -7221 4148 -7219
rect 4173 -7167 4229 -7165
rect 4173 -7219 4175 -7167
rect 4175 -7219 4227 -7167
rect 4227 -7219 4229 -7167
rect 4173 -7221 4229 -7219
rect 4254 -7167 4310 -7165
rect 4254 -7219 4256 -7167
rect 4256 -7219 4308 -7167
rect 4308 -7219 4310 -7167
rect 4254 -7221 4310 -7219
rect 4335 -7167 4391 -7165
rect 4335 -7219 4337 -7167
rect 4337 -7219 4389 -7167
rect 4389 -7219 4391 -7167
rect 4335 -7221 4391 -7219
rect 4416 -7167 4472 -7165
rect 4416 -7219 4418 -7167
rect 4418 -7219 4470 -7167
rect 4470 -7219 4472 -7167
rect 4416 -7221 4472 -7219
rect 4497 -7167 4553 -7165
rect 4497 -7219 4499 -7167
rect 4499 -7219 4551 -7167
rect 4551 -7219 4553 -7167
rect 4497 -7221 4553 -7219
rect 4578 -7167 4634 -7165
rect 4578 -7219 4580 -7167
rect 4580 -7219 4632 -7167
rect 4632 -7219 4634 -7167
rect 4578 -7221 4634 -7219
rect 4660 -7167 4716 -7165
rect 4660 -7219 4662 -7167
rect 4662 -7219 4714 -7167
rect 4714 -7219 4716 -7167
rect 4660 -7221 4716 -7219
rect 4741 -7167 4797 -7165
rect 4741 -7219 4743 -7167
rect 4743 -7219 4795 -7167
rect 4795 -7219 4797 -7167
rect 4741 -7221 4797 -7219
rect 4822 -7167 4878 -7165
rect 4822 -7219 4824 -7167
rect 4824 -7219 4876 -7167
rect 4876 -7219 4878 -7167
rect 4822 -7221 4878 -7219
rect 4903 -7167 4959 -7165
rect 4903 -7219 4905 -7167
rect 4905 -7219 4957 -7167
rect 4957 -7219 4959 -7167
rect 4903 -7221 4959 -7219
rect 4984 -7167 5040 -7165
rect 4984 -7219 4986 -7167
rect 4986 -7219 5038 -7167
rect 5038 -7219 5040 -7167
rect 4984 -7221 5040 -7219
rect 5065 -7167 5121 -7165
rect 5065 -7219 5067 -7167
rect 5067 -7219 5119 -7167
rect 5119 -7219 5121 -7167
rect 5065 -7221 5121 -7219
rect 5146 -7167 5202 -7165
rect 5146 -7219 5148 -7167
rect 5148 -7219 5200 -7167
rect 5200 -7219 5202 -7167
rect 5146 -7221 5202 -7219
rect 5228 -7167 5284 -7165
rect 5228 -7219 5230 -7167
rect 5230 -7219 5282 -7167
rect 5282 -7219 5284 -7167
rect 5228 -7221 5284 -7219
rect 5309 -7167 5365 -7165
rect 5309 -7219 5311 -7167
rect 5311 -7219 5363 -7167
rect 5363 -7219 5365 -7167
rect 5309 -7221 5365 -7219
rect 5390 -7167 5446 -7165
rect 5390 -7219 5392 -7167
rect 5392 -7219 5444 -7167
rect 5444 -7219 5446 -7167
rect 5390 -7221 5446 -7219
rect 4092 -7271 4148 -7269
rect 4092 -7323 4094 -7271
rect 4094 -7323 4146 -7271
rect 4146 -7323 4148 -7271
rect 4092 -7325 4148 -7323
rect 4173 -7271 4229 -7269
rect 4173 -7323 4175 -7271
rect 4175 -7323 4227 -7271
rect 4227 -7323 4229 -7271
rect 4173 -7325 4229 -7323
rect 4254 -7271 4310 -7269
rect 4254 -7323 4256 -7271
rect 4256 -7323 4308 -7271
rect 4308 -7323 4310 -7271
rect 4254 -7325 4310 -7323
rect 4335 -7271 4391 -7269
rect 4335 -7323 4337 -7271
rect 4337 -7323 4389 -7271
rect 4389 -7323 4391 -7271
rect 4335 -7325 4391 -7323
rect 4416 -7271 4472 -7269
rect 4416 -7323 4418 -7271
rect 4418 -7323 4470 -7271
rect 4470 -7323 4472 -7271
rect 4416 -7325 4472 -7323
rect 4497 -7271 4553 -7269
rect 4497 -7323 4499 -7271
rect 4499 -7323 4551 -7271
rect 4551 -7323 4553 -7271
rect 4497 -7325 4553 -7323
rect 4578 -7271 4634 -7269
rect 4578 -7323 4580 -7271
rect 4580 -7323 4632 -7271
rect 4632 -7323 4634 -7271
rect 4578 -7325 4634 -7323
rect 4660 -7271 4716 -7269
rect 4660 -7323 4662 -7271
rect 4662 -7323 4714 -7271
rect 4714 -7323 4716 -7271
rect 4660 -7325 4716 -7323
rect 4741 -7271 4797 -7269
rect 4741 -7323 4743 -7271
rect 4743 -7323 4795 -7271
rect 4795 -7323 4797 -7271
rect 4741 -7325 4797 -7323
rect 4822 -7271 4878 -7269
rect 4822 -7323 4824 -7271
rect 4824 -7323 4876 -7271
rect 4876 -7323 4878 -7271
rect 4822 -7325 4878 -7323
rect 4903 -7271 4959 -7269
rect 4903 -7323 4905 -7271
rect 4905 -7323 4957 -7271
rect 4957 -7323 4959 -7271
rect 4903 -7325 4959 -7323
rect 4984 -7271 5040 -7269
rect 4984 -7323 4986 -7271
rect 4986 -7323 5038 -7271
rect 5038 -7323 5040 -7271
rect 4984 -7325 5040 -7323
rect 5065 -7271 5121 -7269
rect 5065 -7323 5067 -7271
rect 5067 -7323 5119 -7271
rect 5119 -7323 5121 -7271
rect 5065 -7325 5121 -7323
rect 5146 -7271 5202 -7269
rect 5146 -7323 5148 -7271
rect 5148 -7323 5200 -7271
rect 5200 -7323 5202 -7271
rect 5146 -7325 5202 -7323
rect 5228 -7271 5284 -7269
rect 5228 -7323 5230 -7271
rect 5230 -7323 5282 -7271
rect 5282 -7323 5284 -7271
rect 5228 -7325 5284 -7323
rect 5309 -7271 5365 -7269
rect 5309 -7323 5311 -7271
rect 5311 -7323 5363 -7271
rect 5363 -7323 5365 -7271
rect 5309 -7325 5365 -7323
rect 5390 -7271 5446 -7269
rect 5390 -7323 5392 -7271
rect 5392 -7323 5444 -7271
rect 5444 -7323 5446 -7271
rect 5390 -7325 5446 -7323
rect 4092 -7375 4148 -7373
rect 4092 -7427 4094 -7375
rect 4094 -7427 4146 -7375
rect 4146 -7427 4148 -7375
rect 4092 -7429 4148 -7427
rect 4173 -7375 4229 -7373
rect 4173 -7427 4175 -7375
rect 4175 -7427 4227 -7375
rect 4227 -7427 4229 -7375
rect 4173 -7429 4229 -7427
rect 4254 -7375 4310 -7373
rect 4254 -7427 4256 -7375
rect 4256 -7427 4308 -7375
rect 4308 -7427 4310 -7375
rect 4254 -7429 4310 -7427
rect 4335 -7375 4391 -7373
rect 4335 -7427 4337 -7375
rect 4337 -7427 4389 -7375
rect 4389 -7427 4391 -7375
rect 4335 -7429 4391 -7427
rect 4416 -7375 4472 -7373
rect 4416 -7427 4418 -7375
rect 4418 -7427 4470 -7375
rect 4470 -7427 4472 -7375
rect 4416 -7429 4472 -7427
rect 4497 -7375 4553 -7373
rect 4497 -7427 4499 -7375
rect 4499 -7427 4551 -7375
rect 4551 -7427 4553 -7375
rect 4497 -7429 4553 -7427
rect 4578 -7375 4634 -7373
rect 4578 -7427 4580 -7375
rect 4580 -7427 4632 -7375
rect 4632 -7427 4634 -7375
rect 4578 -7429 4634 -7427
rect 4660 -7375 4716 -7373
rect 4660 -7427 4662 -7375
rect 4662 -7427 4714 -7375
rect 4714 -7427 4716 -7375
rect 4660 -7429 4716 -7427
rect 4741 -7375 4797 -7373
rect 4741 -7427 4743 -7375
rect 4743 -7427 4795 -7375
rect 4795 -7427 4797 -7375
rect 4741 -7429 4797 -7427
rect 4822 -7375 4878 -7373
rect 4822 -7427 4824 -7375
rect 4824 -7427 4876 -7375
rect 4876 -7427 4878 -7375
rect 4822 -7429 4878 -7427
rect 4903 -7375 4959 -7373
rect 4903 -7427 4905 -7375
rect 4905 -7427 4957 -7375
rect 4957 -7427 4959 -7375
rect 4903 -7429 4959 -7427
rect 4984 -7375 5040 -7373
rect 4984 -7427 4986 -7375
rect 4986 -7427 5038 -7375
rect 5038 -7427 5040 -7375
rect 4984 -7429 5040 -7427
rect 5065 -7375 5121 -7373
rect 5065 -7427 5067 -7375
rect 5067 -7427 5119 -7375
rect 5119 -7427 5121 -7375
rect 5065 -7429 5121 -7427
rect 5146 -7375 5202 -7373
rect 5146 -7427 5148 -7375
rect 5148 -7427 5200 -7375
rect 5200 -7427 5202 -7375
rect 5146 -7429 5202 -7427
rect 5228 -7375 5284 -7373
rect 5228 -7427 5230 -7375
rect 5230 -7427 5282 -7375
rect 5282 -7427 5284 -7375
rect 5228 -7429 5284 -7427
rect 5309 -7375 5365 -7373
rect 5309 -7427 5311 -7375
rect 5311 -7427 5363 -7375
rect 5363 -7427 5365 -7375
rect 5309 -7429 5365 -7427
rect 5390 -7375 5446 -7373
rect 5390 -7427 5392 -7375
rect 5392 -7427 5444 -7375
rect 5444 -7427 5446 -7375
rect 5390 -7429 5446 -7427
rect 4092 -7479 4148 -7477
rect 4092 -7531 4094 -7479
rect 4094 -7531 4146 -7479
rect 4146 -7531 4148 -7479
rect 4092 -7533 4148 -7531
rect 4173 -7479 4229 -7477
rect 4173 -7531 4175 -7479
rect 4175 -7531 4227 -7479
rect 4227 -7531 4229 -7479
rect 4173 -7533 4229 -7531
rect 4254 -7479 4310 -7477
rect 4254 -7531 4256 -7479
rect 4256 -7531 4308 -7479
rect 4308 -7531 4310 -7479
rect 4254 -7533 4310 -7531
rect 4335 -7479 4391 -7477
rect 4335 -7531 4337 -7479
rect 4337 -7531 4389 -7479
rect 4389 -7531 4391 -7479
rect 4335 -7533 4391 -7531
rect 4416 -7479 4472 -7477
rect 4416 -7531 4418 -7479
rect 4418 -7531 4470 -7479
rect 4470 -7531 4472 -7479
rect 4416 -7533 4472 -7531
rect 4497 -7479 4553 -7477
rect 4497 -7531 4499 -7479
rect 4499 -7531 4551 -7479
rect 4551 -7531 4553 -7479
rect 4497 -7533 4553 -7531
rect 4578 -7479 4634 -7477
rect 4578 -7531 4580 -7479
rect 4580 -7531 4632 -7479
rect 4632 -7531 4634 -7479
rect 4578 -7533 4634 -7531
rect 4660 -7479 4716 -7477
rect 4660 -7531 4662 -7479
rect 4662 -7531 4714 -7479
rect 4714 -7531 4716 -7479
rect 4660 -7533 4716 -7531
rect 4741 -7479 4797 -7477
rect 4741 -7531 4743 -7479
rect 4743 -7531 4795 -7479
rect 4795 -7531 4797 -7479
rect 4741 -7533 4797 -7531
rect 4822 -7479 4878 -7477
rect 4822 -7531 4824 -7479
rect 4824 -7531 4876 -7479
rect 4876 -7531 4878 -7479
rect 4822 -7533 4878 -7531
rect 4903 -7479 4959 -7477
rect 4903 -7531 4905 -7479
rect 4905 -7531 4957 -7479
rect 4957 -7531 4959 -7479
rect 4903 -7533 4959 -7531
rect 4984 -7479 5040 -7477
rect 4984 -7531 4986 -7479
rect 4986 -7531 5038 -7479
rect 5038 -7531 5040 -7479
rect 4984 -7533 5040 -7531
rect 5065 -7479 5121 -7477
rect 5065 -7531 5067 -7479
rect 5067 -7531 5119 -7479
rect 5119 -7531 5121 -7479
rect 5065 -7533 5121 -7531
rect 5146 -7479 5202 -7477
rect 5146 -7531 5148 -7479
rect 5148 -7531 5200 -7479
rect 5200 -7531 5202 -7479
rect 5146 -7533 5202 -7531
rect 5228 -7479 5284 -7477
rect 5228 -7531 5230 -7479
rect 5230 -7531 5282 -7479
rect 5282 -7531 5284 -7479
rect 5228 -7533 5284 -7531
rect 5309 -7479 5365 -7477
rect 5309 -7531 5311 -7479
rect 5311 -7531 5363 -7479
rect 5363 -7531 5365 -7479
rect 5309 -7533 5365 -7531
rect 5390 -7479 5446 -7477
rect 5390 -7531 5392 -7479
rect 5392 -7531 5444 -7479
rect 5444 -7531 5446 -7479
rect 5390 -7533 5446 -7531
rect 4092 -7583 4148 -7581
rect 4092 -7635 4094 -7583
rect 4094 -7635 4146 -7583
rect 4146 -7635 4148 -7583
rect 4092 -7637 4148 -7635
rect 4173 -7583 4229 -7581
rect 4173 -7635 4175 -7583
rect 4175 -7635 4227 -7583
rect 4227 -7635 4229 -7583
rect 4173 -7637 4229 -7635
rect 4254 -7583 4310 -7581
rect 4254 -7635 4256 -7583
rect 4256 -7635 4308 -7583
rect 4308 -7635 4310 -7583
rect 4254 -7637 4310 -7635
rect 4335 -7583 4391 -7581
rect 4335 -7635 4337 -7583
rect 4337 -7635 4389 -7583
rect 4389 -7635 4391 -7583
rect 4335 -7637 4391 -7635
rect 4416 -7583 4472 -7581
rect 4416 -7635 4418 -7583
rect 4418 -7635 4470 -7583
rect 4470 -7635 4472 -7583
rect 4416 -7637 4472 -7635
rect 4497 -7583 4553 -7581
rect 4497 -7635 4499 -7583
rect 4499 -7635 4551 -7583
rect 4551 -7635 4553 -7583
rect 4497 -7637 4553 -7635
rect 4578 -7583 4634 -7581
rect 4578 -7635 4580 -7583
rect 4580 -7635 4632 -7583
rect 4632 -7635 4634 -7583
rect 4578 -7637 4634 -7635
rect 4660 -7583 4716 -7581
rect 4660 -7635 4662 -7583
rect 4662 -7635 4714 -7583
rect 4714 -7635 4716 -7583
rect 4660 -7637 4716 -7635
rect 4741 -7583 4797 -7581
rect 4741 -7635 4743 -7583
rect 4743 -7635 4795 -7583
rect 4795 -7635 4797 -7583
rect 4741 -7637 4797 -7635
rect 4822 -7583 4878 -7581
rect 4822 -7635 4824 -7583
rect 4824 -7635 4876 -7583
rect 4876 -7635 4878 -7583
rect 4822 -7637 4878 -7635
rect 4903 -7583 4959 -7581
rect 4903 -7635 4905 -7583
rect 4905 -7635 4957 -7583
rect 4957 -7635 4959 -7583
rect 4903 -7637 4959 -7635
rect 4984 -7583 5040 -7581
rect 4984 -7635 4986 -7583
rect 4986 -7635 5038 -7583
rect 5038 -7635 5040 -7583
rect 4984 -7637 5040 -7635
rect 5065 -7583 5121 -7581
rect 5065 -7635 5067 -7583
rect 5067 -7635 5119 -7583
rect 5119 -7635 5121 -7583
rect 5065 -7637 5121 -7635
rect 5146 -7583 5202 -7581
rect 5146 -7635 5148 -7583
rect 5148 -7635 5200 -7583
rect 5200 -7635 5202 -7583
rect 5146 -7637 5202 -7635
rect 5228 -7583 5284 -7581
rect 5228 -7635 5230 -7583
rect 5230 -7635 5282 -7583
rect 5282 -7635 5284 -7583
rect 5228 -7637 5284 -7635
rect 5309 -7583 5365 -7581
rect 5309 -7635 5311 -7583
rect 5311 -7635 5363 -7583
rect 5363 -7635 5365 -7583
rect 5309 -7637 5365 -7635
rect 5390 -7583 5446 -7581
rect 5390 -7635 5392 -7583
rect 5392 -7635 5444 -7583
rect 5444 -7635 5446 -7583
rect 5390 -7637 5446 -7635
rect 4092 -7687 4148 -7685
rect 4092 -7739 4094 -7687
rect 4094 -7739 4146 -7687
rect 4146 -7739 4148 -7687
rect 4092 -7741 4148 -7739
rect 4173 -7687 4229 -7685
rect 4173 -7739 4175 -7687
rect 4175 -7739 4227 -7687
rect 4227 -7739 4229 -7687
rect 4173 -7741 4229 -7739
rect 4254 -7687 4310 -7685
rect 4254 -7739 4256 -7687
rect 4256 -7739 4308 -7687
rect 4308 -7739 4310 -7687
rect 4254 -7741 4310 -7739
rect 4335 -7687 4391 -7685
rect 4335 -7739 4337 -7687
rect 4337 -7739 4389 -7687
rect 4389 -7739 4391 -7687
rect 4335 -7741 4391 -7739
rect 4416 -7687 4472 -7685
rect 4416 -7739 4418 -7687
rect 4418 -7739 4470 -7687
rect 4470 -7739 4472 -7687
rect 4416 -7741 4472 -7739
rect 4497 -7687 4553 -7685
rect 4497 -7739 4499 -7687
rect 4499 -7739 4551 -7687
rect 4551 -7739 4553 -7687
rect 4497 -7741 4553 -7739
rect 4578 -7687 4634 -7685
rect 4578 -7739 4580 -7687
rect 4580 -7739 4632 -7687
rect 4632 -7739 4634 -7687
rect 4578 -7741 4634 -7739
rect 4660 -7687 4716 -7685
rect 4660 -7739 4662 -7687
rect 4662 -7739 4714 -7687
rect 4714 -7739 4716 -7687
rect 4660 -7741 4716 -7739
rect 4741 -7687 4797 -7685
rect 4741 -7739 4743 -7687
rect 4743 -7739 4795 -7687
rect 4795 -7739 4797 -7687
rect 4741 -7741 4797 -7739
rect 4822 -7687 4878 -7685
rect 4822 -7739 4824 -7687
rect 4824 -7739 4876 -7687
rect 4876 -7739 4878 -7687
rect 4822 -7741 4878 -7739
rect 4903 -7687 4959 -7685
rect 4903 -7739 4905 -7687
rect 4905 -7739 4957 -7687
rect 4957 -7739 4959 -7687
rect 4903 -7741 4959 -7739
rect 4984 -7687 5040 -7685
rect 4984 -7739 4986 -7687
rect 4986 -7739 5038 -7687
rect 5038 -7739 5040 -7687
rect 4984 -7741 5040 -7739
rect 5065 -7687 5121 -7685
rect 5065 -7739 5067 -7687
rect 5067 -7739 5119 -7687
rect 5119 -7739 5121 -7687
rect 5065 -7741 5121 -7739
rect 5146 -7687 5202 -7685
rect 5146 -7739 5148 -7687
rect 5148 -7739 5200 -7687
rect 5200 -7739 5202 -7687
rect 5146 -7741 5202 -7739
rect 5228 -7687 5284 -7685
rect 5228 -7739 5230 -7687
rect 5230 -7739 5282 -7687
rect 5282 -7739 5284 -7687
rect 5228 -7741 5284 -7739
rect 5309 -7687 5365 -7685
rect 5309 -7739 5311 -7687
rect 5311 -7739 5363 -7687
rect 5363 -7739 5365 -7687
rect 5309 -7741 5365 -7739
rect 5390 -7687 5446 -7685
rect 5390 -7739 5392 -7687
rect 5392 -7739 5444 -7687
rect 5444 -7739 5446 -7687
rect 5390 -7741 5446 -7739
rect 4092 -7791 4148 -7789
rect 4092 -7843 4094 -7791
rect 4094 -7843 4146 -7791
rect 4146 -7843 4148 -7791
rect 4092 -7845 4148 -7843
rect 4173 -7791 4229 -7789
rect 4173 -7843 4175 -7791
rect 4175 -7843 4227 -7791
rect 4227 -7843 4229 -7791
rect 4173 -7845 4229 -7843
rect 4254 -7791 4310 -7789
rect 4254 -7843 4256 -7791
rect 4256 -7843 4308 -7791
rect 4308 -7843 4310 -7791
rect 4254 -7845 4310 -7843
rect 4335 -7791 4391 -7789
rect 4335 -7843 4337 -7791
rect 4337 -7843 4389 -7791
rect 4389 -7843 4391 -7791
rect 4335 -7845 4391 -7843
rect 4416 -7791 4472 -7789
rect 4416 -7843 4418 -7791
rect 4418 -7843 4470 -7791
rect 4470 -7843 4472 -7791
rect 4416 -7845 4472 -7843
rect 4497 -7791 4553 -7789
rect 4497 -7843 4499 -7791
rect 4499 -7843 4551 -7791
rect 4551 -7843 4553 -7791
rect 4497 -7845 4553 -7843
rect 4578 -7791 4634 -7789
rect 4578 -7843 4580 -7791
rect 4580 -7843 4632 -7791
rect 4632 -7843 4634 -7791
rect 4578 -7845 4634 -7843
rect 4660 -7791 4716 -7789
rect 4660 -7843 4662 -7791
rect 4662 -7843 4714 -7791
rect 4714 -7843 4716 -7791
rect 4660 -7845 4716 -7843
rect 4741 -7791 4797 -7789
rect 4741 -7843 4743 -7791
rect 4743 -7843 4795 -7791
rect 4795 -7843 4797 -7791
rect 4741 -7845 4797 -7843
rect 4822 -7791 4878 -7789
rect 4822 -7843 4824 -7791
rect 4824 -7843 4876 -7791
rect 4876 -7843 4878 -7791
rect 4822 -7845 4878 -7843
rect 4903 -7791 4959 -7789
rect 4903 -7843 4905 -7791
rect 4905 -7843 4957 -7791
rect 4957 -7843 4959 -7791
rect 4903 -7845 4959 -7843
rect 4984 -7791 5040 -7789
rect 4984 -7843 4986 -7791
rect 4986 -7843 5038 -7791
rect 5038 -7843 5040 -7791
rect 4984 -7845 5040 -7843
rect 5065 -7791 5121 -7789
rect 5065 -7843 5067 -7791
rect 5067 -7843 5119 -7791
rect 5119 -7843 5121 -7791
rect 5065 -7845 5121 -7843
rect 5146 -7791 5202 -7789
rect 5146 -7843 5148 -7791
rect 5148 -7843 5200 -7791
rect 5200 -7843 5202 -7791
rect 5146 -7845 5202 -7843
rect 5228 -7791 5284 -7789
rect 5228 -7843 5230 -7791
rect 5230 -7843 5282 -7791
rect 5282 -7843 5284 -7791
rect 5228 -7845 5284 -7843
rect 5309 -7791 5365 -7789
rect 5309 -7843 5311 -7791
rect 5311 -7843 5363 -7791
rect 5363 -7843 5365 -7791
rect 5309 -7845 5365 -7843
rect 5390 -7791 5446 -7789
rect 5390 -7843 5392 -7791
rect 5392 -7843 5444 -7791
rect 5444 -7843 5446 -7791
rect 5390 -7845 5446 -7843
rect 5983 -7783 5985 -7223
rect 5985 -7783 6037 -7223
rect 6037 -7783 6039 -7223
rect 6219 -7783 6221 -7223
rect 6221 -7783 6273 -7223
rect 6273 -7783 6275 -7223
rect 6455 -7783 6457 -7223
rect 6457 -7783 6509 -7223
rect 6509 -7783 6511 -7223
rect 6691 -7783 6693 -7223
rect 6693 -7783 6745 -7223
rect 6745 -7783 6747 -7223
rect 6927 -7783 6929 -7223
rect 6929 -7783 6981 -7223
rect 6981 -7783 6983 -7223
rect 7163 -7783 7165 -7223
rect 7165 -7783 7217 -7223
rect 7217 -7783 7219 -7223
rect 7399 -7783 7401 -7223
rect 7401 -7783 7453 -7223
rect 7453 -7783 7455 -7223
rect 7635 -7783 7637 -7223
rect 7637 -7783 7689 -7223
rect 7689 -7783 7691 -7223
rect 7981 -7783 7983 -7223
rect 7983 -7783 8035 -7223
rect 8035 -7783 8037 -7223
rect 8217 -7783 8219 -7223
rect 8219 -7783 8271 -7223
rect 8271 -7783 8273 -7223
rect 8453 -7783 8455 -7223
rect 8455 -7783 8507 -7223
rect 8507 -7783 8509 -7223
rect 8689 -7783 8691 -7223
rect 8691 -7783 8743 -7223
rect 8743 -7783 8745 -7223
rect 8925 -7783 8927 -7223
rect 8927 -7783 8979 -7223
rect 8979 -7783 8981 -7223
rect 9161 -7783 9163 -7223
rect 9163 -7783 9215 -7223
rect 9215 -7783 9217 -7223
rect 9397 -7783 9399 -7223
rect 9399 -7783 9451 -7223
rect 9451 -7783 9453 -7223
rect 9633 -7783 9635 -7223
rect 9635 -7783 9687 -7223
rect 9687 -7783 9689 -7223
rect 4092 -7895 4148 -7893
rect 4092 -7947 4094 -7895
rect 4094 -7947 4146 -7895
rect 4146 -7947 4148 -7895
rect 4092 -7949 4148 -7947
rect 4173 -7895 4229 -7893
rect 4173 -7947 4175 -7895
rect 4175 -7947 4227 -7895
rect 4227 -7947 4229 -7895
rect 4173 -7949 4229 -7947
rect 4254 -7895 4310 -7893
rect 4254 -7947 4256 -7895
rect 4256 -7947 4308 -7895
rect 4308 -7947 4310 -7895
rect 4254 -7949 4310 -7947
rect 4335 -7895 4391 -7893
rect 4335 -7947 4337 -7895
rect 4337 -7947 4389 -7895
rect 4389 -7947 4391 -7895
rect 4335 -7949 4391 -7947
rect 4416 -7895 4472 -7893
rect 4416 -7947 4418 -7895
rect 4418 -7947 4470 -7895
rect 4470 -7947 4472 -7895
rect 4416 -7949 4472 -7947
rect 4497 -7895 4553 -7893
rect 4497 -7947 4499 -7895
rect 4499 -7947 4551 -7895
rect 4551 -7947 4553 -7895
rect 4497 -7949 4553 -7947
rect 4578 -7895 4634 -7893
rect 4578 -7947 4580 -7895
rect 4580 -7947 4632 -7895
rect 4632 -7947 4634 -7895
rect 4578 -7949 4634 -7947
rect 4660 -7895 4716 -7893
rect 4660 -7947 4662 -7895
rect 4662 -7947 4714 -7895
rect 4714 -7947 4716 -7895
rect 4660 -7949 4716 -7947
rect 4741 -7895 4797 -7893
rect 4741 -7947 4743 -7895
rect 4743 -7947 4795 -7895
rect 4795 -7947 4797 -7895
rect 4741 -7949 4797 -7947
rect 4822 -7895 4878 -7893
rect 4822 -7947 4824 -7895
rect 4824 -7947 4876 -7895
rect 4876 -7947 4878 -7895
rect 4822 -7949 4878 -7947
rect 4903 -7895 4959 -7893
rect 4903 -7947 4905 -7895
rect 4905 -7947 4957 -7895
rect 4957 -7947 4959 -7895
rect 4903 -7949 4959 -7947
rect 4984 -7895 5040 -7893
rect 4984 -7947 4986 -7895
rect 4986 -7947 5038 -7895
rect 5038 -7947 5040 -7895
rect 4984 -7949 5040 -7947
rect 5065 -7895 5121 -7893
rect 5065 -7947 5067 -7895
rect 5067 -7947 5119 -7895
rect 5119 -7947 5121 -7895
rect 5065 -7949 5121 -7947
rect 5146 -7895 5202 -7893
rect 5146 -7947 5148 -7895
rect 5148 -7947 5200 -7895
rect 5200 -7947 5202 -7895
rect 5146 -7949 5202 -7947
rect 5228 -7895 5284 -7893
rect 5228 -7947 5230 -7895
rect 5230 -7947 5282 -7895
rect 5282 -7947 5284 -7895
rect 5228 -7949 5284 -7947
rect 5309 -7895 5365 -7893
rect 5309 -7947 5311 -7895
rect 5311 -7947 5363 -7895
rect 5363 -7947 5365 -7895
rect 5309 -7949 5365 -7947
rect 5390 -7895 5446 -7893
rect 5390 -7947 5392 -7895
rect 5392 -7947 5444 -7895
rect 5444 -7947 5446 -7895
rect 5390 -7949 5446 -7947
rect 4092 -7999 4148 -7997
rect 4092 -8051 4094 -7999
rect 4094 -8051 4146 -7999
rect 4146 -8051 4148 -7999
rect 4092 -8053 4148 -8051
rect 4173 -7999 4229 -7997
rect 4173 -8051 4175 -7999
rect 4175 -8051 4227 -7999
rect 4227 -8051 4229 -7999
rect 4173 -8053 4229 -8051
rect 4254 -7999 4310 -7997
rect 4254 -8051 4256 -7999
rect 4256 -8051 4308 -7999
rect 4308 -8051 4310 -7999
rect 4254 -8053 4310 -8051
rect 4335 -7999 4391 -7997
rect 4335 -8051 4337 -7999
rect 4337 -8051 4389 -7999
rect 4389 -8051 4391 -7999
rect 4335 -8053 4391 -8051
rect 4416 -7999 4472 -7997
rect 4416 -8051 4418 -7999
rect 4418 -8051 4470 -7999
rect 4470 -8051 4472 -7999
rect 4416 -8053 4472 -8051
rect 4497 -7999 4553 -7997
rect 4497 -8051 4499 -7999
rect 4499 -8051 4551 -7999
rect 4551 -8051 4553 -7999
rect 4497 -8053 4553 -8051
rect 4578 -7999 4634 -7997
rect 4578 -8051 4580 -7999
rect 4580 -8051 4632 -7999
rect 4632 -8051 4634 -7999
rect 4578 -8053 4634 -8051
rect 4660 -7999 4716 -7997
rect 4660 -8051 4662 -7999
rect 4662 -8051 4714 -7999
rect 4714 -8051 4716 -7999
rect 4660 -8053 4716 -8051
rect 4741 -7999 4797 -7997
rect 4741 -8051 4743 -7999
rect 4743 -8051 4795 -7999
rect 4795 -8051 4797 -7999
rect 4741 -8053 4797 -8051
rect 4822 -7999 4878 -7997
rect 4822 -8051 4824 -7999
rect 4824 -8051 4876 -7999
rect 4876 -8051 4878 -7999
rect 4822 -8053 4878 -8051
rect 4903 -7999 4959 -7997
rect 4903 -8051 4905 -7999
rect 4905 -8051 4957 -7999
rect 4957 -8051 4959 -7999
rect 4903 -8053 4959 -8051
rect 4984 -7999 5040 -7997
rect 4984 -8051 4986 -7999
rect 4986 -8051 5038 -7999
rect 5038 -8051 5040 -7999
rect 4984 -8053 5040 -8051
rect 5065 -7999 5121 -7997
rect 5065 -8051 5067 -7999
rect 5067 -8051 5119 -7999
rect 5119 -8051 5121 -7999
rect 5065 -8053 5121 -8051
rect 5146 -7999 5202 -7997
rect 5146 -8051 5148 -7999
rect 5148 -8051 5200 -7999
rect 5200 -8051 5202 -7999
rect 5146 -8053 5202 -8051
rect 5228 -7999 5284 -7997
rect 5228 -8051 5230 -7999
rect 5230 -8051 5282 -7999
rect 5282 -8051 5284 -7999
rect 5228 -8053 5284 -8051
rect 5309 -7999 5365 -7997
rect 5309 -8051 5311 -7999
rect 5311 -8051 5363 -7999
rect 5363 -8051 5365 -7999
rect 5309 -8053 5365 -8051
rect 5390 -7999 5446 -7997
rect 5390 -8051 5392 -7999
rect 5392 -8051 5444 -7999
rect 5444 -8051 5446 -7999
rect 5390 -8053 5446 -8051
rect 4092 -8103 4148 -8101
rect 4092 -8155 4094 -8103
rect 4094 -8155 4146 -8103
rect 4146 -8155 4148 -8103
rect 4092 -8157 4148 -8155
rect 4173 -8103 4229 -8101
rect 4173 -8155 4175 -8103
rect 4175 -8155 4227 -8103
rect 4227 -8155 4229 -8103
rect 4173 -8157 4229 -8155
rect 4254 -8103 4310 -8101
rect 4254 -8155 4256 -8103
rect 4256 -8155 4308 -8103
rect 4308 -8155 4310 -8103
rect 4254 -8157 4310 -8155
rect 4335 -8103 4391 -8101
rect 4335 -8155 4337 -8103
rect 4337 -8155 4389 -8103
rect 4389 -8155 4391 -8103
rect 4335 -8157 4391 -8155
rect 4416 -8103 4472 -8101
rect 4416 -8155 4418 -8103
rect 4418 -8155 4470 -8103
rect 4470 -8155 4472 -8103
rect 4416 -8157 4472 -8155
rect 4497 -8103 4553 -8101
rect 4497 -8155 4499 -8103
rect 4499 -8155 4551 -8103
rect 4551 -8155 4553 -8103
rect 4497 -8157 4553 -8155
rect 4578 -8103 4634 -8101
rect 4578 -8155 4580 -8103
rect 4580 -8155 4632 -8103
rect 4632 -8155 4634 -8103
rect 4578 -8157 4634 -8155
rect 4660 -8103 4716 -8101
rect 4660 -8155 4662 -8103
rect 4662 -8155 4714 -8103
rect 4714 -8155 4716 -8103
rect 4660 -8157 4716 -8155
rect 4741 -8103 4797 -8101
rect 4741 -8155 4743 -8103
rect 4743 -8155 4795 -8103
rect 4795 -8155 4797 -8103
rect 4741 -8157 4797 -8155
rect 4822 -8103 4878 -8101
rect 4822 -8155 4824 -8103
rect 4824 -8155 4876 -8103
rect 4876 -8155 4878 -8103
rect 4822 -8157 4878 -8155
rect 4903 -8103 4959 -8101
rect 4903 -8155 4905 -8103
rect 4905 -8155 4957 -8103
rect 4957 -8155 4959 -8103
rect 4903 -8157 4959 -8155
rect 4984 -8103 5040 -8101
rect 4984 -8155 4986 -8103
rect 4986 -8155 5038 -8103
rect 5038 -8155 5040 -8103
rect 4984 -8157 5040 -8155
rect 5065 -8103 5121 -8101
rect 5065 -8155 5067 -8103
rect 5067 -8155 5119 -8103
rect 5119 -8155 5121 -8103
rect 5065 -8157 5121 -8155
rect 5146 -8103 5202 -8101
rect 5146 -8155 5148 -8103
rect 5148 -8155 5200 -8103
rect 5200 -8155 5202 -8103
rect 5146 -8157 5202 -8155
rect 5228 -8103 5284 -8101
rect 5228 -8155 5230 -8103
rect 5230 -8155 5282 -8103
rect 5282 -8155 5284 -8103
rect 5228 -8157 5284 -8155
rect 5309 -8103 5365 -8101
rect 5309 -8155 5311 -8103
rect 5311 -8155 5363 -8103
rect 5363 -8155 5365 -8103
rect 5309 -8157 5365 -8155
rect 5390 -8103 5446 -8101
rect 5390 -8155 5392 -8103
rect 5392 -8155 5444 -8103
rect 5444 -8155 5446 -8103
rect 5390 -8157 5446 -8155
rect 4092 -8207 4148 -8205
rect 4092 -8259 4094 -8207
rect 4094 -8259 4146 -8207
rect 4146 -8259 4148 -8207
rect 4092 -8261 4148 -8259
rect 4173 -8207 4229 -8205
rect 4173 -8259 4175 -8207
rect 4175 -8259 4227 -8207
rect 4227 -8259 4229 -8207
rect 4173 -8261 4229 -8259
rect 4254 -8207 4310 -8205
rect 4254 -8259 4256 -8207
rect 4256 -8259 4308 -8207
rect 4308 -8259 4310 -8207
rect 4254 -8261 4310 -8259
rect 4335 -8207 4391 -8205
rect 4335 -8259 4337 -8207
rect 4337 -8259 4389 -8207
rect 4389 -8259 4391 -8207
rect 4335 -8261 4391 -8259
rect 4416 -8207 4472 -8205
rect 4416 -8259 4418 -8207
rect 4418 -8259 4470 -8207
rect 4470 -8259 4472 -8207
rect 4416 -8261 4472 -8259
rect 4497 -8207 4553 -8205
rect 4497 -8259 4499 -8207
rect 4499 -8259 4551 -8207
rect 4551 -8259 4553 -8207
rect 4497 -8261 4553 -8259
rect 4578 -8207 4634 -8205
rect 4578 -8259 4580 -8207
rect 4580 -8259 4632 -8207
rect 4632 -8259 4634 -8207
rect 4578 -8261 4634 -8259
rect 4660 -8207 4716 -8205
rect 4660 -8259 4662 -8207
rect 4662 -8259 4714 -8207
rect 4714 -8259 4716 -8207
rect 4660 -8261 4716 -8259
rect 4741 -8207 4797 -8205
rect 4741 -8259 4743 -8207
rect 4743 -8259 4795 -8207
rect 4795 -8259 4797 -8207
rect 4741 -8261 4797 -8259
rect 4822 -8207 4878 -8205
rect 4822 -8259 4824 -8207
rect 4824 -8259 4876 -8207
rect 4876 -8259 4878 -8207
rect 4822 -8261 4878 -8259
rect 4903 -8207 4959 -8205
rect 4903 -8259 4905 -8207
rect 4905 -8259 4957 -8207
rect 4957 -8259 4959 -8207
rect 4903 -8261 4959 -8259
rect 4984 -8207 5040 -8205
rect 4984 -8259 4986 -8207
rect 4986 -8259 5038 -8207
rect 5038 -8259 5040 -8207
rect 4984 -8261 5040 -8259
rect 5065 -8207 5121 -8205
rect 5065 -8259 5067 -8207
rect 5067 -8259 5119 -8207
rect 5119 -8259 5121 -8207
rect 5065 -8261 5121 -8259
rect 5146 -8207 5202 -8205
rect 5146 -8259 5148 -8207
rect 5148 -8259 5200 -8207
rect 5200 -8259 5202 -8207
rect 5146 -8261 5202 -8259
rect 5228 -8207 5284 -8205
rect 5228 -8259 5230 -8207
rect 5230 -8259 5282 -8207
rect 5282 -8259 5284 -8207
rect 5228 -8261 5284 -8259
rect 5309 -8207 5365 -8205
rect 5309 -8259 5311 -8207
rect 5311 -8259 5363 -8207
rect 5363 -8259 5365 -8207
rect 5309 -8261 5365 -8259
rect 5390 -8207 5446 -8205
rect 5390 -8259 5392 -8207
rect 5392 -8259 5444 -8207
rect 5444 -8259 5446 -8207
rect 5390 -8261 5446 -8259
rect 4092 -8311 4148 -8309
rect 4092 -8363 4094 -8311
rect 4094 -8363 4146 -8311
rect 4146 -8363 4148 -8311
rect 4092 -8365 4148 -8363
rect 4173 -8311 4229 -8309
rect 4173 -8363 4175 -8311
rect 4175 -8363 4227 -8311
rect 4227 -8363 4229 -8311
rect 4173 -8365 4229 -8363
rect 4254 -8311 4310 -8309
rect 4254 -8363 4256 -8311
rect 4256 -8363 4308 -8311
rect 4308 -8363 4310 -8311
rect 4254 -8365 4310 -8363
rect 4335 -8311 4391 -8309
rect 4335 -8363 4337 -8311
rect 4337 -8363 4389 -8311
rect 4389 -8363 4391 -8311
rect 4335 -8365 4391 -8363
rect 4416 -8311 4472 -8309
rect 4416 -8363 4418 -8311
rect 4418 -8363 4470 -8311
rect 4470 -8363 4472 -8311
rect 4416 -8365 4472 -8363
rect 4497 -8311 4553 -8309
rect 4497 -8363 4499 -8311
rect 4499 -8363 4551 -8311
rect 4551 -8363 4553 -8311
rect 4497 -8365 4553 -8363
rect 4578 -8311 4634 -8309
rect 4578 -8363 4580 -8311
rect 4580 -8363 4632 -8311
rect 4632 -8363 4634 -8311
rect 4578 -8365 4634 -8363
rect 4660 -8311 4716 -8309
rect 4660 -8363 4662 -8311
rect 4662 -8363 4714 -8311
rect 4714 -8363 4716 -8311
rect 4660 -8365 4716 -8363
rect 4741 -8311 4797 -8309
rect 4741 -8363 4743 -8311
rect 4743 -8363 4795 -8311
rect 4795 -8363 4797 -8311
rect 4741 -8365 4797 -8363
rect 4822 -8311 4878 -8309
rect 4822 -8363 4824 -8311
rect 4824 -8363 4876 -8311
rect 4876 -8363 4878 -8311
rect 4822 -8365 4878 -8363
rect 4903 -8311 4959 -8309
rect 4903 -8363 4905 -8311
rect 4905 -8363 4957 -8311
rect 4957 -8363 4959 -8311
rect 4903 -8365 4959 -8363
rect 4984 -8311 5040 -8309
rect 4984 -8363 4986 -8311
rect 4986 -8363 5038 -8311
rect 5038 -8363 5040 -8311
rect 4984 -8365 5040 -8363
rect 5065 -8311 5121 -8309
rect 5065 -8363 5067 -8311
rect 5067 -8363 5119 -8311
rect 5119 -8363 5121 -8311
rect 5065 -8365 5121 -8363
rect 5146 -8311 5202 -8309
rect 5146 -8363 5148 -8311
rect 5148 -8363 5200 -8311
rect 5200 -8363 5202 -8311
rect 5146 -8365 5202 -8363
rect 5228 -8311 5284 -8309
rect 5228 -8363 5230 -8311
rect 5230 -8363 5282 -8311
rect 5282 -8363 5284 -8311
rect 5228 -8365 5284 -8363
rect 5309 -8311 5365 -8309
rect 5309 -8363 5311 -8311
rect 5311 -8363 5363 -8311
rect 5363 -8363 5365 -8311
rect 5309 -8365 5365 -8363
rect 5390 -8311 5446 -8309
rect 5390 -8363 5392 -8311
rect 5392 -8363 5444 -8311
rect 5444 -8363 5446 -8311
rect 5390 -8365 5446 -8363
rect 4092 -8415 4148 -8413
rect 4092 -8467 4094 -8415
rect 4094 -8467 4146 -8415
rect 4146 -8467 4148 -8415
rect 4092 -8469 4148 -8467
rect 4173 -8415 4229 -8413
rect 4173 -8467 4175 -8415
rect 4175 -8467 4227 -8415
rect 4227 -8467 4229 -8415
rect 4173 -8469 4229 -8467
rect 4254 -8415 4310 -8413
rect 4254 -8467 4256 -8415
rect 4256 -8467 4308 -8415
rect 4308 -8467 4310 -8415
rect 4254 -8469 4310 -8467
rect 4335 -8415 4391 -8413
rect 4335 -8467 4337 -8415
rect 4337 -8467 4389 -8415
rect 4389 -8467 4391 -8415
rect 4335 -8469 4391 -8467
rect 4416 -8415 4472 -8413
rect 4416 -8467 4418 -8415
rect 4418 -8467 4470 -8415
rect 4470 -8467 4472 -8415
rect 4416 -8469 4472 -8467
rect 4497 -8415 4553 -8413
rect 4497 -8467 4499 -8415
rect 4499 -8467 4551 -8415
rect 4551 -8467 4553 -8415
rect 4497 -8469 4553 -8467
rect 4578 -8415 4634 -8413
rect 4578 -8467 4580 -8415
rect 4580 -8467 4632 -8415
rect 4632 -8467 4634 -8415
rect 4578 -8469 4634 -8467
rect 4660 -8415 4716 -8413
rect 4660 -8467 4662 -8415
rect 4662 -8467 4714 -8415
rect 4714 -8467 4716 -8415
rect 4660 -8469 4716 -8467
rect 4741 -8415 4797 -8413
rect 4741 -8467 4743 -8415
rect 4743 -8467 4795 -8415
rect 4795 -8467 4797 -8415
rect 4741 -8469 4797 -8467
rect 4822 -8415 4878 -8413
rect 4822 -8467 4824 -8415
rect 4824 -8467 4876 -8415
rect 4876 -8467 4878 -8415
rect 4822 -8469 4878 -8467
rect 4903 -8415 4959 -8413
rect 4903 -8467 4905 -8415
rect 4905 -8467 4957 -8415
rect 4957 -8467 4959 -8415
rect 4903 -8469 4959 -8467
rect 4984 -8415 5040 -8413
rect 4984 -8467 4986 -8415
rect 4986 -8467 5038 -8415
rect 5038 -8467 5040 -8415
rect 4984 -8469 5040 -8467
rect 5065 -8415 5121 -8413
rect 5065 -8467 5067 -8415
rect 5067 -8467 5119 -8415
rect 5119 -8467 5121 -8415
rect 5065 -8469 5121 -8467
rect 5146 -8415 5202 -8413
rect 5146 -8467 5148 -8415
rect 5148 -8467 5200 -8415
rect 5200 -8467 5202 -8415
rect 5146 -8469 5202 -8467
rect 5228 -8415 5284 -8413
rect 5228 -8467 5230 -8415
rect 5230 -8467 5282 -8415
rect 5282 -8467 5284 -8415
rect 5228 -8469 5284 -8467
rect 5309 -8415 5365 -8413
rect 5309 -8467 5311 -8415
rect 5311 -8467 5363 -8415
rect 5363 -8467 5365 -8415
rect 5309 -8469 5365 -8467
rect 5390 -8415 5446 -8413
rect 5390 -8467 5392 -8415
rect 5392 -8467 5444 -8415
rect 5444 -8467 5446 -8415
rect 5390 -8469 5446 -8467
rect 4092 -8519 4148 -8517
rect 4092 -8571 4094 -8519
rect 4094 -8571 4146 -8519
rect 4146 -8571 4148 -8519
rect 4092 -8573 4148 -8571
rect 4173 -8519 4229 -8517
rect 4173 -8571 4175 -8519
rect 4175 -8571 4227 -8519
rect 4227 -8571 4229 -8519
rect 4173 -8573 4229 -8571
rect 4254 -8519 4310 -8517
rect 4254 -8571 4256 -8519
rect 4256 -8571 4308 -8519
rect 4308 -8571 4310 -8519
rect 4254 -8573 4310 -8571
rect 4335 -8519 4391 -8517
rect 4335 -8571 4337 -8519
rect 4337 -8571 4389 -8519
rect 4389 -8571 4391 -8519
rect 4335 -8573 4391 -8571
rect 4416 -8519 4472 -8517
rect 4416 -8571 4418 -8519
rect 4418 -8571 4470 -8519
rect 4470 -8571 4472 -8519
rect 4416 -8573 4472 -8571
rect 4497 -8519 4553 -8517
rect 4497 -8571 4499 -8519
rect 4499 -8571 4551 -8519
rect 4551 -8571 4553 -8519
rect 4497 -8573 4553 -8571
rect 4578 -8519 4634 -8517
rect 4578 -8571 4580 -8519
rect 4580 -8571 4632 -8519
rect 4632 -8571 4634 -8519
rect 4578 -8573 4634 -8571
rect 4660 -8519 4716 -8517
rect 4660 -8571 4662 -8519
rect 4662 -8571 4714 -8519
rect 4714 -8571 4716 -8519
rect 4660 -8573 4716 -8571
rect 4741 -8519 4797 -8517
rect 4741 -8571 4743 -8519
rect 4743 -8571 4795 -8519
rect 4795 -8571 4797 -8519
rect 4741 -8573 4797 -8571
rect 4822 -8519 4878 -8517
rect 4822 -8571 4824 -8519
rect 4824 -8571 4876 -8519
rect 4876 -8571 4878 -8519
rect 4822 -8573 4878 -8571
rect 4903 -8519 4959 -8517
rect 4903 -8571 4905 -8519
rect 4905 -8571 4957 -8519
rect 4957 -8571 4959 -8519
rect 4903 -8573 4959 -8571
rect 4984 -8519 5040 -8517
rect 4984 -8571 4986 -8519
rect 4986 -8571 5038 -8519
rect 5038 -8571 5040 -8519
rect 4984 -8573 5040 -8571
rect 5065 -8519 5121 -8517
rect 5065 -8571 5067 -8519
rect 5067 -8571 5119 -8519
rect 5119 -8571 5121 -8519
rect 5065 -8573 5121 -8571
rect 5146 -8519 5202 -8517
rect 5146 -8571 5148 -8519
rect 5148 -8571 5200 -8519
rect 5200 -8571 5202 -8519
rect 5146 -8573 5202 -8571
rect 5228 -8519 5284 -8517
rect 5228 -8571 5230 -8519
rect 5230 -8571 5282 -8519
rect 5282 -8571 5284 -8519
rect 5228 -8573 5284 -8571
rect 5309 -8519 5365 -8517
rect 5309 -8571 5311 -8519
rect 5311 -8571 5363 -8519
rect 5363 -8571 5365 -8519
rect 5309 -8573 5365 -8571
rect 5390 -8519 5446 -8517
rect 5390 -8571 5392 -8519
rect 5392 -8571 5444 -8519
rect 5444 -8571 5446 -8519
rect 5390 -8573 5446 -8571
rect 5983 -8601 5985 -8041
rect 5985 -8601 6037 -8041
rect 6037 -8601 6039 -8041
rect 6219 -8601 6221 -8041
rect 6221 -8601 6273 -8041
rect 6273 -8601 6275 -8041
rect 6455 -8601 6457 -8041
rect 6457 -8601 6509 -8041
rect 6509 -8601 6511 -8041
rect 6691 -8601 6693 -8041
rect 6693 -8601 6745 -8041
rect 6745 -8601 6747 -8041
rect 6927 -8601 6929 -8041
rect 6929 -8601 6981 -8041
rect 6981 -8601 6983 -8041
rect 7163 -8601 7165 -8041
rect 7165 -8601 7217 -8041
rect 7217 -8601 7219 -8041
rect 7399 -8601 7401 -8041
rect 7401 -8601 7453 -8041
rect 7453 -8601 7455 -8041
rect 10625 -7515 10627 -7395
rect 10627 -7515 10679 -7395
rect 10679 -7515 10681 -7395
rect 10941 -7515 10943 -7395
rect 10943 -7515 10995 -7395
rect 10995 -7515 10997 -7395
rect 11257 -7515 11259 -7395
rect 11259 -7515 11311 -7395
rect 11311 -7515 11313 -7395
rect 11573 -7515 11575 -7395
rect 11575 -7515 11627 -7395
rect 11627 -7515 11629 -7395
rect 11889 -7515 11891 -7395
rect 11891 -7515 11943 -7395
rect 11943 -7515 11945 -7395
rect 7635 -8601 7637 -8041
rect 7637 -8601 7689 -8041
rect 7689 -8601 7691 -8041
rect 7981 -8601 7983 -8041
rect 7983 -8601 8035 -8041
rect 8035 -8601 8037 -8041
rect 8217 -8601 8219 -8041
rect 8219 -8601 8271 -8041
rect 8271 -8601 8273 -8041
rect 8453 -8601 8455 -8041
rect 8455 -8601 8507 -8041
rect 8507 -8601 8509 -8041
rect 8689 -8601 8691 -8041
rect 8691 -8601 8743 -8041
rect 8743 -8601 8745 -8041
rect 8925 -8601 8927 -8041
rect 8927 -8601 8979 -8041
rect 8979 -8601 8981 -8041
rect 9161 -8601 9163 -8041
rect 9163 -8601 9215 -8041
rect 9215 -8601 9217 -8041
rect 9397 -8601 9399 -8041
rect 9399 -8601 9451 -8041
rect 9451 -8601 9453 -8041
rect 9633 -8601 9635 -8041
rect 9635 -8601 9687 -8041
rect 9687 -8601 9689 -8041
rect 10834 -8076 10890 -8020
rect 10915 -8076 10971 -8020
rect 10996 -8076 11052 -8020
rect 11077 -8076 11133 -8020
rect 11158 -8076 11214 -8020
rect 11239 -8076 11295 -8020
rect 11320 -8076 11376 -8020
rect 11401 -8076 11457 -8020
rect 11482 -8076 11538 -8020
rect 11563 -8076 11619 -8020
rect 11644 -8076 11700 -8020
rect 11725 -8076 11781 -8020
rect 11806 -8076 11862 -8020
rect 10834 -8180 10890 -8124
rect 10915 -8180 10971 -8124
rect 10996 -8180 11052 -8124
rect 11077 -8180 11133 -8124
rect 11158 -8180 11214 -8124
rect 11239 -8180 11295 -8124
rect 11320 -8180 11376 -8124
rect 11401 -8180 11457 -8124
rect 11482 -8180 11538 -8124
rect 11563 -8180 11619 -8124
rect 11644 -8180 11700 -8124
rect 11725 -8180 11781 -8124
rect 11806 -8180 11862 -8124
rect 12205 -7515 12207 -7395
rect 12207 -7515 12259 -7395
rect 12259 -7515 12261 -7395
rect 12523 -8059 12525 -7219
rect 12525 -8059 12577 -7219
rect 12577 -8059 12579 -7219
rect 12671 -8059 12673 -7219
rect 12673 -8059 12725 -7219
rect 12725 -8059 12727 -7219
rect 12819 -8059 12821 -7219
rect 12821 -8059 12873 -7219
rect 12873 -8059 12875 -7219
rect 12967 -8059 12969 -7219
rect 12969 -8059 13021 -7219
rect 13021 -8059 13023 -7219
rect 13115 -8059 13117 -7219
rect 13117 -8059 13169 -7219
rect 13169 -8059 13171 -7219
rect 13263 -8059 13265 -7219
rect 13265 -8059 13317 -7219
rect 13317 -8059 13319 -7219
rect 13411 -8059 13413 -7219
rect 13413 -8059 13465 -7219
rect 13465 -8059 13467 -7219
rect 13559 -8059 13561 -7219
rect 13561 -8059 13613 -7219
rect 13613 -8059 13615 -7219
rect 13707 -8059 13709 -7219
rect 13709 -8059 13761 -7219
rect 13761 -8059 13763 -7219
rect 13855 -8059 13857 -7219
rect 13857 -8059 13909 -7219
rect 13909 -8059 13911 -7219
rect 14003 -8059 14005 -7219
rect 14005 -8059 14057 -7219
rect 14057 -8059 14059 -7219
rect 14151 -8059 14153 -7219
rect 14153 -8059 14205 -7219
rect 14205 -8059 14207 -7219
rect 14299 -8059 14301 -7219
rect 14301 -8059 14353 -7219
rect 14353 -8059 14355 -7219
rect 14447 -8059 14449 -7219
rect 14449 -8059 14501 -7219
rect 14501 -8059 14503 -7219
rect 14595 -8059 14597 -7219
rect 14597 -8059 14649 -7219
rect 14649 -8059 14651 -7219
rect 14743 -8059 14745 -7219
rect 14745 -8059 14797 -7219
rect 14797 -8059 14799 -7219
rect 14891 -8059 14893 -7219
rect 14893 -8059 14945 -7219
rect 14945 -8059 14947 -7219
rect 15039 -8059 15041 -7219
rect 15041 -8059 15093 -7219
rect 15093 -8059 15095 -7219
rect 15187 -8059 15189 -7219
rect 15189 -8059 15241 -7219
rect 15241 -8059 15243 -7219
rect 15335 -8059 15337 -7219
rect 15337 -8059 15389 -7219
rect 15389 -8059 15391 -7219
rect 15483 -8059 15485 -7219
rect 15485 -8059 15537 -7219
rect 15537 -8059 15539 -7219
rect 15631 -8059 15633 -7219
rect 15633 -8059 15685 -7219
rect 15685 -8059 15687 -7219
rect 15779 -8059 15781 -7219
rect 15781 -8059 15833 -7219
rect 15833 -8059 15835 -7219
rect 15927 -8059 15929 -7219
rect 15929 -8059 15981 -7219
rect 15981 -8059 15983 -7219
rect 16075 -8059 16077 -7219
rect 16077 -8059 16129 -7219
rect 16129 -8059 16131 -7219
rect 16223 -8059 16225 -7219
rect 16225 -8059 16277 -7219
rect 16277 -8059 16279 -7219
rect 16371 -8059 16373 -7219
rect 16373 -8059 16425 -7219
rect 16425 -8059 16427 -7219
rect 16519 -8059 16521 -7219
rect 16521 -8059 16573 -7219
rect 16573 -8059 16575 -7219
rect 16667 -8059 16669 -7219
rect 16669 -8059 16721 -7219
rect 16721 -8059 16723 -7219
rect 16815 -8059 16817 -7219
rect 16817 -8059 16869 -7219
rect 16869 -8059 16871 -7219
rect 16963 -8059 16965 -7219
rect 16965 -8059 17017 -7219
rect 17017 -8059 17019 -7219
rect 17111 -8059 17113 -7219
rect 17113 -8059 17165 -7219
rect 17165 -8059 17167 -7219
rect 17259 -8059 17261 -7219
rect 17261 -8059 17313 -7219
rect 17313 -8059 17315 -7219
rect 17407 -8059 17409 -7219
rect 17409 -8059 17461 -7219
rect 17461 -8059 17463 -7219
rect 17555 -8059 17557 -7219
rect 17557 -8059 17609 -7219
rect 17609 -8059 17611 -7219
rect 17703 -8059 17705 -7219
rect 17705 -8059 17757 -7219
rect 17757 -8059 17759 -7219
rect 17851 -8059 17853 -7219
rect 17853 -8059 17905 -7219
rect 17905 -8059 17907 -7219
rect 17999 -8059 18001 -7219
rect 18001 -8059 18053 -7219
rect 18053 -8059 18055 -7219
rect 18147 -8059 18149 -7219
rect 18149 -8059 18201 -7219
rect 18201 -8059 18203 -7219
rect 18295 -8059 18297 -7219
rect 18297 -8059 18349 -7219
rect 18349 -8059 18351 -7219
rect 18443 -8059 18445 -7219
rect 18445 -8059 18497 -7219
rect 18497 -8059 18499 -7219
rect 18591 -8059 18593 -7219
rect 18593 -8059 18645 -7219
rect 18645 -8059 18647 -7219
rect 18739 -8059 18741 -7219
rect 18741 -8059 18793 -7219
rect 18793 -8059 18795 -7219
rect 18887 -8059 18889 -7219
rect 18889 -8059 18941 -7219
rect 18941 -8059 18943 -7219
rect 19035 -8059 19037 -7219
rect 19037 -8059 19089 -7219
rect 19089 -8059 19091 -7219
rect 19183 -8059 19185 -7219
rect 19185 -8059 19237 -7219
rect 19237 -8059 19239 -7219
rect 19331 -8059 19333 -7219
rect 19333 -8059 19385 -7219
rect 19385 -8059 19387 -7219
rect 19479 -8059 19481 -7219
rect 19481 -8059 19533 -7219
rect 19533 -8059 19535 -7219
rect 19627 -8059 19629 -7219
rect 19629 -8059 19681 -7219
rect 19681 -8059 19683 -7219
rect 19775 -8059 19777 -7219
rect 19777 -8059 19829 -7219
rect 19829 -8059 19831 -7219
rect 19923 -8059 19925 -7219
rect 19925 -8059 19977 -7219
rect 19977 -8059 19979 -7219
rect 20071 -8059 20073 -7219
rect 20073 -8059 20125 -7219
rect 20125 -8059 20127 -7219
rect 20219 -8059 20221 -7219
rect 20221 -8059 20273 -7219
rect 20273 -8059 20275 -7219
rect 20367 -8059 20369 -7219
rect 20369 -8059 20421 -7219
rect 20421 -8059 20423 -7219
rect 20515 -8059 20517 -7219
rect 20517 -8059 20569 -7219
rect 20569 -8059 20571 -7219
rect 20663 -8059 20665 -7219
rect 20665 -8059 20717 -7219
rect 20717 -8059 20719 -7219
rect 20811 -8059 20813 -7219
rect 20813 -8059 20865 -7219
rect 20865 -8059 20867 -7219
rect 20959 -8059 20961 -7219
rect 20961 -8059 21013 -7219
rect 21013 -8059 21015 -7219
rect 21107 -8059 21109 -7219
rect 21109 -8059 21161 -7219
rect 21161 -8059 21163 -7219
rect 21255 -8059 21257 -7219
rect 21257 -8059 21309 -7219
rect 21309 -8059 21311 -7219
rect 21403 -8059 21405 -7219
rect 21405 -8059 21457 -7219
rect 21457 -8059 21459 -7219
rect 21551 -8059 21553 -7219
rect 21553 -8059 21605 -7219
rect 21605 -8059 21607 -7219
rect 21699 -8059 21701 -7219
rect 21701 -8059 21753 -7219
rect 21753 -8059 21755 -7219
rect 21847 -8059 21849 -7219
rect 21849 -8059 21901 -7219
rect 21901 -8059 21903 -7219
rect 21995 -8059 21997 -7219
rect 21997 -8059 22049 -7219
rect 22049 -8059 22051 -7219
rect 22143 -8059 22145 -7219
rect 22145 -8059 22197 -7219
rect 22197 -8059 22199 -7219
rect 22291 -8059 22293 -7219
rect 22293 -8059 22345 -7219
rect 22345 -8059 22347 -7219
rect 22439 -8059 22441 -7219
rect 22441 -8059 22493 -7219
rect 22493 -8059 22495 -7219
rect 22587 -8059 22589 -7219
rect 22589 -8059 22641 -7219
rect 22641 -8059 22643 -7219
rect 22735 -8059 22737 -7219
rect 22737 -8059 22789 -7219
rect 22789 -8059 22791 -7219
rect 22883 -8059 22885 -7219
rect 22885 -8059 22937 -7219
rect 22937 -8059 22939 -7219
rect 23031 -8059 23033 -7219
rect 23033 -8059 23085 -7219
rect 23085 -8059 23087 -7219
rect 23179 -8059 23181 -7219
rect 23181 -8059 23233 -7219
rect 23233 -8059 23235 -7219
rect 23327 -8059 23329 -7219
rect 23329 -8059 23381 -7219
rect 23381 -8059 23383 -7219
rect 23475 -8059 23477 -7219
rect 23477 -8059 23529 -7219
rect 23529 -8059 23531 -7219
rect 23623 -8059 23625 -7219
rect 23625 -8059 23677 -7219
rect 23677 -8059 23679 -7219
rect 10834 -8284 10890 -8228
rect 10915 -8284 10971 -8228
rect 10996 -8284 11052 -8228
rect 11077 -8284 11133 -8228
rect 11158 -8284 11214 -8228
rect 11239 -8284 11295 -8228
rect 11320 -8284 11376 -8228
rect 11401 -8284 11457 -8228
rect 11482 -8284 11538 -8228
rect 11563 -8284 11619 -8228
rect 11644 -8284 11700 -8228
rect 11725 -8284 11781 -8228
rect 11806 -8284 11862 -8228
rect 10834 -8388 10890 -8332
rect 10915 -8388 10971 -8332
rect 10996 -8388 11052 -8332
rect 11077 -8388 11133 -8332
rect 11158 -8388 11214 -8332
rect 11239 -8388 11295 -8332
rect 11320 -8388 11376 -8332
rect 11401 -8388 11457 -8332
rect 11482 -8388 11538 -8332
rect 11563 -8388 11619 -8332
rect 11644 -8388 11700 -8332
rect 11725 -8388 11781 -8332
rect 11806 -8388 11862 -8332
rect 12523 -9205 12525 -8365
rect 12525 -9205 12577 -8365
rect 12577 -9205 12579 -8365
rect 12671 -9205 12673 -8365
rect 12673 -9205 12725 -8365
rect 12725 -9205 12727 -8365
rect 12819 -9205 12821 -8365
rect 12821 -9205 12873 -8365
rect 12873 -9205 12875 -8365
rect 12967 -9205 12969 -8365
rect 12969 -9205 13021 -8365
rect 13021 -9205 13023 -8365
rect 13115 -9205 13117 -8365
rect 13117 -9205 13169 -8365
rect 13169 -9205 13171 -8365
rect 13263 -9205 13265 -8365
rect 13265 -9205 13317 -8365
rect 13317 -9205 13319 -8365
rect 13411 -9205 13413 -8365
rect 13413 -9205 13465 -8365
rect 13465 -9205 13467 -8365
rect 13559 -9205 13561 -8365
rect 13561 -9205 13613 -8365
rect 13613 -9205 13615 -8365
rect 13707 -9205 13709 -8365
rect 13709 -9205 13761 -8365
rect 13761 -9205 13763 -8365
rect 13855 -9205 13857 -8365
rect 13857 -9205 13909 -8365
rect 13909 -9205 13911 -8365
rect 14003 -9205 14005 -8365
rect 14005 -9205 14057 -8365
rect 14057 -9205 14059 -8365
rect 14151 -9205 14153 -8365
rect 14153 -9205 14205 -8365
rect 14205 -9205 14207 -8365
rect 14299 -9205 14301 -8365
rect 14301 -9205 14353 -8365
rect 14353 -9205 14355 -8365
rect 14447 -9205 14449 -8365
rect 14449 -9205 14501 -8365
rect 14501 -9205 14503 -8365
rect 14595 -9205 14597 -8365
rect 14597 -9205 14649 -8365
rect 14649 -9205 14651 -8365
rect 14743 -9205 14745 -8365
rect 14745 -9205 14797 -8365
rect 14797 -9205 14799 -8365
rect 14891 -9205 14893 -8365
rect 14893 -9205 14945 -8365
rect 14945 -9205 14947 -8365
rect 15039 -9205 15041 -8365
rect 15041 -9205 15093 -8365
rect 15093 -9205 15095 -8365
rect 15187 -9205 15189 -8365
rect 15189 -9205 15241 -8365
rect 15241 -9205 15243 -8365
rect 15335 -9205 15337 -8365
rect 15337 -9205 15389 -8365
rect 15389 -9205 15391 -8365
rect 15483 -9205 15485 -8365
rect 15485 -9205 15537 -8365
rect 15537 -9205 15539 -8365
rect 15631 -9205 15633 -8365
rect 15633 -9205 15685 -8365
rect 15685 -9205 15687 -8365
rect 15779 -9205 15781 -8365
rect 15781 -9205 15833 -8365
rect 15833 -9205 15835 -8365
rect 15927 -9205 15929 -8365
rect 15929 -9205 15981 -8365
rect 15981 -9205 15983 -8365
rect 16075 -9205 16077 -8365
rect 16077 -9205 16129 -8365
rect 16129 -9205 16131 -8365
rect 16223 -9205 16225 -8365
rect 16225 -9205 16277 -8365
rect 16277 -9205 16279 -8365
rect 16371 -9205 16373 -8365
rect 16373 -9205 16425 -8365
rect 16425 -9205 16427 -8365
rect 16519 -9205 16521 -8365
rect 16521 -9205 16573 -8365
rect 16573 -9205 16575 -8365
rect 16667 -9205 16669 -8365
rect 16669 -9205 16721 -8365
rect 16721 -9205 16723 -8365
rect 16815 -9205 16817 -8365
rect 16817 -9205 16869 -8365
rect 16869 -9205 16871 -8365
rect 16963 -9205 16965 -8365
rect 16965 -9205 17017 -8365
rect 17017 -9205 17019 -8365
rect 17111 -9205 17113 -8365
rect 17113 -9205 17165 -8365
rect 17165 -9205 17167 -8365
rect 17259 -9205 17261 -8365
rect 17261 -9205 17313 -8365
rect 17313 -9205 17315 -8365
rect 17407 -9205 17409 -8365
rect 17409 -9205 17461 -8365
rect 17461 -9205 17463 -8365
rect 17555 -9205 17557 -8365
rect 17557 -9205 17609 -8365
rect 17609 -9205 17611 -8365
rect 17703 -9205 17705 -8365
rect 17705 -9205 17757 -8365
rect 17757 -9205 17759 -8365
rect 17851 -9205 17853 -8365
rect 17853 -9205 17905 -8365
rect 17905 -9205 17907 -8365
rect 17999 -9205 18001 -8365
rect 18001 -9205 18053 -8365
rect 18053 -9205 18055 -8365
rect 18147 -9205 18149 -8365
rect 18149 -9205 18201 -8365
rect 18201 -9205 18203 -8365
rect 18295 -9205 18297 -8365
rect 18297 -9205 18349 -8365
rect 18349 -9205 18351 -8365
rect 18443 -9205 18445 -8365
rect 18445 -9205 18497 -8365
rect 18497 -9205 18499 -8365
rect 18591 -9205 18593 -8365
rect 18593 -9205 18645 -8365
rect 18645 -9205 18647 -8365
rect 18739 -9205 18741 -8365
rect 18741 -9205 18793 -8365
rect 18793 -9205 18795 -8365
rect 18887 -9205 18889 -8365
rect 18889 -9205 18941 -8365
rect 18941 -9205 18943 -8365
rect 19035 -9205 19037 -8365
rect 19037 -9205 19089 -8365
rect 19089 -9205 19091 -8365
rect 19183 -9205 19185 -8365
rect 19185 -9205 19237 -8365
rect 19237 -9205 19239 -8365
rect 19331 -9205 19333 -8365
rect 19333 -9205 19385 -8365
rect 19385 -9205 19387 -8365
rect 19479 -9205 19481 -8365
rect 19481 -9205 19533 -8365
rect 19533 -9205 19535 -8365
rect 19627 -9205 19629 -8365
rect 19629 -9205 19681 -8365
rect 19681 -9205 19683 -8365
rect 19775 -9205 19777 -8365
rect 19777 -9205 19829 -8365
rect 19829 -9205 19831 -8365
rect 19923 -9205 19925 -8365
rect 19925 -9205 19977 -8365
rect 19977 -9205 19979 -8365
rect 20071 -9205 20073 -8365
rect 20073 -9205 20125 -8365
rect 20125 -9205 20127 -8365
rect 20219 -9205 20221 -8365
rect 20221 -9205 20273 -8365
rect 20273 -9205 20275 -8365
rect 20367 -9205 20369 -8365
rect 20369 -9205 20421 -8365
rect 20421 -9205 20423 -8365
rect 20515 -9205 20517 -8365
rect 20517 -9205 20569 -8365
rect 20569 -9205 20571 -8365
rect 20663 -9205 20665 -8365
rect 20665 -9205 20717 -8365
rect 20717 -9205 20719 -8365
rect 20811 -9205 20813 -8365
rect 20813 -9205 20865 -8365
rect 20865 -9205 20867 -8365
rect 20959 -9205 20961 -8365
rect 20961 -9205 21013 -8365
rect 21013 -9205 21015 -8365
rect 21107 -9205 21109 -8365
rect 21109 -9205 21161 -8365
rect 21161 -9205 21163 -8365
rect 21255 -9205 21257 -8365
rect 21257 -9205 21309 -8365
rect 21309 -9205 21311 -8365
rect 21403 -9205 21405 -8365
rect 21405 -9205 21457 -8365
rect 21457 -9205 21459 -8365
rect 21551 -9205 21553 -8365
rect 21553 -9205 21605 -8365
rect 21605 -9205 21607 -8365
rect 21699 -9205 21701 -8365
rect 21701 -9205 21753 -8365
rect 21753 -9205 21755 -8365
rect 21847 -9205 21849 -8365
rect 21849 -9205 21901 -8365
rect 21901 -9205 21903 -8365
rect 21995 -9205 21997 -8365
rect 21997 -9205 22049 -8365
rect 22049 -9205 22051 -8365
rect 22143 -9205 22145 -8365
rect 22145 -9205 22197 -8365
rect 22197 -9205 22199 -8365
rect 22291 -9205 22293 -8365
rect 22293 -9205 22345 -8365
rect 22345 -9205 22347 -8365
rect 22439 -9205 22441 -8365
rect 22441 -9205 22493 -8365
rect 22493 -9205 22495 -8365
rect 22587 -9205 22589 -8365
rect 22589 -9205 22641 -8365
rect 22641 -9205 22643 -8365
rect 22735 -9205 22737 -8365
rect 22737 -9205 22789 -8365
rect 22789 -9205 22791 -8365
rect 22883 -9205 22885 -8365
rect 22885 -9205 22937 -8365
rect 22937 -9205 22939 -8365
rect 23031 -9205 23033 -8365
rect 23033 -9205 23085 -8365
rect 23085 -9205 23087 -8365
rect 23179 -9205 23181 -8365
rect 23181 -9205 23233 -8365
rect 23233 -9205 23235 -8365
rect 23327 -9205 23329 -8365
rect 23329 -9205 23381 -8365
rect 23381 -9205 23383 -8365
rect 23475 -9205 23477 -8365
rect 23477 -9205 23529 -8365
rect 23529 -9205 23531 -8365
rect 23623 -9205 23625 -8365
rect 23625 -9205 23677 -8365
rect 23677 -9205 23679 -8365
rect 4053 -9683 4109 -9681
rect 4053 -9735 4055 -9683
rect 4055 -9735 4107 -9683
rect 4107 -9735 4109 -9683
rect 4053 -9737 4109 -9735
rect 4134 -9683 4190 -9681
rect 4134 -9735 4136 -9683
rect 4136 -9735 4188 -9683
rect 4188 -9735 4190 -9683
rect 4134 -9737 4190 -9735
rect 4215 -9683 4271 -9681
rect 4215 -9735 4217 -9683
rect 4217 -9735 4269 -9683
rect 4269 -9735 4271 -9683
rect 4215 -9737 4271 -9735
rect 4296 -9683 4352 -9681
rect 4296 -9735 4298 -9683
rect 4298 -9735 4350 -9683
rect 4350 -9735 4352 -9683
rect 4296 -9737 4352 -9735
rect 4377 -9683 4433 -9681
rect 4377 -9735 4379 -9683
rect 4379 -9735 4431 -9683
rect 4431 -9735 4433 -9683
rect 4377 -9737 4433 -9735
rect 4458 -9683 4514 -9681
rect 4458 -9735 4460 -9683
rect 4460 -9735 4512 -9683
rect 4512 -9735 4514 -9683
rect 4458 -9737 4514 -9735
rect 4539 -9683 4595 -9681
rect 4539 -9735 4541 -9683
rect 4541 -9735 4593 -9683
rect 4593 -9735 4595 -9683
rect 4539 -9737 4595 -9735
rect 4621 -9683 4677 -9681
rect 4621 -9735 4623 -9683
rect 4623 -9735 4675 -9683
rect 4675 -9735 4677 -9683
rect 4621 -9737 4677 -9735
rect 4702 -9683 4758 -9681
rect 4702 -9735 4704 -9683
rect 4704 -9735 4756 -9683
rect 4756 -9735 4758 -9683
rect 4702 -9737 4758 -9735
rect 4783 -9683 4839 -9681
rect 4783 -9735 4785 -9683
rect 4785 -9735 4837 -9683
rect 4837 -9735 4839 -9683
rect 4783 -9737 4839 -9735
rect 4864 -9683 4920 -9681
rect 4864 -9735 4866 -9683
rect 4866 -9735 4918 -9683
rect 4918 -9735 4920 -9683
rect 4864 -9737 4920 -9735
rect 4945 -9683 5001 -9681
rect 4945 -9735 4947 -9683
rect 4947 -9735 4999 -9683
rect 4999 -9735 5001 -9683
rect 4945 -9737 5001 -9735
rect 5026 -9683 5082 -9681
rect 5026 -9735 5028 -9683
rect 5028 -9735 5080 -9683
rect 5080 -9735 5082 -9683
rect 5026 -9737 5082 -9735
rect 5107 -9683 5163 -9681
rect 5107 -9735 5109 -9683
rect 5109 -9735 5161 -9683
rect 5161 -9735 5163 -9683
rect 5107 -9737 5163 -9735
rect 5189 -9683 5245 -9681
rect 5189 -9735 5191 -9683
rect 5191 -9735 5243 -9683
rect 5243 -9735 5245 -9683
rect 5189 -9737 5245 -9735
rect 5270 -9683 5326 -9681
rect 5270 -9735 5272 -9683
rect 5272 -9735 5324 -9683
rect 5324 -9735 5326 -9683
rect 5270 -9737 5326 -9735
rect 5351 -9683 5407 -9681
rect 5351 -9735 5353 -9683
rect 5353 -9735 5405 -9683
rect 5405 -9735 5407 -9683
rect 5351 -9737 5407 -9735
rect 5432 -9683 5488 -9681
rect 5432 -9735 5434 -9683
rect 5434 -9735 5486 -9683
rect 5486 -9735 5488 -9683
rect 5432 -9737 5488 -9735
rect 5513 -9683 5569 -9681
rect 5513 -9735 5515 -9683
rect 5515 -9735 5567 -9683
rect 5567 -9735 5569 -9683
rect 5513 -9737 5569 -9735
rect 5594 -9683 5650 -9681
rect 5594 -9735 5596 -9683
rect 5596 -9735 5648 -9683
rect 5648 -9735 5650 -9683
rect 5594 -9737 5650 -9735
rect 5675 -9683 5731 -9681
rect 5675 -9735 5677 -9683
rect 5677 -9735 5729 -9683
rect 5729 -9735 5731 -9683
rect 5675 -9737 5731 -9735
rect 5757 -9683 5813 -9681
rect 5757 -9735 5759 -9683
rect 5759 -9735 5811 -9683
rect 5811 -9735 5813 -9683
rect 5757 -9737 5813 -9735
rect 5838 -9683 5894 -9681
rect 5838 -9735 5840 -9683
rect 5840 -9735 5892 -9683
rect 5892 -9735 5894 -9683
rect 5838 -9737 5894 -9735
rect 5919 -9683 5975 -9681
rect 5919 -9735 5921 -9683
rect 5921 -9735 5973 -9683
rect 5973 -9735 5975 -9683
rect 5919 -9737 5975 -9735
rect 6000 -9683 6056 -9681
rect 6000 -9735 6002 -9683
rect 6002 -9735 6054 -9683
rect 6054 -9735 6056 -9683
rect 6000 -9737 6056 -9735
rect 6081 -9683 6137 -9681
rect 6081 -9735 6083 -9683
rect 6083 -9735 6135 -9683
rect 6135 -9735 6137 -9683
rect 6081 -9737 6137 -9735
rect 6162 -9683 6218 -9681
rect 6162 -9735 6164 -9683
rect 6164 -9735 6216 -9683
rect 6216 -9735 6218 -9683
rect 6162 -9737 6218 -9735
rect 6243 -9683 6299 -9681
rect 6243 -9735 6245 -9683
rect 6245 -9735 6297 -9683
rect 6297 -9735 6299 -9683
rect 6243 -9737 6299 -9735
rect 6325 -9683 6381 -9681
rect 6325 -9735 6327 -9683
rect 6327 -9735 6379 -9683
rect 6379 -9735 6381 -9683
rect 6325 -9737 6381 -9735
rect 6406 -9683 6462 -9681
rect 6406 -9735 6408 -9683
rect 6408 -9735 6460 -9683
rect 6460 -9735 6462 -9683
rect 6406 -9737 6462 -9735
rect 6487 -9683 6543 -9681
rect 6487 -9735 6489 -9683
rect 6489 -9735 6541 -9683
rect 6541 -9735 6543 -9683
rect 6487 -9737 6543 -9735
rect 6568 -9683 6624 -9681
rect 6568 -9735 6570 -9683
rect 6570 -9735 6622 -9683
rect 6622 -9735 6624 -9683
rect 6568 -9737 6624 -9735
rect 6649 -9683 6705 -9681
rect 6649 -9735 6651 -9683
rect 6651 -9735 6703 -9683
rect 6703 -9735 6705 -9683
rect 6649 -9737 6705 -9735
rect 6730 -9683 6786 -9681
rect 6730 -9735 6732 -9683
rect 6732 -9735 6784 -9683
rect 6784 -9735 6786 -9683
rect 6730 -9737 6786 -9735
rect 6811 -9683 6867 -9681
rect 6811 -9735 6813 -9683
rect 6813 -9735 6865 -9683
rect 6865 -9735 6867 -9683
rect 6811 -9737 6867 -9735
rect 6893 -9683 6949 -9681
rect 6893 -9735 6895 -9683
rect 6895 -9735 6947 -9683
rect 6947 -9735 6949 -9683
rect 6893 -9737 6949 -9735
rect 6974 -9683 7030 -9681
rect 6974 -9735 6976 -9683
rect 6976 -9735 7028 -9683
rect 7028 -9735 7030 -9683
rect 6974 -9737 7030 -9735
rect 7055 -9683 7111 -9681
rect 7055 -9735 7057 -9683
rect 7057 -9735 7109 -9683
rect 7109 -9735 7111 -9683
rect 7055 -9737 7111 -9735
rect 7136 -9683 7192 -9681
rect 7136 -9735 7138 -9683
rect 7138 -9735 7190 -9683
rect 7190 -9735 7192 -9683
rect 7136 -9737 7192 -9735
rect 7217 -9683 7273 -9681
rect 7217 -9735 7219 -9683
rect 7219 -9735 7271 -9683
rect 7271 -9735 7273 -9683
rect 7217 -9737 7273 -9735
rect 7298 -9683 7354 -9681
rect 7298 -9735 7300 -9683
rect 7300 -9735 7352 -9683
rect 7352 -9735 7354 -9683
rect 7298 -9737 7354 -9735
rect 7379 -9683 7435 -9681
rect 7379 -9735 7381 -9683
rect 7381 -9735 7433 -9683
rect 7433 -9735 7435 -9683
rect 7379 -9737 7435 -9735
rect 7461 -9683 7517 -9681
rect 7461 -9735 7463 -9683
rect 7463 -9735 7515 -9683
rect 7515 -9735 7517 -9683
rect 7461 -9737 7517 -9735
rect 7542 -9683 7598 -9681
rect 7542 -9735 7544 -9683
rect 7544 -9735 7596 -9683
rect 7596 -9735 7598 -9683
rect 7542 -9737 7598 -9735
rect 7623 -9683 7679 -9681
rect 7623 -9735 7625 -9683
rect 7625 -9735 7677 -9683
rect 7677 -9735 7679 -9683
rect 7623 -9737 7679 -9735
rect 7704 -9683 7760 -9681
rect 7704 -9735 7706 -9683
rect 7706 -9735 7758 -9683
rect 7758 -9735 7760 -9683
rect 7704 -9737 7760 -9735
rect 7785 -9683 7841 -9681
rect 7785 -9735 7787 -9683
rect 7787 -9735 7839 -9683
rect 7839 -9735 7841 -9683
rect 7785 -9737 7841 -9735
rect 7866 -9683 7922 -9681
rect 7866 -9735 7868 -9683
rect 7868 -9735 7920 -9683
rect 7920 -9735 7922 -9683
rect 7866 -9737 7922 -9735
rect 7947 -9683 8003 -9681
rect 7947 -9735 7949 -9683
rect 7949 -9735 8001 -9683
rect 8001 -9735 8003 -9683
rect 7947 -9737 8003 -9735
rect 8029 -9683 8085 -9681
rect 8029 -9735 8031 -9683
rect 8031 -9735 8083 -9683
rect 8083 -9735 8085 -9683
rect 8029 -9737 8085 -9735
rect 8110 -9683 8166 -9681
rect 8110 -9735 8112 -9683
rect 8112 -9735 8164 -9683
rect 8164 -9735 8166 -9683
rect 8110 -9737 8166 -9735
rect 8191 -9683 8247 -9681
rect 8191 -9735 8193 -9683
rect 8193 -9735 8245 -9683
rect 8245 -9735 8247 -9683
rect 8191 -9737 8247 -9735
rect 8272 -9683 8328 -9681
rect 8272 -9735 8274 -9683
rect 8274 -9735 8326 -9683
rect 8326 -9735 8328 -9683
rect 8272 -9737 8328 -9735
rect 8353 -9683 8409 -9681
rect 8353 -9735 8355 -9683
rect 8355 -9735 8407 -9683
rect 8407 -9735 8409 -9683
rect 8353 -9737 8409 -9735
rect 8434 -9683 8490 -9681
rect 8434 -9735 8436 -9683
rect 8436 -9735 8488 -9683
rect 8488 -9735 8490 -9683
rect 8434 -9737 8490 -9735
rect 8515 -9683 8571 -9681
rect 8515 -9735 8517 -9683
rect 8517 -9735 8569 -9683
rect 8569 -9735 8571 -9683
rect 8515 -9737 8571 -9735
rect 8597 -9683 8653 -9681
rect 8597 -9735 8599 -9683
rect 8599 -9735 8651 -9683
rect 8651 -9735 8653 -9683
rect 8597 -9737 8653 -9735
rect 8678 -9683 8734 -9681
rect 8678 -9735 8680 -9683
rect 8680 -9735 8732 -9683
rect 8732 -9735 8734 -9683
rect 8678 -9737 8734 -9735
rect 8759 -9683 8815 -9681
rect 8759 -9735 8761 -9683
rect 8761 -9735 8813 -9683
rect 8813 -9735 8815 -9683
rect 8759 -9737 8815 -9735
rect 8840 -9683 8896 -9681
rect 8840 -9735 8842 -9683
rect 8842 -9735 8894 -9683
rect 8894 -9735 8896 -9683
rect 8840 -9737 8896 -9735
rect 8921 -9683 8977 -9681
rect 8921 -9735 8923 -9683
rect 8923 -9735 8975 -9683
rect 8975 -9735 8977 -9683
rect 8921 -9737 8977 -9735
rect 9002 -9683 9058 -9681
rect 9002 -9735 9004 -9683
rect 9004 -9735 9056 -9683
rect 9056 -9735 9058 -9683
rect 9002 -9737 9058 -9735
rect 9083 -9683 9139 -9681
rect 9083 -9735 9085 -9683
rect 9085 -9735 9137 -9683
rect 9137 -9735 9139 -9683
rect 9083 -9737 9139 -9735
rect 9165 -9683 9221 -9681
rect 9165 -9735 9167 -9683
rect 9167 -9735 9219 -9683
rect 9219 -9735 9221 -9683
rect 9165 -9737 9221 -9735
rect 9246 -9683 9302 -9681
rect 9246 -9735 9248 -9683
rect 9248 -9735 9300 -9683
rect 9300 -9735 9302 -9683
rect 9246 -9737 9302 -9735
rect 9327 -9683 9383 -9681
rect 9327 -9735 9329 -9683
rect 9329 -9735 9381 -9683
rect 9381 -9735 9383 -9683
rect 9327 -9737 9383 -9735
rect 9408 -9683 9464 -9681
rect 9408 -9735 9410 -9683
rect 9410 -9735 9462 -9683
rect 9462 -9735 9464 -9683
rect 9408 -9737 9464 -9735
rect 9489 -9683 9545 -9681
rect 9489 -9735 9491 -9683
rect 9491 -9735 9543 -9683
rect 9543 -9735 9545 -9683
rect 9489 -9737 9545 -9735
rect 9570 -9683 9626 -9681
rect 9570 -9735 9572 -9683
rect 9572 -9735 9624 -9683
rect 9624 -9735 9626 -9683
rect 9570 -9737 9626 -9735
rect 9651 -9683 9707 -9681
rect 9651 -9735 9653 -9683
rect 9653 -9735 9705 -9683
rect 9705 -9735 9707 -9683
rect 9651 -9737 9707 -9735
rect 9733 -9683 9789 -9681
rect 9733 -9735 9735 -9683
rect 9735 -9735 9787 -9683
rect 9787 -9735 9789 -9683
rect 9733 -9737 9789 -9735
rect 9814 -9683 9870 -9681
rect 9814 -9735 9816 -9683
rect 9816 -9735 9868 -9683
rect 9868 -9735 9870 -9683
rect 9814 -9737 9870 -9735
rect 9895 -9683 9951 -9681
rect 9895 -9735 9897 -9683
rect 9897 -9735 9949 -9683
rect 9949 -9735 9951 -9683
rect 9895 -9737 9951 -9735
rect 9976 -9683 10032 -9681
rect 9976 -9735 9978 -9683
rect 9978 -9735 10030 -9683
rect 10030 -9735 10032 -9683
rect 9976 -9737 10032 -9735
rect 10057 -9683 10113 -9681
rect 10057 -9735 10059 -9683
rect 10059 -9735 10111 -9683
rect 10111 -9735 10113 -9683
rect 10057 -9737 10113 -9735
rect 10138 -9683 10194 -9681
rect 10138 -9735 10140 -9683
rect 10140 -9735 10192 -9683
rect 10192 -9735 10194 -9683
rect 10138 -9737 10194 -9735
rect 10219 -9683 10275 -9681
rect 10219 -9735 10221 -9683
rect 10221 -9735 10273 -9683
rect 10273 -9735 10275 -9683
rect 10219 -9737 10275 -9735
rect 10301 -9683 10357 -9681
rect 10301 -9735 10303 -9683
rect 10303 -9735 10355 -9683
rect 10355 -9735 10357 -9683
rect 10301 -9737 10357 -9735
rect 10382 -9683 10438 -9681
rect 10382 -9735 10384 -9683
rect 10384 -9735 10436 -9683
rect 10436 -9735 10438 -9683
rect 10382 -9737 10438 -9735
rect 10463 -9683 10519 -9681
rect 10463 -9735 10465 -9683
rect 10465 -9735 10517 -9683
rect 10517 -9735 10519 -9683
rect 10463 -9737 10519 -9735
rect 10544 -9683 10600 -9681
rect 10544 -9735 10546 -9683
rect 10546 -9735 10598 -9683
rect 10598 -9735 10600 -9683
rect 10544 -9737 10600 -9735
rect 10625 -9683 10681 -9681
rect 10625 -9735 10627 -9683
rect 10627 -9735 10679 -9683
rect 10679 -9735 10681 -9683
rect 10625 -9737 10681 -9735
rect 10706 -9683 10762 -9681
rect 10706 -9735 10708 -9683
rect 10708 -9735 10760 -9683
rect 10760 -9735 10762 -9683
rect 10706 -9737 10762 -9735
rect 10787 -9683 10843 -9681
rect 10787 -9735 10789 -9683
rect 10789 -9735 10841 -9683
rect 10841 -9735 10843 -9683
rect 10787 -9737 10843 -9735
rect 10869 -9683 10925 -9681
rect 10869 -9735 10871 -9683
rect 10871 -9735 10923 -9683
rect 10923 -9735 10925 -9683
rect 10869 -9737 10925 -9735
rect 10950 -9683 11006 -9681
rect 10950 -9735 10952 -9683
rect 10952 -9735 11004 -9683
rect 11004 -9735 11006 -9683
rect 10950 -9737 11006 -9735
rect 11031 -9683 11087 -9681
rect 11031 -9735 11033 -9683
rect 11033 -9735 11085 -9683
rect 11085 -9735 11087 -9683
rect 11031 -9737 11087 -9735
rect 11112 -9683 11168 -9681
rect 11112 -9735 11114 -9683
rect 11114 -9735 11166 -9683
rect 11166 -9735 11168 -9683
rect 11112 -9737 11168 -9735
rect 11193 -9683 11249 -9681
rect 11193 -9735 11195 -9683
rect 11195 -9735 11247 -9683
rect 11247 -9735 11249 -9683
rect 11193 -9737 11249 -9735
rect 11274 -9683 11330 -9681
rect 11274 -9735 11276 -9683
rect 11276 -9735 11328 -9683
rect 11328 -9735 11330 -9683
rect 11274 -9737 11330 -9735
rect 11355 -9683 11411 -9681
rect 11355 -9735 11357 -9683
rect 11357 -9735 11409 -9683
rect 11409 -9735 11411 -9683
rect 11355 -9737 11411 -9735
rect 11437 -9683 11493 -9681
rect 11437 -9735 11439 -9683
rect 11439 -9735 11491 -9683
rect 11491 -9735 11493 -9683
rect 11437 -9737 11493 -9735
rect 11518 -9683 11574 -9681
rect 11518 -9735 11520 -9683
rect 11520 -9735 11572 -9683
rect 11572 -9735 11574 -9683
rect 11518 -9737 11574 -9735
rect 11599 -9683 11655 -9681
rect 11599 -9735 11601 -9683
rect 11601 -9735 11653 -9683
rect 11653 -9735 11655 -9683
rect 11599 -9737 11655 -9735
rect 11680 -9683 11736 -9681
rect 11680 -9735 11682 -9683
rect 11682 -9735 11734 -9683
rect 11734 -9735 11736 -9683
rect 11680 -9737 11736 -9735
rect 11761 -9683 11817 -9681
rect 11761 -9735 11763 -9683
rect 11763 -9735 11815 -9683
rect 11815 -9735 11817 -9683
rect 11761 -9737 11817 -9735
rect 11842 -9683 11898 -9681
rect 11842 -9735 11844 -9683
rect 11844 -9735 11896 -9683
rect 11896 -9735 11898 -9683
rect 11842 -9737 11898 -9735
rect 11923 -9683 11979 -9681
rect 11923 -9735 11925 -9683
rect 11925 -9735 11977 -9683
rect 11977 -9735 11979 -9683
rect 11923 -9737 11979 -9735
rect 12005 -9683 12061 -9681
rect 12005 -9735 12007 -9683
rect 12007 -9735 12059 -9683
rect 12059 -9735 12061 -9683
rect 12005 -9737 12061 -9735
rect 12086 -9683 12142 -9681
rect 12086 -9735 12088 -9683
rect 12088 -9735 12140 -9683
rect 12140 -9735 12142 -9683
rect 12086 -9737 12142 -9735
rect 12167 -9683 12223 -9681
rect 12167 -9735 12169 -9683
rect 12169 -9735 12221 -9683
rect 12221 -9735 12223 -9683
rect 12167 -9737 12223 -9735
rect 12248 -9683 12304 -9681
rect 12248 -9735 12250 -9683
rect 12250 -9735 12302 -9683
rect 12302 -9735 12304 -9683
rect 12248 -9737 12304 -9735
rect 12329 -9683 12385 -9681
rect 12329 -9735 12331 -9683
rect 12331 -9735 12383 -9683
rect 12383 -9735 12385 -9683
rect 12329 -9737 12385 -9735
rect 12410 -9683 12466 -9681
rect 12410 -9735 12412 -9683
rect 12412 -9735 12464 -9683
rect 12464 -9735 12466 -9683
rect 12410 -9737 12466 -9735
rect 12491 -9683 12547 -9681
rect 12491 -9735 12493 -9683
rect 12493 -9735 12545 -9683
rect 12545 -9735 12547 -9683
rect 12491 -9737 12547 -9735
rect 12573 -9683 12629 -9681
rect 12573 -9735 12575 -9683
rect 12575 -9735 12627 -9683
rect 12627 -9735 12629 -9683
rect 12573 -9737 12629 -9735
rect 12654 -9683 12710 -9681
rect 12654 -9735 12656 -9683
rect 12656 -9735 12708 -9683
rect 12708 -9735 12710 -9683
rect 12654 -9737 12710 -9735
rect 12735 -9683 12791 -9681
rect 12735 -9735 12737 -9683
rect 12737 -9735 12789 -9683
rect 12789 -9735 12791 -9683
rect 12735 -9737 12791 -9735
rect 12816 -9683 12872 -9681
rect 12816 -9735 12818 -9683
rect 12818 -9735 12870 -9683
rect 12870 -9735 12872 -9683
rect 12816 -9737 12872 -9735
rect 12897 -9683 12953 -9681
rect 12897 -9735 12899 -9683
rect 12899 -9735 12951 -9683
rect 12951 -9735 12953 -9683
rect 12897 -9737 12953 -9735
rect 12978 -9683 13034 -9681
rect 12978 -9735 12980 -9683
rect 12980 -9735 13032 -9683
rect 13032 -9735 13034 -9683
rect 12978 -9737 13034 -9735
rect 13059 -9683 13115 -9681
rect 13059 -9735 13061 -9683
rect 13061 -9735 13113 -9683
rect 13113 -9735 13115 -9683
rect 13059 -9737 13115 -9735
rect 13141 -9683 13197 -9681
rect 13141 -9735 13143 -9683
rect 13143 -9735 13195 -9683
rect 13195 -9735 13197 -9683
rect 13141 -9737 13197 -9735
rect 13222 -9683 13278 -9681
rect 13222 -9735 13224 -9683
rect 13224 -9735 13276 -9683
rect 13276 -9735 13278 -9683
rect 13222 -9737 13278 -9735
rect 13303 -9683 13359 -9681
rect 13303 -9735 13305 -9683
rect 13305 -9735 13357 -9683
rect 13357 -9735 13359 -9683
rect 13303 -9737 13359 -9735
rect 13384 -9683 13440 -9681
rect 13384 -9735 13386 -9683
rect 13386 -9735 13438 -9683
rect 13438 -9735 13440 -9683
rect 13384 -9737 13440 -9735
rect 13465 -9683 13521 -9681
rect 13465 -9735 13467 -9683
rect 13467 -9735 13519 -9683
rect 13519 -9735 13521 -9683
rect 13465 -9737 13521 -9735
rect 13546 -9683 13602 -9681
rect 13546 -9735 13548 -9683
rect 13548 -9735 13600 -9683
rect 13600 -9735 13602 -9683
rect 13546 -9737 13602 -9735
rect 13627 -9683 13683 -9681
rect 13627 -9735 13629 -9683
rect 13629 -9735 13681 -9683
rect 13681 -9735 13683 -9683
rect 13627 -9737 13683 -9735
rect 13709 -9683 13765 -9681
rect 13709 -9735 13711 -9683
rect 13711 -9735 13763 -9683
rect 13763 -9735 13765 -9683
rect 13709 -9737 13765 -9735
rect 13790 -9683 13846 -9681
rect 13790 -9735 13792 -9683
rect 13792 -9735 13844 -9683
rect 13844 -9735 13846 -9683
rect 13790 -9737 13846 -9735
rect 13871 -9683 13927 -9681
rect 13871 -9735 13873 -9683
rect 13873 -9735 13925 -9683
rect 13925 -9735 13927 -9683
rect 13871 -9737 13927 -9735
rect 13952 -9683 14008 -9681
rect 13952 -9735 13954 -9683
rect 13954 -9735 14006 -9683
rect 14006 -9735 14008 -9683
rect 13952 -9737 14008 -9735
rect 14033 -9683 14089 -9681
rect 14033 -9735 14035 -9683
rect 14035 -9735 14087 -9683
rect 14087 -9735 14089 -9683
rect 14033 -9737 14089 -9735
rect 14114 -9683 14170 -9681
rect 14114 -9735 14116 -9683
rect 14116 -9735 14168 -9683
rect 14168 -9735 14170 -9683
rect 14114 -9737 14170 -9735
rect 14195 -9683 14251 -9681
rect 14195 -9735 14197 -9683
rect 14197 -9735 14249 -9683
rect 14249 -9735 14251 -9683
rect 14195 -9737 14251 -9735
rect 14277 -9683 14333 -9681
rect 14277 -9735 14279 -9683
rect 14279 -9735 14331 -9683
rect 14331 -9735 14333 -9683
rect 14277 -9737 14333 -9735
rect 14358 -9683 14414 -9681
rect 14358 -9735 14360 -9683
rect 14360 -9735 14412 -9683
rect 14412 -9735 14414 -9683
rect 14358 -9737 14414 -9735
rect 14439 -9683 14495 -9681
rect 14439 -9735 14441 -9683
rect 14441 -9735 14493 -9683
rect 14493 -9735 14495 -9683
rect 14439 -9737 14495 -9735
rect 14520 -9683 14576 -9681
rect 14520 -9735 14522 -9683
rect 14522 -9735 14574 -9683
rect 14574 -9735 14576 -9683
rect 14520 -9737 14576 -9735
rect 14601 -9683 14657 -9681
rect 14601 -9735 14603 -9683
rect 14603 -9735 14655 -9683
rect 14655 -9735 14657 -9683
rect 14601 -9737 14657 -9735
rect 14682 -9683 14738 -9681
rect 14682 -9735 14684 -9683
rect 14684 -9735 14736 -9683
rect 14736 -9735 14738 -9683
rect 14682 -9737 14738 -9735
rect 14763 -9683 14819 -9681
rect 14763 -9735 14765 -9683
rect 14765 -9735 14817 -9683
rect 14817 -9735 14819 -9683
rect 14763 -9737 14819 -9735
rect 14845 -9683 14901 -9681
rect 14845 -9735 14847 -9683
rect 14847 -9735 14899 -9683
rect 14899 -9735 14901 -9683
rect 14845 -9737 14901 -9735
rect 14926 -9683 14982 -9681
rect 14926 -9735 14928 -9683
rect 14928 -9735 14980 -9683
rect 14980 -9735 14982 -9683
rect 14926 -9737 14982 -9735
rect 15007 -9683 15063 -9681
rect 15007 -9735 15009 -9683
rect 15009 -9735 15061 -9683
rect 15061 -9735 15063 -9683
rect 15007 -9737 15063 -9735
rect 15088 -9683 15144 -9681
rect 15088 -9735 15090 -9683
rect 15090 -9735 15142 -9683
rect 15142 -9735 15144 -9683
rect 15088 -9737 15144 -9735
rect 15169 -9683 15225 -9681
rect 15169 -9735 15171 -9683
rect 15171 -9735 15223 -9683
rect 15223 -9735 15225 -9683
rect 15169 -9737 15225 -9735
rect 15250 -9683 15306 -9681
rect 15250 -9735 15252 -9683
rect 15252 -9735 15304 -9683
rect 15304 -9735 15306 -9683
rect 15250 -9737 15306 -9735
rect 15331 -9683 15387 -9681
rect 15331 -9735 15333 -9683
rect 15333 -9735 15385 -9683
rect 15385 -9735 15387 -9683
rect 15331 -9737 15387 -9735
rect 15413 -9683 15469 -9681
rect 15413 -9735 15415 -9683
rect 15415 -9735 15467 -9683
rect 15467 -9735 15469 -9683
rect 15413 -9737 15469 -9735
rect 15494 -9683 15550 -9681
rect 15494 -9735 15496 -9683
rect 15496 -9735 15548 -9683
rect 15548 -9735 15550 -9683
rect 15494 -9737 15550 -9735
rect 15575 -9683 15631 -9681
rect 15575 -9735 15577 -9683
rect 15577 -9735 15629 -9683
rect 15629 -9735 15631 -9683
rect 15575 -9737 15631 -9735
rect 15656 -9683 15712 -9681
rect 15656 -9735 15658 -9683
rect 15658 -9735 15710 -9683
rect 15710 -9735 15712 -9683
rect 15656 -9737 15712 -9735
rect 15737 -9683 15793 -9681
rect 15737 -9735 15739 -9683
rect 15739 -9735 15791 -9683
rect 15791 -9735 15793 -9683
rect 15737 -9737 15793 -9735
rect 15818 -9683 15874 -9681
rect 15818 -9735 15820 -9683
rect 15820 -9735 15872 -9683
rect 15872 -9735 15874 -9683
rect 15818 -9737 15874 -9735
rect 15899 -9683 15955 -9681
rect 15899 -9735 15901 -9683
rect 15901 -9735 15953 -9683
rect 15953 -9735 15955 -9683
rect 15899 -9737 15955 -9735
rect 15981 -9683 16037 -9681
rect 15981 -9735 15983 -9683
rect 15983 -9735 16035 -9683
rect 16035 -9735 16037 -9683
rect 15981 -9737 16037 -9735
rect 16062 -9683 16118 -9681
rect 16062 -9735 16064 -9683
rect 16064 -9735 16116 -9683
rect 16116 -9735 16118 -9683
rect 16062 -9737 16118 -9735
rect 16143 -9683 16199 -9681
rect 16143 -9735 16145 -9683
rect 16145 -9735 16197 -9683
rect 16197 -9735 16199 -9683
rect 16143 -9737 16199 -9735
rect 16224 -9683 16280 -9681
rect 16224 -9735 16226 -9683
rect 16226 -9735 16278 -9683
rect 16278 -9735 16280 -9683
rect 16224 -9737 16280 -9735
rect 16305 -9683 16361 -9681
rect 16305 -9735 16307 -9683
rect 16307 -9735 16359 -9683
rect 16359 -9735 16361 -9683
rect 16305 -9737 16361 -9735
rect 16386 -9683 16442 -9681
rect 16386 -9735 16388 -9683
rect 16388 -9735 16440 -9683
rect 16440 -9735 16442 -9683
rect 16386 -9737 16442 -9735
rect 16467 -9683 16523 -9681
rect 16467 -9735 16469 -9683
rect 16469 -9735 16521 -9683
rect 16521 -9735 16523 -9683
rect 16467 -9737 16523 -9735
rect 16549 -9683 16605 -9681
rect 16549 -9735 16551 -9683
rect 16551 -9735 16603 -9683
rect 16603 -9735 16605 -9683
rect 16549 -9737 16605 -9735
rect 16630 -9683 16686 -9681
rect 16630 -9735 16632 -9683
rect 16632 -9735 16684 -9683
rect 16684 -9735 16686 -9683
rect 16630 -9737 16686 -9735
rect 16711 -9683 16767 -9681
rect 16711 -9735 16713 -9683
rect 16713 -9735 16765 -9683
rect 16765 -9735 16767 -9683
rect 16711 -9737 16767 -9735
rect 16792 -9683 16848 -9681
rect 16792 -9735 16794 -9683
rect 16794 -9735 16846 -9683
rect 16846 -9735 16848 -9683
rect 16792 -9737 16848 -9735
rect 16873 -9683 16929 -9681
rect 16873 -9735 16875 -9683
rect 16875 -9735 16927 -9683
rect 16927 -9735 16929 -9683
rect 16873 -9737 16929 -9735
rect 16954 -9683 17010 -9681
rect 16954 -9735 16956 -9683
rect 16956 -9735 17008 -9683
rect 17008 -9735 17010 -9683
rect 16954 -9737 17010 -9735
rect 17035 -9683 17091 -9681
rect 17035 -9735 17037 -9683
rect 17037 -9735 17089 -9683
rect 17089 -9735 17091 -9683
rect 17035 -9737 17091 -9735
rect 17117 -9683 17173 -9681
rect 17117 -9735 17119 -9683
rect 17119 -9735 17171 -9683
rect 17171 -9735 17173 -9683
rect 17117 -9737 17173 -9735
rect 17198 -9683 17254 -9681
rect 17198 -9735 17200 -9683
rect 17200 -9735 17252 -9683
rect 17252 -9735 17254 -9683
rect 17198 -9737 17254 -9735
rect 17279 -9683 17335 -9681
rect 17279 -9735 17281 -9683
rect 17281 -9735 17333 -9683
rect 17333 -9735 17335 -9683
rect 17279 -9737 17335 -9735
rect 17360 -9683 17416 -9681
rect 17360 -9735 17362 -9683
rect 17362 -9735 17414 -9683
rect 17414 -9735 17416 -9683
rect 17360 -9737 17416 -9735
rect 17441 -9683 17497 -9681
rect 17441 -9735 17443 -9683
rect 17443 -9735 17495 -9683
rect 17495 -9735 17497 -9683
rect 17441 -9737 17497 -9735
rect 17522 -9683 17578 -9681
rect 17522 -9735 17524 -9683
rect 17524 -9735 17576 -9683
rect 17576 -9735 17578 -9683
rect 17522 -9737 17578 -9735
rect 17603 -9683 17659 -9681
rect 17603 -9735 17605 -9683
rect 17605 -9735 17657 -9683
rect 17657 -9735 17659 -9683
rect 17603 -9737 17659 -9735
rect 17684 -9683 17740 -9681
rect 17684 -9735 17686 -9683
rect 17686 -9735 17738 -9683
rect 17738 -9735 17740 -9683
rect 17684 -9737 17740 -9735
rect 17765 -9683 17821 -9681
rect 17765 -9735 17767 -9683
rect 17767 -9735 17819 -9683
rect 17819 -9735 17821 -9683
rect 17765 -9737 17821 -9735
rect 17846 -9683 17902 -9681
rect 17846 -9735 17848 -9683
rect 17848 -9735 17900 -9683
rect 17900 -9735 17902 -9683
rect 17846 -9737 17902 -9735
rect 17927 -9683 17983 -9681
rect 17927 -9735 17929 -9683
rect 17929 -9735 17981 -9683
rect 17981 -9735 17983 -9683
rect 17927 -9737 17983 -9735
rect 18008 -9683 18064 -9681
rect 18008 -9735 18010 -9683
rect 18010 -9735 18062 -9683
rect 18062 -9735 18064 -9683
rect 18008 -9737 18064 -9735
rect 18089 -9683 18145 -9681
rect 18089 -9735 18091 -9683
rect 18091 -9735 18143 -9683
rect 18143 -9735 18145 -9683
rect 18089 -9737 18145 -9735
rect 18171 -9683 18227 -9681
rect 18171 -9735 18173 -9683
rect 18173 -9735 18225 -9683
rect 18225 -9735 18227 -9683
rect 18171 -9737 18227 -9735
rect 18252 -9683 18308 -9681
rect 18252 -9735 18254 -9683
rect 18254 -9735 18306 -9683
rect 18306 -9735 18308 -9683
rect 18252 -9737 18308 -9735
rect 18333 -9683 18389 -9681
rect 18333 -9735 18335 -9683
rect 18335 -9735 18387 -9683
rect 18387 -9735 18389 -9683
rect 18333 -9737 18389 -9735
rect 18414 -9683 18470 -9681
rect 18414 -9735 18416 -9683
rect 18416 -9735 18468 -9683
rect 18468 -9735 18470 -9683
rect 18414 -9737 18470 -9735
rect 18495 -9683 18551 -9681
rect 18495 -9735 18497 -9683
rect 18497 -9735 18549 -9683
rect 18549 -9735 18551 -9683
rect 18495 -9737 18551 -9735
rect 18576 -9683 18632 -9681
rect 18576 -9735 18578 -9683
rect 18578 -9735 18630 -9683
rect 18630 -9735 18632 -9683
rect 18576 -9737 18632 -9735
rect 18657 -9683 18713 -9681
rect 18657 -9735 18659 -9683
rect 18659 -9735 18711 -9683
rect 18711 -9735 18713 -9683
rect 18657 -9737 18713 -9735
rect 18739 -9683 18795 -9681
rect 18739 -9735 18741 -9683
rect 18741 -9735 18793 -9683
rect 18793 -9735 18795 -9683
rect 18739 -9737 18795 -9735
rect 18820 -9683 18876 -9681
rect 18820 -9735 18822 -9683
rect 18822 -9735 18874 -9683
rect 18874 -9735 18876 -9683
rect 18820 -9737 18876 -9735
rect 18901 -9683 18957 -9681
rect 18901 -9735 18903 -9683
rect 18903 -9735 18955 -9683
rect 18955 -9735 18957 -9683
rect 18901 -9737 18957 -9735
rect 18982 -9683 19038 -9681
rect 18982 -9735 18984 -9683
rect 18984 -9735 19036 -9683
rect 19036 -9735 19038 -9683
rect 18982 -9737 19038 -9735
rect 19063 -9683 19119 -9681
rect 19063 -9735 19065 -9683
rect 19065 -9735 19117 -9683
rect 19117 -9735 19119 -9683
rect 19063 -9737 19119 -9735
rect 19144 -9683 19200 -9681
rect 19144 -9735 19146 -9683
rect 19146 -9735 19198 -9683
rect 19198 -9735 19200 -9683
rect 19144 -9737 19200 -9735
rect 19225 -9683 19281 -9681
rect 19225 -9735 19227 -9683
rect 19227 -9735 19279 -9683
rect 19279 -9735 19281 -9683
rect 19225 -9737 19281 -9735
rect 19307 -9683 19363 -9681
rect 19307 -9735 19309 -9683
rect 19309 -9735 19361 -9683
rect 19361 -9735 19363 -9683
rect 19307 -9737 19363 -9735
rect 19388 -9683 19444 -9681
rect 19388 -9735 19390 -9683
rect 19390 -9735 19442 -9683
rect 19442 -9735 19444 -9683
rect 19388 -9737 19444 -9735
rect 19469 -9683 19525 -9681
rect 19469 -9735 19471 -9683
rect 19471 -9735 19523 -9683
rect 19523 -9735 19525 -9683
rect 19469 -9737 19525 -9735
rect 19550 -9683 19606 -9681
rect 19550 -9735 19552 -9683
rect 19552 -9735 19604 -9683
rect 19604 -9735 19606 -9683
rect 19550 -9737 19606 -9735
rect 19631 -9683 19687 -9681
rect 19631 -9735 19633 -9683
rect 19633 -9735 19685 -9683
rect 19685 -9735 19687 -9683
rect 19631 -9737 19687 -9735
rect 19712 -9683 19768 -9681
rect 19712 -9735 19714 -9683
rect 19714 -9735 19766 -9683
rect 19766 -9735 19768 -9683
rect 19712 -9737 19768 -9735
rect 19793 -9683 19849 -9681
rect 19793 -9735 19795 -9683
rect 19795 -9735 19847 -9683
rect 19847 -9735 19849 -9683
rect 19793 -9737 19849 -9735
rect 19875 -9683 19931 -9681
rect 19875 -9735 19877 -9683
rect 19877 -9735 19929 -9683
rect 19929 -9735 19931 -9683
rect 19875 -9737 19931 -9735
rect 19956 -9683 20012 -9681
rect 19956 -9735 19958 -9683
rect 19958 -9735 20010 -9683
rect 20010 -9735 20012 -9683
rect 19956 -9737 20012 -9735
rect 20037 -9683 20093 -9681
rect 20037 -9735 20039 -9683
rect 20039 -9735 20091 -9683
rect 20091 -9735 20093 -9683
rect 20037 -9737 20093 -9735
rect 20118 -9683 20174 -9681
rect 20118 -9735 20120 -9683
rect 20120 -9735 20172 -9683
rect 20172 -9735 20174 -9683
rect 20118 -9737 20174 -9735
rect 20199 -9683 20255 -9681
rect 20199 -9735 20201 -9683
rect 20201 -9735 20253 -9683
rect 20253 -9735 20255 -9683
rect 20199 -9737 20255 -9735
rect 20280 -9683 20336 -9681
rect 20280 -9735 20282 -9683
rect 20282 -9735 20334 -9683
rect 20334 -9735 20336 -9683
rect 20280 -9737 20336 -9735
rect 20361 -9683 20417 -9681
rect 20361 -9735 20363 -9683
rect 20363 -9735 20415 -9683
rect 20415 -9735 20417 -9683
rect 20361 -9737 20417 -9735
rect 20443 -9683 20499 -9681
rect 20443 -9735 20445 -9683
rect 20445 -9735 20497 -9683
rect 20497 -9735 20499 -9683
rect 20443 -9737 20499 -9735
rect 20524 -9683 20580 -9681
rect 20524 -9735 20526 -9683
rect 20526 -9735 20578 -9683
rect 20578 -9735 20580 -9683
rect 20524 -9737 20580 -9735
rect 20605 -9683 20661 -9681
rect 20605 -9735 20607 -9683
rect 20607 -9735 20659 -9683
rect 20659 -9735 20661 -9683
rect 20605 -9737 20661 -9735
rect 20686 -9683 20742 -9681
rect 20686 -9735 20688 -9683
rect 20688 -9735 20740 -9683
rect 20740 -9735 20742 -9683
rect 20686 -9737 20742 -9735
rect 20767 -9683 20823 -9681
rect 20767 -9735 20769 -9683
rect 20769 -9735 20821 -9683
rect 20821 -9735 20823 -9683
rect 20767 -9737 20823 -9735
rect 20848 -9683 20904 -9681
rect 20848 -9735 20850 -9683
rect 20850 -9735 20902 -9683
rect 20902 -9735 20904 -9683
rect 20848 -9737 20904 -9735
rect 20929 -9683 20985 -9681
rect 20929 -9735 20931 -9683
rect 20931 -9735 20983 -9683
rect 20983 -9735 20985 -9683
rect 20929 -9737 20985 -9735
rect 21011 -9683 21067 -9681
rect 21011 -9735 21013 -9683
rect 21013 -9735 21065 -9683
rect 21065 -9735 21067 -9683
rect 21011 -9737 21067 -9735
rect 21092 -9683 21148 -9681
rect 21092 -9735 21094 -9683
rect 21094 -9735 21146 -9683
rect 21146 -9735 21148 -9683
rect 21092 -9737 21148 -9735
rect 21173 -9683 21229 -9681
rect 21173 -9735 21175 -9683
rect 21175 -9735 21227 -9683
rect 21227 -9735 21229 -9683
rect 21173 -9737 21229 -9735
rect 21254 -9683 21310 -9681
rect 21254 -9735 21256 -9683
rect 21256 -9735 21308 -9683
rect 21308 -9735 21310 -9683
rect 21254 -9737 21310 -9735
rect 21335 -9683 21391 -9681
rect 21335 -9735 21337 -9683
rect 21337 -9735 21389 -9683
rect 21389 -9735 21391 -9683
rect 21335 -9737 21391 -9735
rect 21416 -9683 21472 -9681
rect 21416 -9735 21418 -9683
rect 21418 -9735 21470 -9683
rect 21470 -9735 21472 -9683
rect 21416 -9737 21472 -9735
rect 21497 -9683 21553 -9681
rect 21497 -9735 21499 -9683
rect 21499 -9735 21551 -9683
rect 21551 -9735 21553 -9683
rect 21497 -9737 21553 -9735
rect 21579 -9683 21635 -9681
rect 21579 -9735 21581 -9683
rect 21581 -9735 21633 -9683
rect 21633 -9735 21635 -9683
rect 21579 -9737 21635 -9735
rect 21660 -9683 21716 -9681
rect 21660 -9735 21662 -9683
rect 21662 -9735 21714 -9683
rect 21714 -9735 21716 -9683
rect 21660 -9737 21716 -9735
rect 21741 -9683 21797 -9681
rect 21741 -9735 21743 -9683
rect 21743 -9735 21795 -9683
rect 21795 -9735 21797 -9683
rect 21741 -9737 21797 -9735
rect 21822 -9683 21878 -9681
rect 21822 -9735 21824 -9683
rect 21824 -9735 21876 -9683
rect 21876 -9735 21878 -9683
rect 21822 -9737 21878 -9735
rect 21903 -9683 21959 -9681
rect 21903 -9735 21905 -9683
rect 21905 -9735 21957 -9683
rect 21957 -9735 21959 -9683
rect 21903 -9737 21959 -9735
rect 21984 -9683 22040 -9681
rect 21984 -9735 21986 -9683
rect 21986 -9735 22038 -9683
rect 22038 -9735 22040 -9683
rect 21984 -9737 22040 -9735
rect 22065 -9683 22121 -9681
rect 22065 -9735 22067 -9683
rect 22067 -9735 22119 -9683
rect 22119 -9735 22121 -9683
rect 22065 -9737 22121 -9735
rect 22147 -9683 22203 -9681
rect 22147 -9735 22149 -9683
rect 22149 -9735 22201 -9683
rect 22201 -9735 22203 -9683
rect 22147 -9737 22203 -9735
rect 22228 -9683 22284 -9681
rect 22228 -9735 22230 -9683
rect 22230 -9735 22282 -9683
rect 22282 -9735 22284 -9683
rect 22228 -9737 22284 -9735
rect 22309 -9683 22365 -9681
rect 22309 -9735 22311 -9683
rect 22311 -9735 22363 -9683
rect 22363 -9735 22365 -9683
rect 22309 -9737 22365 -9735
rect 22390 -9683 22446 -9681
rect 22390 -9735 22392 -9683
rect 22392 -9735 22444 -9683
rect 22444 -9735 22446 -9683
rect 22390 -9737 22446 -9735
rect 22471 -9683 22527 -9681
rect 22471 -9735 22473 -9683
rect 22473 -9735 22525 -9683
rect 22525 -9735 22527 -9683
rect 22471 -9737 22527 -9735
rect 22552 -9683 22608 -9681
rect 22552 -9735 22554 -9683
rect 22554 -9735 22606 -9683
rect 22606 -9735 22608 -9683
rect 22552 -9737 22608 -9735
rect 22633 -9683 22689 -9681
rect 22633 -9735 22635 -9683
rect 22635 -9735 22687 -9683
rect 22687 -9735 22689 -9683
rect 22633 -9737 22689 -9735
rect 22715 -9683 22771 -9681
rect 22715 -9735 22717 -9683
rect 22717 -9735 22769 -9683
rect 22769 -9735 22771 -9683
rect 22715 -9737 22771 -9735
rect 22796 -9683 22852 -9681
rect 22796 -9735 22798 -9683
rect 22798 -9735 22850 -9683
rect 22850 -9735 22852 -9683
rect 22796 -9737 22852 -9735
rect 22877 -9683 22933 -9681
rect 22877 -9735 22879 -9683
rect 22879 -9735 22931 -9683
rect 22931 -9735 22933 -9683
rect 22877 -9737 22933 -9735
rect 22958 -9683 23014 -9681
rect 22958 -9735 22960 -9683
rect 22960 -9735 23012 -9683
rect 23012 -9735 23014 -9683
rect 22958 -9737 23014 -9735
rect 23039 -9683 23095 -9681
rect 23039 -9735 23041 -9683
rect 23041 -9735 23093 -9683
rect 23093 -9735 23095 -9683
rect 23039 -9737 23095 -9735
rect 23120 -9683 23176 -9681
rect 23120 -9735 23122 -9683
rect 23122 -9735 23174 -9683
rect 23174 -9735 23176 -9683
rect 23120 -9737 23176 -9735
rect 23201 -9683 23257 -9681
rect 23201 -9735 23203 -9683
rect 23203 -9735 23255 -9683
rect 23255 -9735 23257 -9683
rect 23201 -9737 23257 -9735
rect 23283 -9683 23339 -9681
rect 23283 -9735 23285 -9683
rect 23285 -9735 23337 -9683
rect 23337 -9735 23339 -9683
rect 23283 -9737 23339 -9735
rect 23364 -9683 23420 -9681
rect 23364 -9735 23366 -9683
rect 23366 -9735 23418 -9683
rect 23418 -9735 23420 -9683
rect 23364 -9737 23420 -9735
rect 23445 -9683 23501 -9681
rect 23445 -9735 23447 -9683
rect 23447 -9735 23499 -9683
rect 23499 -9735 23501 -9683
rect 23445 -9737 23501 -9735
rect 23526 -9683 23582 -9681
rect 23526 -9735 23528 -9683
rect 23528 -9735 23580 -9683
rect 23580 -9735 23582 -9683
rect 23526 -9737 23582 -9735
rect 23607 -9683 23663 -9681
rect 23607 -9735 23609 -9683
rect 23609 -9735 23661 -9683
rect 23661 -9735 23663 -9683
rect 23607 -9737 23663 -9735
rect 23688 -9683 23744 -9681
rect 23688 -9735 23690 -9683
rect 23690 -9735 23742 -9683
rect 23742 -9735 23744 -9683
rect 23688 -9737 23744 -9735
rect 23769 -9683 23825 -9681
rect 23769 -9735 23771 -9683
rect 23771 -9735 23823 -9683
rect 23823 -9735 23825 -9683
rect 23769 -9737 23825 -9735
rect 23851 -9683 23907 -9681
rect 23851 -9735 23853 -9683
rect 23853 -9735 23905 -9683
rect 23905 -9735 23907 -9683
rect 23851 -9737 23907 -9735
rect 23932 -9683 23988 -9681
rect 23932 -9735 23934 -9683
rect 23934 -9735 23986 -9683
rect 23986 -9735 23988 -9683
rect 23932 -9737 23988 -9735
rect 24013 -9683 24069 -9681
rect 24013 -9735 24015 -9683
rect 24015 -9735 24067 -9683
rect 24067 -9735 24069 -9683
rect 24013 -9737 24069 -9735
rect 24094 -9683 24150 -9681
rect 24094 -9735 24096 -9683
rect 24096 -9735 24148 -9683
rect 24148 -9735 24150 -9683
rect 24094 -9737 24150 -9735
rect 24175 -9683 24231 -9681
rect 24175 -9735 24177 -9683
rect 24177 -9735 24229 -9683
rect 24229 -9735 24231 -9683
rect 24175 -9737 24231 -9735
rect 24256 -9683 24312 -9681
rect 24256 -9735 24258 -9683
rect 24258 -9735 24310 -9683
rect 24310 -9735 24312 -9683
rect 24256 -9737 24312 -9735
rect 24337 -9683 24393 -9681
rect 24337 -9735 24339 -9683
rect 24339 -9735 24391 -9683
rect 24391 -9735 24393 -9683
rect 24337 -9737 24393 -9735
rect 24419 -9683 24475 -9681
rect 24419 -9735 24421 -9683
rect 24421 -9735 24473 -9683
rect 24473 -9735 24475 -9683
rect 24419 -9737 24475 -9735
rect 24500 -9683 24556 -9681
rect 24500 -9735 24502 -9683
rect 24502 -9735 24554 -9683
rect 24554 -9735 24556 -9683
rect 24500 -9737 24556 -9735
rect 24581 -9683 24637 -9681
rect 24581 -9735 24583 -9683
rect 24583 -9735 24635 -9683
rect 24635 -9735 24637 -9683
rect 24581 -9737 24637 -9735
rect 24662 -9683 24718 -9681
rect 24662 -9735 24664 -9683
rect 24664 -9735 24716 -9683
rect 24716 -9735 24718 -9683
rect 24662 -9737 24718 -9735
rect 24743 -9683 24799 -9681
rect 24743 -9735 24745 -9683
rect 24745 -9735 24797 -9683
rect 24797 -9735 24799 -9683
rect 24743 -9737 24799 -9735
rect 24824 -9683 24880 -9681
rect 24824 -9735 24826 -9683
rect 24826 -9735 24878 -9683
rect 24878 -9735 24880 -9683
rect 24824 -9737 24880 -9735
rect 24905 -9683 24961 -9681
rect 24905 -9735 24907 -9683
rect 24907 -9735 24959 -9683
rect 24959 -9735 24961 -9683
rect 24905 -9737 24961 -9735
rect 24987 -9683 25043 -9681
rect 24987 -9735 24989 -9683
rect 24989 -9735 25041 -9683
rect 25041 -9735 25043 -9683
rect 24987 -9737 25043 -9735
rect 25068 -9683 25124 -9681
rect 25068 -9735 25070 -9683
rect 25070 -9735 25122 -9683
rect 25122 -9735 25124 -9683
rect 25068 -9737 25124 -9735
rect 25149 -9683 25205 -9681
rect 25149 -9735 25151 -9683
rect 25151 -9735 25203 -9683
rect 25203 -9735 25205 -9683
rect 25149 -9737 25205 -9735
rect 25230 -9683 25286 -9681
rect 25230 -9735 25232 -9683
rect 25232 -9735 25284 -9683
rect 25284 -9735 25286 -9683
rect 25230 -9737 25286 -9735
rect 25311 -9683 25367 -9681
rect 25311 -9735 25313 -9683
rect 25313 -9735 25365 -9683
rect 25365 -9735 25367 -9683
rect 25311 -9737 25367 -9735
rect 25392 -9683 25448 -9681
rect 25392 -9735 25394 -9683
rect 25394 -9735 25446 -9683
rect 25446 -9735 25448 -9683
rect 25392 -9737 25448 -9735
rect 25473 -9683 25529 -9681
rect 25473 -9735 25475 -9683
rect 25475 -9735 25527 -9683
rect 25527 -9735 25529 -9683
rect 25473 -9737 25529 -9735
rect 25555 -9683 25611 -9681
rect 25555 -9735 25557 -9683
rect 25557 -9735 25609 -9683
rect 25609 -9735 25611 -9683
rect 25555 -9737 25611 -9735
rect 25636 -9683 25692 -9681
rect 25636 -9735 25638 -9683
rect 25638 -9735 25690 -9683
rect 25690 -9735 25692 -9683
rect 25636 -9737 25692 -9735
rect 25717 -9683 25773 -9681
rect 25717 -9735 25719 -9683
rect 25719 -9735 25771 -9683
rect 25771 -9735 25773 -9683
rect 25717 -9737 25773 -9735
rect 25798 -9683 25854 -9681
rect 25798 -9735 25800 -9683
rect 25800 -9735 25852 -9683
rect 25852 -9735 25854 -9683
rect 25798 -9737 25854 -9735
rect 25879 -9683 25935 -9681
rect 25879 -9735 25881 -9683
rect 25881 -9735 25933 -9683
rect 25933 -9735 25935 -9683
rect 25879 -9737 25935 -9735
rect 25960 -9683 26016 -9681
rect 25960 -9735 25962 -9683
rect 25962 -9735 26014 -9683
rect 26014 -9735 26016 -9683
rect 25960 -9737 26016 -9735
rect 26041 -9683 26097 -9681
rect 26041 -9735 26043 -9683
rect 26043 -9735 26095 -9683
rect 26095 -9735 26097 -9683
rect 26041 -9737 26097 -9735
rect 26123 -9683 26179 -9681
rect 26123 -9735 26125 -9683
rect 26125 -9735 26177 -9683
rect 26177 -9735 26179 -9683
rect 26123 -9737 26179 -9735
rect 26204 -9683 26260 -9681
rect 26204 -9735 26206 -9683
rect 26206 -9735 26258 -9683
rect 26258 -9735 26260 -9683
rect 26204 -9737 26260 -9735
rect 4053 -9787 4109 -9785
rect 4053 -9839 4055 -9787
rect 4055 -9839 4107 -9787
rect 4107 -9839 4109 -9787
rect 4053 -9841 4109 -9839
rect 4134 -9787 4190 -9785
rect 4134 -9839 4136 -9787
rect 4136 -9839 4188 -9787
rect 4188 -9839 4190 -9787
rect 4134 -9841 4190 -9839
rect 4215 -9787 4271 -9785
rect 4215 -9839 4217 -9787
rect 4217 -9839 4269 -9787
rect 4269 -9839 4271 -9787
rect 4215 -9841 4271 -9839
rect 4296 -9787 4352 -9785
rect 4296 -9839 4298 -9787
rect 4298 -9839 4350 -9787
rect 4350 -9839 4352 -9787
rect 4296 -9841 4352 -9839
rect 4377 -9787 4433 -9785
rect 4377 -9839 4379 -9787
rect 4379 -9839 4431 -9787
rect 4431 -9839 4433 -9787
rect 4377 -9841 4433 -9839
rect 4458 -9787 4514 -9785
rect 4458 -9839 4460 -9787
rect 4460 -9839 4512 -9787
rect 4512 -9839 4514 -9787
rect 4458 -9841 4514 -9839
rect 4539 -9787 4595 -9785
rect 4539 -9839 4541 -9787
rect 4541 -9839 4593 -9787
rect 4593 -9839 4595 -9787
rect 4539 -9841 4595 -9839
rect 4621 -9787 4677 -9785
rect 4621 -9839 4623 -9787
rect 4623 -9839 4675 -9787
rect 4675 -9839 4677 -9787
rect 4621 -9841 4677 -9839
rect 4702 -9787 4758 -9785
rect 4702 -9839 4704 -9787
rect 4704 -9839 4756 -9787
rect 4756 -9839 4758 -9787
rect 4702 -9841 4758 -9839
rect 4783 -9787 4839 -9785
rect 4783 -9839 4785 -9787
rect 4785 -9839 4837 -9787
rect 4837 -9839 4839 -9787
rect 4783 -9841 4839 -9839
rect 4864 -9787 4920 -9785
rect 4864 -9839 4866 -9787
rect 4866 -9839 4918 -9787
rect 4918 -9839 4920 -9787
rect 4864 -9841 4920 -9839
rect 4945 -9787 5001 -9785
rect 4945 -9839 4947 -9787
rect 4947 -9839 4999 -9787
rect 4999 -9839 5001 -9787
rect 4945 -9841 5001 -9839
rect 5026 -9787 5082 -9785
rect 5026 -9839 5028 -9787
rect 5028 -9839 5080 -9787
rect 5080 -9839 5082 -9787
rect 5026 -9841 5082 -9839
rect 5107 -9787 5163 -9785
rect 5107 -9839 5109 -9787
rect 5109 -9839 5161 -9787
rect 5161 -9839 5163 -9787
rect 5107 -9841 5163 -9839
rect 5189 -9787 5245 -9785
rect 5189 -9839 5191 -9787
rect 5191 -9839 5243 -9787
rect 5243 -9839 5245 -9787
rect 5189 -9841 5245 -9839
rect 5270 -9787 5326 -9785
rect 5270 -9839 5272 -9787
rect 5272 -9839 5324 -9787
rect 5324 -9839 5326 -9787
rect 5270 -9841 5326 -9839
rect 5351 -9787 5407 -9785
rect 5351 -9839 5353 -9787
rect 5353 -9839 5405 -9787
rect 5405 -9839 5407 -9787
rect 5351 -9841 5407 -9839
rect 5432 -9787 5488 -9785
rect 5432 -9839 5434 -9787
rect 5434 -9839 5486 -9787
rect 5486 -9839 5488 -9787
rect 5432 -9841 5488 -9839
rect 5513 -9787 5569 -9785
rect 5513 -9839 5515 -9787
rect 5515 -9839 5567 -9787
rect 5567 -9839 5569 -9787
rect 5513 -9841 5569 -9839
rect 5594 -9787 5650 -9785
rect 5594 -9839 5596 -9787
rect 5596 -9839 5648 -9787
rect 5648 -9839 5650 -9787
rect 5594 -9841 5650 -9839
rect 5675 -9787 5731 -9785
rect 5675 -9839 5677 -9787
rect 5677 -9839 5729 -9787
rect 5729 -9839 5731 -9787
rect 5675 -9841 5731 -9839
rect 5757 -9787 5813 -9785
rect 5757 -9839 5759 -9787
rect 5759 -9839 5811 -9787
rect 5811 -9839 5813 -9787
rect 5757 -9841 5813 -9839
rect 5838 -9787 5894 -9785
rect 5838 -9839 5840 -9787
rect 5840 -9839 5892 -9787
rect 5892 -9839 5894 -9787
rect 5838 -9841 5894 -9839
rect 5919 -9787 5975 -9785
rect 5919 -9839 5921 -9787
rect 5921 -9839 5973 -9787
rect 5973 -9839 5975 -9787
rect 5919 -9841 5975 -9839
rect 6000 -9787 6056 -9785
rect 6000 -9839 6002 -9787
rect 6002 -9839 6054 -9787
rect 6054 -9839 6056 -9787
rect 6000 -9841 6056 -9839
rect 6081 -9787 6137 -9785
rect 6081 -9839 6083 -9787
rect 6083 -9839 6135 -9787
rect 6135 -9839 6137 -9787
rect 6081 -9841 6137 -9839
rect 6162 -9787 6218 -9785
rect 6162 -9839 6164 -9787
rect 6164 -9839 6216 -9787
rect 6216 -9839 6218 -9787
rect 6162 -9841 6218 -9839
rect 6243 -9787 6299 -9785
rect 6243 -9839 6245 -9787
rect 6245 -9839 6297 -9787
rect 6297 -9839 6299 -9787
rect 6243 -9841 6299 -9839
rect 6325 -9787 6381 -9785
rect 6325 -9839 6327 -9787
rect 6327 -9839 6379 -9787
rect 6379 -9839 6381 -9787
rect 6325 -9841 6381 -9839
rect 6406 -9787 6462 -9785
rect 6406 -9839 6408 -9787
rect 6408 -9839 6460 -9787
rect 6460 -9839 6462 -9787
rect 6406 -9841 6462 -9839
rect 6487 -9787 6543 -9785
rect 6487 -9839 6489 -9787
rect 6489 -9839 6541 -9787
rect 6541 -9839 6543 -9787
rect 6487 -9841 6543 -9839
rect 6568 -9787 6624 -9785
rect 6568 -9839 6570 -9787
rect 6570 -9839 6622 -9787
rect 6622 -9839 6624 -9787
rect 6568 -9841 6624 -9839
rect 6649 -9787 6705 -9785
rect 6649 -9839 6651 -9787
rect 6651 -9839 6703 -9787
rect 6703 -9839 6705 -9787
rect 6649 -9841 6705 -9839
rect 6730 -9787 6786 -9785
rect 6730 -9839 6732 -9787
rect 6732 -9839 6784 -9787
rect 6784 -9839 6786 -9787
rect 6730 -9841 6786 -9839
rect 6811 -9787 6867 -9785
rect 6811 -9839 6813 -9787
rect 6813 -9839 6865 -9787
rect 6865 -9839 6867 -9787
rect 6811 -9841 6867 -9839
rect 6893 -9787 6949 -9785
rect 6893 -9839 6895 -9787
rect 6895 -9839 6947 -9787
rect 6947 -9839 6949 -9787
rect 6893 -9841 6949 -9839
rect 6974 -9787 7030 -9785
rect 6974 -9839 6976 -9787
rect 6976 -9839 7028 -9787
rect 7028 -9839 7030 -9787
rect 6974 -9841 7030 -9839
rect 7055 -9787 7111 -9785
rect 7055 -9839 7057 -9787
rect 7057 -9839 7109 -9787
rect 7109 -9839 7111 -9787
rect 7055 -9841 7111 -9839
rect 7136 -9787 7192 -9785
rect 7136 -9839 7138 -9787
rect 7138 -9839 7190 -9787
rect 7190 -9839 7192 -9787
rect 7136 -9841 7192 -9839
rect 7217 -9787 7273 -9785
rect 7217 -9839 7219 -9787
rect 7219 -9839 7271 -9787
rect 7271 -9839 7273 -9787
rect 7217 -9841 7273 -9839
rect 7298 -9787 7354 -9785
rect 7298 -9839 7300 -9787
rect 7300 -9839 7352 -9787
rect 7352 -9839 7354 -9787
rect 7298 -9841 7354 -9839
rect 7379 -9787 7435 -9785
rect 7379 -9839 7381 -9787
rect 7381 -9839 7433 -9787
rect 7433 -9839 7435 -9787
rect 7379 -9841 7435 -9839
rect 7461 -9787 7517 -9785
rect 7461 -9839 7463 -9787
rect 7463 -9839 7515 -9787
rect 7515 -9839 7517 -9787
rect 7461 -9841 7517 -9839
rect 7542 -9787 7598 -9785
rect 7542 -9839 7544 -9787
rect 7544 -9839 7596 -9787
rect 7596 -9839 7598 -9787
rect 7542 -9841 7598 -9839
rect 7623 -9787 7679 -9785
rect 7623 -9839 7625 -9787
rect 7625 -9839 7677 -9787
rect 7677 -9839 7679 -9787
rect 7623 -9841 7679 -9839
rect 7704 -9787 7760 -9785
rect 7704 -9839 7706 -9787
rect 7706 -9839 7758 -9787
rect 7758 -9839 7760 -9787
rect 7704 -9841 7760 -9839
rect 7785 -9787 7841 -9785
rect 7785 -9839 7787 -9787
rect 7787 -9839 7839 -9787
rect 7839 -9839 7841 -9787
rect 7785 -9841 7841 -9839
rect 7866 -9787 7922 -9785
rect 7866 -9839 7868 -9787
rect 7868 -9839 7920 -9787
rect 7920 -9839 7922 -9787
rect 7866 -9841 7922 -9839
rect 7947 -9787 8003 -9785
rect 7947 -9839 7949 -9787
rect 7949 -9839 8001 -9787
rect 8001 -9839 8003 -9787
rect 7947 -9841 8003 -9839
rect 8029 -9787 8085 -9785
rect 8029 -9839 8031 -9787
rect 8031 -9839 8083 -9787
rect 8083 -9839 8085 -9787
rect 8029 -9841 8085 -9839
rect 8110 -9787 8166 -9785
rect 8110 -9839 8112 -9787
rect 8112 -9839 8164 -9787
rect 8164 -9839 8166 -9787
rect 8110 -9841 8166 -9839
rect 8191 -9787 8247 -9785
rect 8191 -9839 8193 -9787
rect 8193 -9839 8245 -9787
rect 8245 -9839 8247 -9787
rect 8191 -9841 8247 -9839
rect 8272 -9787 8328 -9785
rect 8272 -9839 8274 -9787
rect 8274 -9839 8326 -9787
rect 8326 -9839 8328 -9787
rect 8272 -9841 8328 -9839
rect 8353 -9787 8409 -9785
rect 8353 -9839 8355 -9787
rect 8355 -9839 8407 -9787
rect 8407 -9839 8409 -9787
rect 8353 -9841 8409 -9839
rect 8434 -9787 8490 -9785
rect 8434 -9839 8436 -9787
rect 8436 -9839 8488 -9787
rect 8488 -9839 8490 -9787
rect 8434 -9841 8490 -9839
rect 8515 -9787 8571 -9785
rect 8515 -9839 8517 -9787
rect 8517 -9839 8569 -9787
rect 8569 -9839 8571 -9787
rect 8515 -9841 8571 -9839
rect 8597 -9787 8653 -9785
rect 8597 -9839 8599 -9787
rect 8599 -9839 8651 -9787
rect 8651 -9839 8653 -9787
rect 8597 -9841 8653 -9839
rect 8678 -9787 8734 -9785
rect 8678 -9839 8680 -9787
rect 8680 -9839 8732 -9787
rect 8732 -9839 8734 -9787
rect 8678 -9841 8734 -9839
rect 8759 -9787 8815 -9785
rect 8759 -9839 8761 -9787
rect 8761 -9839 8813 -9787
rect 8813 -9839 8815 -9787
rect 8759 -9841 8815 -9839
rect 8840 -9787 8896 -9785
rect 8840 -9839 8842 -9787
rect 8842 -9839 8894 -9787
rect 8894 -9839 8896 -9787
rect 8840 -9841 8896 -9839
rect 8921 -9787 8977 -9785
rect 8921 -9839 8923 -9787
rect 8923 -9839 8975 -9787
rect 8975 -9839 8977 -9787
rect 8921 -9841 8977 -9839
rect 9002 -9787 9058 -9785
rect 9002 -9839 9004 -9787
rect 9004 -9839 9056 -9787
rect 9056 -9839 9058 -9787
rect 9002 -9841 9058 -9839
rect 9083 -9787 9139 -9785
rect 9083 -9839 9085 -9787
rect 9085 -9839 9137 -9787
rect 9137 -9839 9139 -9787
rect 9083 -9841 9139 -9839
rect 9165 -9787 9221 -9785
rect 9165 -9839 9167 -9787
rect 9167 -9839 9219 -9787
rect 9219 -9839 9221 -9787
rect 9165 -9841 9221 -9839
rect 9246 -9787 9302 -9785
rect 9246 -9839 9248 -9787
rect 9248 -9839 9300 -9787
rect 9300 -9839 9302 -9787
rect 9246 -9841 9302 -9839
rect 9327 -9787 9383 -9785
rect 9327 -9839 9329 -9787
rect 9329 -9839 9381 -9787
rect 9381 -9839 9383 -9787
rect 9327 -9841 9383 -9839
rect 9408 -9787 9464 -9785
rect 9408 -9839 9410 -9787
rect 9410 -9839 9462 -9787
rect 9462 -9839 9464 -9787
rect 9408 -9841 9464 -9839
rect 9489 -9787 9545 -9785
rect 9489 -9839 9491 -9787
rect 9491 -9839 9543 -9787
rect 9543 -9839 9545 -9787
rect 9489 -9841 9545 -9839
rect 9570 -9787 9626 -9785
rect 9570 -9839 9572 -9787
rect 9572 -9839 9624 -9787
rect 9624 -9839 9626 -9787
rect 9570 -9841 9626 -9839
rect 9651 -9787 9707 -9785
rect 9651 -9839 9653 -9787
rect 9653 -9839 9705 -9787
rect 9705 -9839 9707 -9787
rect 9651 -9841 9707 -9839
rect 9733 -9787 9789 -9785
rect 9733 -9839 9735 -9787
rect 9735 -9839 9787 -9787
rect 9787 -9839 9789 -9787
rect 9733 -9841 9789 -9839
rect 9814 -9787 9870 -9785
rect 9814 -9839 9816 -9787
rect 9816 -9839 9868 -9787
rect 9868 -9839 9870 -9787
rect 9814 -9841 9870 -9839
rect 9895 -9787 9951 -9785
rect 9895 -9839 9897 -9787
rect 9897 -9839 9949 -9787
rect 9949 -9839 9951 -9787
rect 9895 -9841 9951 -9839
rect 9976 -9787 10032 -9785
rect 9976 -9839 9978 -9787
rect 9978 -9839 10030 -9787
rect 10030 -9839 10032 -9787
rect 9976 -9841 10032 -9839
rect 10057 -9787 10113 -9785
rect 10057 -9839 10059 -9787
rect 10059 -9839 10111 -9787
rect 10111 -9839 10113 -9787
rect 10057 -9841 10113 -9839
rect 10138 -9787 10194 -9785
rect 10138 -9839 10140 -9787
rect 10140 -9839 10192 -9787
rect 10192 -9839 10194 -9787
rect 10138 -9841 10194 -9839
rect 10219 -9787 10275 -9785
rect 10219 -9839 10221 -9787
rect 10221 -9839 10273 -9787
rect 10273 -9839 10275 -9787
rect 10219 -9841 10275 -9839
rect 10301 -9787 10357 -9785
rect 10301 -9839 10303 -9787
rect 10303 -9839 10355 -9787
rect 10355 -9839 10357 -9787
rect 10301 -9841 10357 -9839
rect 10382 -9787 10438 -9785
rect 10382 -9839 10384 -9787
rect 10384 -9839 10436 -9787
rect 10436 -9839 10438 -9787
rect 10382 -9841 10438 -9839
rect 10463 -9787 10519 -9785
rect 10463 -9839 10465 -9787
rect 10465 -9839 10517 -9787
rect 10517 -9839 10519 -9787
rect 10463 -9841 10519 -9839
rect 10544 -9787 10600 -9785
rect 10544 -9839 10546 -9787
rect 10546 -9839 10598 -9787
rect 10598 -9839 10600 -9787
rect 10544 -9841 10600 -9839
rect 10625 -9787 10681 -9785
rect 10625 -9839 10627 -9787
rect 10627 -9839 10679 -9787
rect 10679 -9839 10681 -9787
rect 10625 -9841 10681 -9839
rect 10706 -9787 10762 -9785
rect 10706 -9839 10708 -9787
rect 10708 -9839 10760 -9787
rect 10760 -9839 10762 -9787
rect 10706 -9841 10762 -9839
rect 10787 -9787 10843 -9785
rect 10787 -9839 10789 -9787
rect 10789 -9839 10841 -9787
rect 10841 -9839 10843 -9787
rect 10787 -9841 10843 -9839
rect 10869 -9787 10925 -9785
rect 10869 -9839 10871 -9787
rect 10871 -9839 10923 -9787
rect 10923 -9839 10925 -9787
rect 10869 -9841 10925 -9839
rect 10950 -9787 11006 -9785
rect 10950 -9839 10952 -9787
rect 10952 -9839 11004 -9787
rect 11004 -9839 11006 -9787
rect 10950 -9841 11006 -9839
rect 11031 -9787 11087 -9785
rect 11031 -9839 11033 -9787
rect 11033 -9839 11085 -9787
rect 11085 -9839 11087 -9787
rect 11031 -9841 11087 -9839
rect 11112 -9787 11168 -9785
rect 11112 -9839 11114 -9787
rect 11114 -9839 11166 -9787
rect 11166 -9839 11168 -9787
rect 11112 -9841 11168 -9839
rect 11193 -9787 11249 -9785
rect 11193 -9839 11195 -9787
rect 11195 -9839 11247 -9787
rect 11247 -9839 11249 -9787
rect 11193 -9841 11249 -9839
rect 11274 -9787 11330 -9785
rect 11274 -9839 11276 -9787
rect 11276 -9839 11328 -9787
rect 11328 -9839 11330 -9787
rect 11274 -9841 11330 -9839
rect 11355 -9787 11411 -9785
rect 11355 -9839 11357 -9787
rect 11357 -9839 11409 -9787
rect 11409 -9839 11411 -9787
rect 11355 -9841 11411 -9839
rect 11437 -9787 11493 -9785
rect 11437 -9839 11439 -9787
rect 11439 -9839 11491 -9787
rect 11491 -9839 11493 -9787
rect 11437 -9841 11493 -9839
rect 11518 -9787 11574 -9785
rect 11518 -9839 11520 -9787
rect 11520 -9839 11572 -9787
rect 11572 -9839 11574 -9787
rect 11518 -9841 11574 -9839
rect 11599 -9787 11655 -9785
rect 11599 -9839 11601 -9787
rect 11601 -9839 11653 -9787
rect 11653 -9839 11655 -9787
rect 11599 -9841 11655 -9839
rect 11680 -9787 11736 -9785
rect 11680 -9839 11682 -9787
rect 11682 -9839 11734 -9787
rect 11734 -9839 11736 -9787
rect 11680 -9841 11736 -9839
rect 11761 -9787 11817 -9785
rect 11761 -9839 11763 -9787
rect 11763 -9839 11815 -9787
rect 11815 -9839 11817 -9787
rect 11761 -9841 11817 -9839
rect 11842 -9787 11898 -9785
rect 11842 -9839 11844 -9787
rect 11844 -9839 11896 -9787
rect 11896 -9839 11898 -9787
rect 11842 -9841 11898 -9839
rect 11923 -9787 11979 -9785
rect 11923 -9839 11925 -9787
rect 11925 -9839 11977 -9787
rect 11977 -9839 11979 -9787
rect 11923 -9841 11979 -9839
rect 12005 -9787 12061 -9785
rect 12005 -9839 12007 -9787
rect 12007 -9839 12059 -9787
rect 12059 -9839 12061 -9787
rect 12005 -9841 12061 -9839
rect 12086 -9787 12142 -9785
rect 12086 -9839 12088 -9787
rect 12088 -9839 12140 -9787
rect 12140 -9839 12142 -9787
rect 12086 -9841 12142 -9839
rect 12167 -9787 12223 -9785
rect 12167 -9839 12169 -9787
rect 12169 -9839 12221 -9787
rect 12221 -9839 12223 -9787
rect 12167 -9841 12223 -9839
rect 12248 -9787 12304 -9785
rect 12248 -9839 12250 -9787
rect 12250 -9839 12302 -9787
rect 12302 -9839 12304 -9787
rect 12248 -9841 12304 -9839
rect 12329 -9787 12385 -9785
rect 12329 -9839 12331 -9787
rect 12331 -9839 12383 -9787
rect 12383 -9839 12385 -9787
rect 12329 -9841 12385 -9839
rect 12410 -9787 12466 -9785
rect 12410 -9839 12412 -9787
rect 12412 -9839 12464 -9787
rect 12464 -9839 12466 -9787
rect 12410 -9841 12466 -9839
rect 12491 -9787 12547 -9785
rect 12491 -9839 12493 -9787
rect 12493 -9839 12545 -9787
rect 12545 -9839 12547 -9787
rect 12491 -9841 12547 -9839
rect 12573 -9787 12629 -9785
rect 12573 -9839 12575 -9787
rect 12575 -9839 12627 -9787
rect 12627 -9839 12629 -9787
rect 12573 -9841 12629 -9839
rect 12654 -9787 12710 -9785
rect 12654 -9839 12656 -9787
rect 12656 -9839 12708 -9787
rect 12708 -9839 12710 -9787
rect 12654 -9841 12710 -9839
rect 12735 -9787 12791 -9785
rect 12735 -9839 12737 -9787
rect 12737 -9839 12789 -9787
rect 12789 -9839 12791 -9787
rect 12735 -9841 12791 -9839
rect 12816 -9787 12872 -9785
rect 12816 -9839 12818 -9787
rect 12818 -9839 12870 -9787
rect 12870 -9839 12872 -9787
rect 12816 -9841 12872 -9839
rect 12897 -9787 12953 -9785
rect 12897 -9839 12899 -9787
rect 12899 -9839 12951 -9787
rect 12951 -9839 12953 -9787
rect 12897 -9841 12953 -9839
rect 12978 -9787 13034 -9785
rect 12978 -9839 12980 -9787
rect 12980 -9839 13032 -9787
rect 13032 -9839 13034 -9787
rect 12978 -9841 13034 -9839
rect 13059 -9787 13115 -9785
rect 13059 -9839 13061 -9787
rect 13061 -9839 13113 -9787
rect 13113 -9839 13115 -9787
rect 13059 -9841 13115 -9839
rect 13141 -9787 13197 -9785
rect 13141 -9839 13143 -9787
rect 13143 -9839 13195 -9787
rect 13195 -9839 13197 -9787
rect 13141 -9841 13197 -9839
rect 13222 -9787 13278 -9785
rect 13222 -9839 13224 -9787
rect 13224 -9839 13276 -9787
rect 13276 -9839 13278 -9787
rect 13222 -9841 13278 -9839
rect 13303 -9787 13359 -9785
rect 13303 -9839 13305 -9787
rect 13305 -9839 13357 -9787
rect 13357 -9839 13359 -9787
rect 13303 -9841 13359 -9839
rect 13384 -9787 13440 -9785
rect 13384 -9839 13386 -9787
rect 13386 -9839 13438 -9787
rect 13438 -9839 13440 -9787
rect 13384 -9841 13440 -9839
rect 13465 -9787 13521 -9785
rect 13465 -9839 13467 -9787
rect 13467 -9839 13519 -9787
rect 13519 -9839 13521 -9787
rect 13465 -9841 13521 -9839
rect 13546 -9787 13602 -9785
rect 13546 -9839 13548 -9787
rect 13548 -9839 13600 -9787
rect 13600 -9839 13602 -9787
rect 13546 -9841 13602 -9839
rect 13627 -9787 13683 -9785
rect 13627 -9839 13629 -9787
rect 13629 -9839 13681 -9787
rect 13681 -9839 13683 -9787
rect 13627 -9841 13683 -9839
rect 13709 -9787 13765 -9785
rect 13709 -9839 13711 -9787
rect 13711 -9839 13763 -9787
rect 13763 -9839 13765 -9787
rect 13709 -9841 13765 -9839
rect 13790 -9787 13846 -9785
rect 13790 -9839 13792 -9787
rect 13792 -9839 13844 -9787
rect 13844 -9839 13846 -9787
rect 13790 -9841 13846 -9839
rect 13871 -9787 13927 -9785
rect 13871 -9839 13873 -9787
rect 13873 -9839 13925 -9787
rect 13925 -9839 13927 -9787
rect 13871 -9841 13927 -9839
rect 13952 -9787 14008 -9785
rect 13952 -9839 13954 -9787
rect 13954 -9839 14006 -9787
rect 14006 -9839 14008 -9787
rect 13952 -9841 14008 -9839
rect 14033 -9787 14089 -9785
rect 14033 -9839 14035 -9787
rect 14035 -9839 14087 -9787
rect 14087 -9839 14089 -9787
rect 14033 -9841 14089 -9839
rect 14114 -9787 14170 -9785
rect 14114 -9839 14116 -9787
rect 14116 -9839 14168 -9787
rect 14168 -9839 14170 -9787
rect 14114 -9841 14170 -9839
rect 14195 -9787 14251 -9785
rect 14195 -9839 14197 -9787
rect 14197 -9839 14249 -9787
rect 14249 -9839 14251 -9787
rect 14195 -9841 14251 -9839
rect 14277 -9787 14333 -9785
rect 14277 -9839 14279 -9787
rect 14279 -9839 14331 -9787
rect 14331 -9839 14333 -9787
rect 14277 -9841 14333 -9839
rect 14358 -9787 14414 -9785
rect 14358 -9839 14360 -9787
rect 14360 -9839 14412 -9787
rect 14412 -9839 14414 -9787
rect 14358 -9841 14414 -9839
rect 14439 -9787 14495 -9785
rect 14439 -9839 14441 -9787
rect 14441 -9839 14493 -9787
rect 14493 -9839 14495 -9787
rect 14439 -9841 14495 -9839
rect 14520 -9787 14576 -9785
rect 14520 -9839 14522 -9787
rect 14522 -9839 14574 -9787
rect 14574 -9839 14576 -9787
rect 14520 -9841 14576 -9839
rect 14601 -9787 14657 -9785
rect 14601 -9839 14603 -9787
rect 14603 -9839 14655 -9787
rect 14655 -9839 14657 -9787
rect 14601 -9841 14657 -9839
rect 14682 -9787 14738 -9785
rect 14682 -9839 14684 -9787
rect 14684 -9839 14736 -9787
rect 14736 -9839 14738 -9787
rect 14682 -9841 14738 -9839
rect 14763 -9787 14819 -9785
rect 14763 -9839 14765 -9787
rect 14765 -9839 14817 -9787
rect 14817 -9839 14819 -9787
rect 14763 -9841 14819 -9839
rect 14845 -9787 14901 -9785
rect 14845 -9839 14847 -9787
rect 14847 -9839 14899 -9787
rect 14899 -9839 14901 -9787
rect 14845 -9841 14901 -9839
rect 14926 -9787 14982 -9785
rect 14926 -9839 14928 -9787
rect 14928 -9839 14980 -9787
rect 14980 -9839 14982 -9787
rect 14926 -9841 14982 -9839
rect 15007 -9787 15063 -9785
rect 15007 -9839 15009 -9787
rect 15009 -9839 15061 -9787
rect 15061 -9839 15063 -9787
rect 15007 -9841 15063 -9839
rect 15088 -9787 15144 -9785
rect 15088 -9839 15090 -9787
rect 15090 -9839 15142 -9787
rect 15142 -9839 15144 -9787
rect 15088 -9841 15144 -9839
rect 15169 -9787 15225 -9785
rect 15169 -9839 15171 -9787
rect 15171 -9839 15223 -9787
rect 15223 -9839 15225 -9787
rect 15169 -9841 15225 -9839
rect 15250 -9787 15306 -9785
rect 15250 -9839 15252 -9787
rect 15252 -9839 15304 -9787
rect 15304 -9839 15306 -9787
rect 15250 -9841 15306 -9839
rect 15331 -9787 15387 -9785
rect 15331 -9839 15333 -9787
rect 15333 -9839 15385 -9787
rect 15385 -9839 15387 -9787
rect 15331 -9841 15387 -9839
rect 15413 -9787 15469 -9785
rect 15413 -9839 15415 -9787
rect 15415 -9839 15467 -9787
rect 15467 -9839 15469 -9787
rect 15413 -9841 15469 -9839
rect 15494 -9787 15550 -9785
rect 15494 -9839 15496 -9787
rect 15496 -9839 15548 -9787
rect 15548 -9839 15550 -9787
rect 15494 -9841 15550 -9839
rect 15575 -9787 15631 -9785
rect 15575 -9839 15577 -9787
rect 15577 -9839 15629 -9787
rect 15629 -9839 15631 -9787
rect 15575 -9841 15631 -9839
rect 15656 -9787 15712 -9785
rect 15656 -9839 15658 -9787
rect 15658 -9839 15710 -9787
rect 15710 -9839 15712 -9787
rect 15656 -9841 15712 -9839
rect 15737 -9787 15793 -9785
rect 15737 -9839 15739 -9787
rect 15739 -9839 15791 -9787
rect 15791 -9839 15793 -9787
rect 15737 -9841 15793 -9839
rect 15818 -9787 15874 -9785
rect 15818 -9839 15820 -9787
rect 15820 -9839 15872 -9787
rect 15872 -9839 15874 -9787
rect 15818 -9841 15874 -9839
rect 15899 -9787 15955 -9785
rect 15899 -9839 15901 -9787
rect 15901 -9839 15953 -9787
rect 15953 -9839 15955 -9787
rect 15899 -9841 15955 -9839
rect 15981 -9787 16037 -9785
rect 15981 -9839 15983 -9787
rect 15983 -9839 16035 -9787
rect 16035 -9839 16037 -9787
rect 15981 -9841 16037 -9839
rect 16062 -9787 16118 -9785
rect 16062 -9839 16064 -9787
rect 16064 -9839 16116 -9787
rect 16116 -9839 16118 -9787
rect 16062 -9841 16118 -9839
rect 16143 -9787 16199 -9785
rect 16143 -9839 16145 -9787
rect 16145 -9839 16197 -9787
rect 16197 -9839 16199 -9787
rect 16143 -9841 16199 -9839
rect 16224 -9787 16280 -9785
rect 16224 -9839 16226 -9787
rect 16226 -9839 16278 -9787
rect 16278 -9839 16280 -9787
rect 16224 -9841 16280 -9839
rect 16305 -9787 16361 -9785
rect 16305 -9839 16307 -9787
rect 16307 -9839 16359 -9787
rect 16359 -9839 16361 -9787
rect 16305 -9841 16361 -9839
rect 16386 -9787 16442 -9785
rect 16386 -9839 16388 -9787
rect 16388 -9839 16440 -9787
rect 16440 -9839 16442 -9787
rect 16386 -9841 16442 -9839
rect 16467 -9787 16523 -9785
rect 16467 -9839 16469 -9787
rect 16469 -9839 16521 -9787
rect 16521 -9839 16523 -9787
rect 16467 -9841 16523 -9839
rect 16549 -9787 16605 -9785
rect 16549 -9839 16551 -9787
rect 16551 -9839 16603 -9787
rect 16603 -9839 16605 -9787
rect 16549 -9841 16605 -9839
rect 16630 -9787 16686 -9785
rect 16630 -9839 16632 -9787
rect 16632 -9839 16684 -9787
rect 16684 -9839 16686 -9787
rect 16630 -9841 16686 -9839
rect 16711 -9787 16767 -9785
rect 16711 -9839 16713 -9787
rect 16713 -9839 16765 -9787
rect 16765 -9839 16767 -9787
rect 16711 -9841 16767 -9839
rect 16792 -9787 16848 -9785
rect 16792 -9839 16794 -9787
rect 16794 -9839 16846 -9787
rect 16846 -9839 16848 -9787
rect 16792 -9841 16848 -9839
rect 16873 -9787 16929 -9785
rect 16873 -9839 16875 -9787
rect 16875 -9839 16927 -9787
rect 16927 -9839 16929 -9787
rect 16873 -9841 16929 -9839
rect 16954 -9787 17010 -9785
rect 16954 -9839 16956 -9787
rect 16956 -9839 17008 -9787
rect 17008 -9839 17010 -9787
rect 16954 -9841 17010 -9839
rect 17035 -9787 17091 -9785
rect 17035 -9839 17037 -9787
rect 17037 -9839 17089 -9787
rect 17089 -9839 17091 -9787
rect 17035 -9841 17091 -9839
rect 17117 -9787 17173 -9785
rect 17117 -9839 17119 -9787
rect 17119 -9839 17171 -9787
rect 17171 -9839 17173 -9787
rect 17117 -9841 17173 -9839
rect 17198 -9787 17254 -9785
rect 17198 -9839 17200 -9787
rect 17200 -9839 17252 -9787
rect 17252 -9839 17254 -9787
rect 17198 -9841 17254 -9839
rect 17279 -9787 17335 -9785
rect 17279 -9839 17281 -9787
rect 17281 -9839 17333 -9787
rect 17333 -9839 17335 -9787
rect 17279 -9841 17335 -9839
rect 17360 -9787 17416 -9785
rect 17360 -9839 17362 -9787
rect 17362 -9839 17414 -9787
rect 17414 -9839 17416 -9787
rect 17360 -9841 17416 -9839
rect 17441 -9787 17497 -9785
rect 17441 -9839 17443 -9787
rect 17443 -9839 17495 -9787
rect 17495 -9839 17497 -9787
rect 17441 -9841 17497 -9839
rect 17522 -9787 17578 -9785
rect 17522 -9839 17524 -9787
rect 17524 -9839 17576 -9787
rect 17576 -9839 17578 -9787
rect 17522 -9841 17578 -9839
rect 17603 -9787 17659 -9785
rect 17603 -9839 17605 -9787
rect 17605 -9839 17657 -9787
rect 17657 -9839 17659 -9787
rect 17603 -9841 17659 -9839
rect 17684 -9787 17740 -9785
rect 17684 -9839 17686 -9787
rect 17686 -9839 17738 -9787
rect 17738 -9839 17740 -9787
rect 17684 -9841 17740 -9839
rect 17765 -9787 17821 -9785
rect 17765 -9839 17767 -9787
rect 17767 -9839 17819 -9787
rect 17819 -9839 17821 -9787
rect 17765 -9841 17821 -9839
rect 17846 -9787 17902 -9785
rect 17846 -9839 17848 -9787
rect 17848 -9839 17900 -9787
rect 17900 -9839 17902 -9787
rect 17846 -9841 17902 -9839
rect 17927 -9787 17983 -9785
rect 17927 -9839 17929 -9787
rect 17929 -9839 17981 -9787
rect 17981 -9839 17983 -9787
rect 17927 -9841 17983 -9839
rect 18008 -9787 18064 -9785
rect 18008 -9839 18010 -9787
rect 18010 -9839 18062 -9787
rect 18062 -9839 18064 -9787
rect 18008 -9841 18064 -9839
rect 18089 -9787 18145 -9785
rect 18089 -9839 18091 -9787
rect 18091 -9839 18143 -9787
rect 18143 -9839 18145 -9787
rect 18089 -9841 18145 -9839
rect 18171 -9787 18227 -9785
rect 18171 -9839 18173 -9787
rect 18173 -9839 18225 -9787
rect 18225 -9839 18227 -9787
rect 18171 -9841 18227 -9839
rect 18252 -9787 18308 -9785
rect 18252 -9839 18254 -9787
rect 18254 -9839 18306 -9787
rect 18306 -9839 18308 -9787
rect 18252 -9841 18308 -9839
rect 18333 -9787 18389 -9785
rect 18333 -9839 18335 -9787
rect 18335 -9839 18387 -9787
rect 18387 -9839 18389 -9787
rect 18333 -9841 18389 -9839
rect 18414 -9787 18470 -9785
rect 18414 -9839 18416 -9787
rect 18416 -9839 18468 -9787
rect 18468 -9839 18470 -9787
rect 18414 -9841 18470 -9839
rect 18495 -9787 18551 -9785
rect 18495 -9839 18497 -9787
rect 18497 -9839 18549 -9787
rect 18549 -9839 18551 -9787
rect 18495 -9841 18551 -9839
rect 18576 -9787 18632 -9785
rect 18576 -9839 18578 -9787
rect 18578 -9839 18630 -9787
rect 18630 -9839 18632 -9787
rect 18576 -9841 18632 -9839
rect 18657 -9787 18713 -9785
rect 18657 -9839 18659 -9787
rect 18659 -9839 18711 -9787
rect 18711 -9839 18713 -9787
rect 18657 -9841 18713 -9839
rect 18739 -9787 18795 -9785
rect 18739 -9839 18741 -9787
rect 18741 -9839 18793 -9787
rect 18793 -9839 18795 -9787
rect 18739 -9841 18795 -9839
rect 18820 -9787 18876 -9785
rect 18820 -9839 18822 -9787
rect 18822 -9839 18874 -9787
rect 18874 -9839 18876 -9787
rect 18820 -9841 18876 -9839
rect 18901 -9787 18957 -9785
rect 18901 -9839 18903 -9787
rect 18903 -9839 18955 -9787
rect 18955 -9839 18957 -9787
rect 18901 -9841 18957 -9839
rect 18982 -9787 19038 -9785
rect 18982 -9839 18984 -9787
rect 18984 -9839 19036 -9787
rect 19036 -9839 19038 -9787
rect 18982 -9841 19038 -9839
rect 19063 -9787 19119 -9785
rect 19063 -9839 19065 -9787
rect 19065 -9839 19117 -9787
rect 19117 -9839 19119 -9787
rect 19063 -9841 19119 -9839
rect 19144 -9787 19200 -9785
rect 19144 -9839 19146 -9787
rect 19146 -9839 19198 -9787
rect 19198 -9839 19200 -9787
rect 19144 -9841 19200 -9839
rect 19225 -9787 19281 -9785
rect 19225 -9839 19227 -9787
rect 19227 -9839 19279 -9787
rect 19279 -9839 19281 -9787
rect 19225 -9841 19281 -9839
rect 19307 -9787 19363 -9785
rect 19307 -9839 19309 -9787
rect 19309 -9839 19361 -9787
rect 19361 -9839 19363 -9787
rect 19307 -9841 19363 -9839
rect 19388 -9787 19444 -9785
rect 19388 -9839 19390 -9787
rect 19390 -9839 19442 -9787
rect 19442 -9839 19444 -9787
rect 19388 -9841 19444 -9839
rect 19469 -9787 19525 -9785
rect 19469 -9839 19471 -9787
rect 19471 -9839 19523 -9787
rect 19523 -9839 19525 -9787
rect 19469 -9841 19525 -9839
rect 19550 -9787 19606 -9785
rect 19550 -9839 19552 -9787
rect 19552 -9839 19604 -9787
rect 19604 -9839 19606 -9787
rect 19550 -9841 19606 -9839
rect 19631 -9787 19687 -9785
rect 19631 -9839 19633 -9787
rect 19633 -9839 19685 -9787
rect 19685 -9839 19687 -9787
rect 19631 -9841 19687 -9839
rect 19712 -9787 19768 -9785
rect 19712 -9839 19714 -9787
rect 19714 -9839 19766 -9787
rect 19766 -9839 19768 -9787
rect 19712 -9841 19768 -9839
rect 19793 -9787 19849 -9785
rect 19793 -9839 19795 -9787
rect 19795 -9839 19847 -9787
rect 19847 -9839 19849 -9787
rect 19793 -9841 19849 -9839
rect 19875 -9787 19931 -9785
rect 19875 -9839 19877 -9787
rect 19877 -9839 19929 -9787
rect 19929 -9839 19931 -9787
rect 19875 -9841 19931 -9839
rect 19956 -9787 20012 -9785
rect 19956 -9839 19958 -9787
rect 19958 -9839 20010 -9787
rect 20010 -9839 20012 -9787
rect 19956 -9841 20012 -9839
rect 20037 -9787 20093 -9785
rect 20037 -9839 20039 -9787
rect 20039 -9839 20091 -9787
rect 20091 -9839 20093 -9787
rect 20037 -9841 20093 -9839
rect 20118 -9787 20174 -9785
rect 20118 -9839 20120 -9787
rect 20120 -9839 20172 -9787
rect 20172 -9839 20174 -9787
rect 20118 -9841 20174 -9839
rect 20199 -9787 20255 -9785
rect 20199 -9839 20201 -9787
rect 20201 -9839 20253 -9787
rect 20253 -9839 20255 -9787
rect 20199 -9841 20255 -9839
rect 20280 -9787 20336 -9785
rect 20280 -9839 20282 -9787
rect 20282 -9839 20334 -9787
rect 20334 -9839 20336 -9787
rect 20280 -9841 20336 -9839
rect 20361 -9787 20417 -9785
rect 20361 -9839 20363 -9787
rect 20363 -9839 20415 -9787
rect 20415 -9839 20417 -9787
rect 20361 -9841 20417 -9839
rect 20443 -9787 20499 -9785
rect 20443 -9839 20445 -9787
rect 20445 -9839 20497 -9787
rect 20497 -9839 20499 -9787
rect 20443 -9841 20499 -9839
rect 20524 -9787 20580 -9785
rect 20524 -9839 20526 -9787
rect 20526 -9839 20578 -9787
rect 20578 -9839 20580 -9787
rect 20524 -9841 20580 -9839
rect 20605 -9787 20661 -9785
rect 20605 -9839 20607 -9787
rect 20607 -9839 20659 -9787
rect 20659 -9839 20661 -9787
rect 20605 -9841 20661 -9839
rect 20686 -9787 20742 -9785
rect 20686 -9839 20688 -9787
rect 20688 -9839 20740 -9787
rect 20740 -9839 20742 -9787
rect 20686 -9841 20742 -9839
rect 20767 -9787 20823 -9785
rect 20767 -9839 20769 -9787
rect 20769 -9839 20821 -9787
rect 20821 -9839 20823 -9787
rect 20767 -9841 20823 -9839
rect 20848 -9787 20904 -9785
rect 20848 -9839 20850 -9787
rect 20850 -9839 20902 -9787
rect 20902 -9839 20904 -9787
rect 20848 -9841 20904 -9839
rect 20929 -9787 20985 -9785
rect 20929 -9839 20931 -9787
rect 20931 -9839 20983 -9787
rect 20983 -9839 20985 -9787
rect 20929 -9841 20985 -9839
rect 21011 -9787 21067 -9785
rect 21011 -9839 21013 -9787
rect 21013 -9839 21065 -9787
rect 21065 -9839 21067 -9787
rect 21011 -9841 21067 -9839
rect 21092 -9787 21148 -9785
rect 21092 -9839 21094 -9787
rect 21094 -9839 21146 -9787
rect 21146 -9839 21148 -9787
rect 21092 -9841 21148 -9839
rect 21173 -9787 21229 -9785
rect 21173 -9839 21175 -9787
rect 21175 -9839 21227 -9787
rect 21227 -9839 21229 -9787
rect 21173 -9841 21229 -9839
rect 21254 -9787 21310 -9785
rect 21254 -9839 21256 -9787
rect 21256 -9839 21308 -9787
rect 21308 -9839 21310 -9787
rect 21254 -9841 21310 -9839
rect 21335 -9787 21391 -9785
rect 21335 -9839 21337 -9787
rect 21337 -9839 21389 -9787
rect 21389 -9839 21391 -9787
rect 21335 -9841 21391 -9839
rect 21416 -9787 21472 -9785
rect 21416 -9839 21418 -9787
rect 21418 -9839 21470 -9787
rect 21470 -9839 21472 -9787
rect 21416 -9841 21472 -9839
rect 21497 -9787 21553 -9785
rect 21497 -9839 21499 -9787
rect 21499 -9839 21551 -9787
rect 21551 -9839 21553 -9787
rect 21497 -9841 21553 -9839
rect 21579 -9787 21635 -9785
rect 21579 -9839 21581 -9787
rect 21581 -9839 21633 -9787
rect 21633 -9839 21635 -9787
rect 21579 -9841 21635 -9839
rect 21660 -9787 21716 -9785
rect 21660 -9839 21662 -9787
rect 21662 -9839 21714 -9787
rect 21714 -9839 21716 -9787
rect 21660 -9841 21716 -9839
rect 21741 -9787 21797 -9785
rect 21741 -9839 21743 -9787
rect 21743 -9839 21795 -9787
rect 21795 -9839 21797 -9787
rect 21741 -9841 21797 -9839
rect 21822 -9787 21878 -9785
rect 21822 -9839 21824 -9787
rect 21824 -9839 21876 -9787
rect 21876 -9839 21878 -9787
rect 21822 -9841 21878 -9839
rect 21903 -9787 21959 -9785
rect 21903 -9839 21905 -9787
rect 21905 -9839 21957 -9787
rect 21957 -9839 21959 -9787
rect 21903 -9841 21959 -9839
rect 21984 -9787 22040 -9785
rect 21984 -9839 21986 -9787
rect 21986 -9839 22038 -9787
rect 22038 -9839 22040 -9787
rect 21984 -9841 22040 -9839
rect 22065 -9787 22121 -9785
rect 22065 -9839 22067 -9787
rect 22067 -9839 22119 -9787
rect 22119 -9839 22121 -9787
rect 22065 -9841 22121 -9839
rect 22147 -9787 22203 -9785
rect 22147 -9839 22149 -9787
rect 22149 -9839 22201 -9787
rect 22201 -9839 22203 -9787
rect 22147 -9841 22203 -9839
rect 22228 -9787 22284 -9785
rect 22228 -9839 22230 -9787
rect 22230 -9839 22282 -9787
rect 22282 -9839 22284 -9787
rect 22228 -9841 22284 -9839
rect 22309 -9787 22365 -9785
rect 22309 -9839 22311 -9787
rect 22311 -9839 22363 -9787
rect 22363 -9839 22365 -9787
rect 22309 -9841 22365 -9839
rect 22390 -9787 22446 -9785
rect 22390 -9839 22392 -9787
rect 22392 -9839 22444 -9787
rect 22444 -9839 22446 -9787
rect 22390 -9841 22446 -9839
rect 22471 -9787 22527 -9785
rect 22471 -9839 22473 -9787
rect 22473 -9839 22525 -9787
rect 22525 -9839 22527 -9787
rect 22471 -9841 22527 -9839
rect 22552 -9787 22608 -9785
rect 22552 -9839 22554 -9787
rect 22554 -9839 22606 -9787
rect 22606 -9839 22608 -9787
rect 22552 -9841 22608 -9839
rect 22633 -9787 22689 -9785
rect 22633 -9839 22635 -9787
rect 22635 -9839 22687 -9787
rect 22687 -9839 22689 -9787
rect 22633 -9841 22689 -9839
rect 22715 -9787 22771 -9785
rect 22715 -9839 22717 -9787
rect 22717 -9839 22769 -9787
rect 22769 -9839 22771 -9787
rect 22715 -9841 22771 -9839
rect 22796 -9787 22852 -9785
rect 22796 -9839 22798 -9787
rect 22798 -9839 22850 -9787
rect 22850 -9839 22852 -9787
rect 22796 -9841 22852 -9839
rect 22877 -9787 22933 -9785
rect 22877 -9839 22879 -9787
rect 22879 -9839 22931 -9787
rect 22931 -9839 22933 -9787
rect 22877 -9841 22933 -9839
rect 22958 -9787 23014 -9785
rect 22958 -9839 22960 -9787
rect 22960 -9839 23012 -9787
rect 23012 -9839 23014 -9787
rect 22958 -9841 23014 -9839
rect 23039 -9787 23095 -9785
rect 23039 -9839 23041 -9787
rect 23041 -9839 23093 -9787
rect 23093 -9839 23095 -9787
rect 23039 -9841 23095 -9839
rect 23120 -9787 23176 -9785
rect 23120 -9839 23122 -9787
rect 23122 -9839 23174 -9787
rect 23174 -9839 23176 -9787
rect 23120 -9841 23176 -9839
rect 23201 -9787 23257 -9785
rect 23201 -9839 23203 -9787
rect 23203 -9839 23255 -9787
rect 23255 -9839 23257 -9787
rect 23201 -9841 23257 -9839
rect 23283 -9787 23339 -9785
rect 23283 -9839 23285 -9787
rect 23285 -9839 23337 -9787
rect 23337 -9839 23339 -9787
rect 23283 -9841 23339 -9839
rect 23364 -9787 23420 -9785
rect 23364 -9839 23366 -9787
rect 23366 -9839 23418 -9787
rect 23418 -9839 23420 -9787
rect 23364 -9841 23420 -9839
rect 23445 -9787 23501 -9785
rect 23445 -9839 23447 -9787
rect 23447 -9839 23499 -9787
rect 23499 -9839 23501 -9787
rect 23445 -9841 23501 -9839
rect 23526 -9787 23582 -9785
rect 23526 -9839 23528 -9787
rect 23528 -9839 23580 -9787
rect 23580 -9839 23582 -9787
rect 23526 -9841 23582 -9839
rect 23607 -9787 23663 -9785
rect 23607 -9839 23609 -9787
rect 23609 -9839 23661 -9787
rect 23661 -9839 23663 -9787
rect 23607 -9841 23663 -9839
rect 23688 -9787 23744 -9785
rect 23688 -9839 23690 -9787
rect 23690 -9839 23742 -9787
rect 23742 -9839 23744 -9787
rect 23688 -9841 23744 -9839
rect 23769 -9787 23825 -9785
rect 23769 -9839 23771 -9787
rect 23771 -9839 23823 -9787
rect 23823 -9839 23825 -9787
rect 23769 -9841 23825 -9839
rect 23851 -9787 23907 -9785
rect 23851 -9839 23853 -9787
rect 23853 -9839 23905 -9787
rect 23905 -9839 23907 -9787
rect 23851 -9841 23907 -9839
rect 23932 -9787 23988 -9785
rect 23932 -9839 23934 -9787
rect 23934 -9839 23986 -9787
rect 23986 -9839 23988 -9787
rect 23932 -9841 23988 -9839
rect 24013 -9787 24069 -9785
rect 24013 -9839 24015 -9787
rect 24015 -9839 24067 -9787
rect 24067 -9839 24069 -9787
rect 24013 -9841 24069 -9839
rect 24094 -9787 24150 -9785
rect 24094 -9839 24096 -9787
rect 24096 -9839 24148 -9787
rect 24148 -9839 24150 -9787
rect 24094 -9841 24150 -9839
rect 24175 -9787 24231 -9785
rect 24175 -9839 24177 -9787
rect 24177 -9839 24229 -9787
rect 24229 -9839 24231 -9787
rect 24175 -9841 24231 -9839
rect 24256 -9787 24312 -9785
rect 24256 -9839 24258 -9787
rect 24258 -9839 24310 -9787
rect 24310 -9839 24312 -9787
rect 24256 -9841 24312 -9839
rect 24337 -9787 24393 -9785
rect 24337 -9839 24339 -9787
rect 24339 -9839 24391 -9787
rect 24391 -9839 24393 -9787
rect 24337 -9841 24393 -9839
rect 24419 -9787 24475 -9785
rect 24419 -9839 24421 -9787
rect 24421 -9839 24473 -9787
rect 24473 -9839 24475 -9787
rect 24419 -9841 24475 -9839
rect 24500 -9787 24556 -9785
rect 24500 -9839 24502 -9787
rect 24502 -9839 24554 -9787
rect 24554 -9839 24556 -9787
rect 24500 -9841 24556 -9839
rect 24581 -9787 24637 -9785
rect 24581 -9839 24583 -9787
rect 24583 -9839 24635 -9787
rect 24635 -9839 24637 -9787
rect 24581 -9841 24637 -9839
rect 24662 -9787 24718 -9785
rect 24662 -9839 24664 -9787
rect 24664 -9839 24716 -9787
rect 24716 -9839 24718 -9787
rect 24662 -9841 24718 -9839
rect 24743 -9787 24799 -9785
rect 24743 -9839 24745 -9787
rect 24745 -9839 24797 -9787
rect 24797 -9839 24799 -9787
rect 24743 -9841 24799 -9839
rect 24824 -9787 24880 -9785
rect 24824 -9839 24826 -9787
rect 24826 -9839 24878 -9787
rect 24878 -9839 24880 -9787
rect 24824 -9841 24880 -9839
rect 24905 -9787 24961 -9785
rect 24905 -9839 24907 -9787
rect 24907 -9839 24959 -9787
rect 24959 -9839 24961 -9787
rect 24905 -9841 24961 -9839
rect 24987 -9787 25043 -9785
rect 24987 -9839 24989 -9787
rect 24989 -9839 25041 -9787
rect 25041 -9839 25043 -9787
rect 24987 -9841 25043 -9839
rect 25068 -9787 25124 -9785
rect 25068 -9839 25070 -9787
rect 25070 -9839 25122 -9787
rect 25122 -9839 25124 -9787
rect 25068 -9841 25124 -9839
rect 25149 -9787 25205 -9785
rect 25149 -9839 25151 -9787
rect 25151 -9839 25203 -9787
rect 25203 -9839 25205 -9787
rect 25149 -9841 25205 -9839
rect 25230 -9787 25286 -9785
rect 25230 -9839 25232 -9787
rect 25232 -9839 25284 -9787
rect 25284 -9839 25286 -9787
rect 25230 -9841 25286 -9839
rect 25311 -9787 25367 -9785
rect 25311 -9839 25313 -9787
rect 25313 -9839 25365 -9787
rect 25365 -9839 25367 -9787
rect 25311 -9841 25367 -9839
rect 25392 -9787 25448 -9785
rect 25392 -9839 25394 -9787
rect 25394 -9839 25446 -9787
rect 25446 -9839 25448 -9787
rect 25392 -9841 25448 -9839
rect 25473 -9787 25529 -9785
rect 25473 -9839 25475 -9787
rect 25475 -9839 25527 -9787
rect 25527 -9839 25529 -9787
rect 25473 -9841 25529 -9839
rect 25555 -9787 25611 -9785
rect 25555 -9839 25557 -9787
rect 25557 -9839 25609 -9787
rect 25609 -9839 25611 -9787
rect 25555 -9841 25611 -9839
rect 25636 -9787 25692 -9785
rect 25636 -9839 25638 -9787
rect 25638 -9839 25690 -9787
rect 25690 -9839 25692 -9787
rect 25636 -9841 25692 -9839
rect 25717 -9787 25773 -9785
rect 25717 -9839 25719 -9787
rect 25719 -9839 25771 -9787
rect 25771 -9839 25773 -9787
rect 25717 -9841 25773 -9839
rect 25798 -9787 25854 -9785
rect 25798 -9839 25800 -9787
rect 25800 -9839 25852 -9787
rect 25852 -9839 25854 -9787
rect 25798 -9841 25854 -9839
rect 25879 -9787 25935 -9785
rect 25879 -9839 25881 -9787
rect 25881 -9839 25933 -9787
rect 25933 -9839 25935 -9787
rect 25879 -9841 25935 -9839
rect 25960 -9787 26016 -9785
rect 25960 -9839 25962 -9787
rect 25962 -9839 26014 -9787
rect 26014 -9839 26016 -9787
rect 25960 -9841 26016 -9839
rect 26041 -9787 26097 -9785
rect 26041 -9839 26043 -9787
rect 26043 -9839 26095 -9787
rect 26095 -9839 26097 -9787
rect 26041 -9841 26097 -9839
rect 26123 -9787 26179 -9785
rect 26123 -9839 26125 -9787
rect 26125 -9839 26177 -9787
rect 26177 -9839 26179 -9787
rect 26123 -9841 26179 -9839
rect 26204 -9787 26260 -9785
rect 26204 -9839 26206 -9787
rect 26206 -9839 26258 -9787
rect 26258 -9839 26260 -9787
rect 26204 -9841 26260 -9839
rect 4053 -9891 4109 -9889
rect 4053 -9943 4055 -9891
rect 4055 -9943 4107 -9891
rect 4107 -9943 4109 -9891
rect 4053 -9945 4109 -9943
rect 4134 -9891 4190 -9889
rect 4134 -9943 4136 -9891
rect 4136 -9943 4188 -9891
rect 4188 -9943 4190 -9891
rect 4134 -9945 4190 -9943
rect 4215 -9891 4271 -9889
rect 4215 -9943 4217 -9891
rect 4217 -9943 4269 -9891
rect 4269 -9943 4271 -9891
rect 4215 -9945 4271 -9943
rect 4296 -9891 4352 -9889
rect 4296 -9943 4298 -9891
rect 4298 -9943 4350 -9891
rect 4350 -9943 4352 -9891
rect 4296 -9945 4352 -9943
rect 4377 -9891 4433 -9889
rect 4377 -9943 4379 -9891
rect 4379 -9943 4431 -9891
rect 4431 -9943 4433 -9891
rect 4377 -9945 4433 -9943
rect 4458 -9891 4514 -9889
rect 4458 -9943 4460 -9891
rect 4460 -9943 4512 -9891
rect 4512 -9943 4514 -9891
rect 4458 -9945 4514 -9943
rect 4539 -9891 4595 -9889
rect 4539 -9943 4541 -9891
rect 4541 -9943 4593 -9891
rect 4593 -9943 4595 -9891
rect 4539 -9945 4595 -9943
rect 4621 -9891 4677 -9889
rect 4621 -9943 4623 -9891
rect 4623 -9943 4675 -9891
rect 4675 -9943 4677 -9891
rect 4621 -9945 4677 -9943
rect 4702 -9891 4758 -9889
rect 4702 -9943 4704 -9891
rect 4704 -9943 4756 -9891
rect 4756 -9943 4758 -9891
rect 4702 -9945 4758 -9943
rect 4783 -9891 4839 -9889
rect 4783 -9943 4785 -9891
rect 4785 -9943 4837 -9891
rect 4837 -9943 4839 -9891
rect 4783 -9945 4839 -9943
rect 4864 -9891 4920 -9889
rect 4864 -9943 4866 -9891
rect 4866 -9943 4918 -9891
rect 4918 -9943 4920 -9891
rect 4864 -9945 4920 -9943
rect 4945 -9891 5001 -9889
rect 4945 -9943 4947 -9891
rect 4947 -9943 4999 -9891
rect 4999 -9943 5001 -9891
rect 4945 -9945 5001 -9943
rect 5026 -9891 5082 -9889
rect 5026 -9943 5028 -9891
rect 5028 -9943 5080 -9891
rect 5080 -9943 5082 -9891
rect 5026 -9945 5082 -9943
rect 5107 -9891 5163 -9889
rect 5107 -9943 5109 -9891
rect 5109 -9943 5161 -9891
rect 5161 -9943 5163 -9891
rect 5107 -9945 5163 -9943
rect 5189 -9891 5245 -9889
rect 5189 -9943 5191 -9891
rect 5191 -9943 5243 -9891
rect 5243 -9943 5245 -9891
rect 5189 -9945 5245 -9943
rect 5270 -9891 5326 -9889
rect 5270 -9943 5272 -9891
rect 5272 -9943 5324 -9891
rect 5324 -9943 5326 -9891
rect 5270 -9945 5326 -9943
rect 5351 -9891 5407 -9889
rect 5351 -9943 5353 -9891
rect 5353 -9943 5405 -9891
rect 5405 -9943 5407 -9891
rect 5351 -9945 5407 -9943
rect 5432 -9891 5488 -9889
rect 5432 -9943 5434 -9891
rect 5434 -9943 5486 -9891
rect 5486 -9943 5488 -9891
rect 5432 -9945 5488 -9943
rect 5513 -9891 5569 -9889
rect 5513 -9943 5515 -9891
rect 5515 -9943 5567 -9891
rect 5567 -9943 5569 -9891
rect 5513 -9945 5569 -9943
rect 5594 -9891 5650 -9889
rect 5594 -9943 5596 -9891
rect 5596 -9943 5648 -9891
rect 5648 -9943 5650 -9891
rect 5594 -9945 5650 -9943
rect 5675 -9891 5731 -9889
rect 5675 -9943 5677 -9891
rect 5677 -9943 5729 -9891
rect 5729 -9943 5731 -9891
rect 5675 -9945 5731 -9943
rect 5757 -9891 5813 -9889
rect 5757 -9943 5759 -9891
rect 5759 -9943 5811 -9891
rect 5811 -9943 5813 -9891
rect 5757 -9945 5813 -9943
rect 5838 -9891 5894 -9889
rect 5838 -9943 5840 -9891
rect 5840 -9943 5892 -9891
rect 5892 -9943 5894 -9891
rect 5838 -9945 5894 -9943
rect 5919 -9891 5975 -9889
rect 5919 -9943 5921 -9891
rect 5921 -9943 5973 -9891
rect 5973 -9943 5975 -9891
rect 5919 -9945 5975 -9943
rect 6000 -9891 6056 -9889
rect 6000 -9943 6002 -9891
rect 6002 -9943 6054 -9891
rect 6054 -9943 6056 -9891
rect 6000 -9945 6056 -9943
rect 6081 -9891 6137 -9889
rect 6081 -9943 6083 -9891
rect 6083 -9943 6135 -9891
rect 6135 -9943 6137 -9891
rect 6081 -9945 6137 -9943
rect 6162 -9891 6218 -9889
rect 6162 -9943 6164 -9891
rect 6164 -9943 6216 -9891
rect 6216 -9943 6218 -9891
rect 6162 -9945 6218 -9943
rect 6243 -9891 6299 -9889
rect 6243 -9943 6245 -9891
rect 6245 -9943 6297 -9891
rect 6297 -9943 6299 -9891
rect 6243 -9945 6299 -9943
rect 6325 -9891 6381 -9889
rect 6325 -9943 6327 -9891
rect 6327 -9943 6379 -9891
rect 6379 -9943 6381 -9891
rect 6325 -9945 6381 -9943
rect 6406 -9891 6462 -9889
rect 6406 -9943 6408 -9891
rect 6408 -9943 6460 -9891
rect 6460 -9943 6462 -9891
rect 6406 -9945 6462 -9943
rect 6487 -9891 6543 -9889
rect 6487 -9943 6489 -9891
rect 6489 -9943 6541 -9891
rect 6541 -9943 6543 -9891
rect 6487 -9945 6543 -9943
rect 6568 -9891 6624 -9889
rect 6568 -9943 6570 -9891
rect 6570 -9943 6622 -9891
rect 6622 -9943 6624 -9891
rect 6568 -9945 6624 -9943
rect 6649 -9891 6705 -9889
rect 6649 -9943 6651 -9891
rect 6651 -9943 6703 -9891
rect 6703 -9943 6705 -9891
rect 6649 -9945 6705 -9943
rect 6730 -9891 6786 -9889
rect 6730 -9943 6732 -9891
rect 6732 -9943 6784 -9891
rect 6784 -9943 6786 -9891
rect 6730 -9945 6786 -9943
rect 6811 -9891 6867 -9889
rect 6811 -9943 6813 -9891
rect 6813 -9943 6865 -9891
rect 6865 -9943 6867 -9891
rect 6811 -9945 6867 -9943
rect 6893 -9891 6949 -9889
rect 6893 -9943 6895 -9891
rect 6895 -9943 6947 -9891
rect 6947 -9943 6949 -9891
rect 6893 -9945 6949 -9943
rect 6974 -9891 7030 -9889
rect 6974 -9943 6976 -9891
rect 6976 -9943 7028 -9891
rect 7028 -9943 7030 -9891
rect 6974 -9945 7030 -9943
rect 7055 -9891 7111 -9889
rect 7055 -9943 7057 -9891
rect 7057 -9943 7109 -9891
rect 7109 -9943 7111 -9891
rect 7055 -9945 7111 -9943
rect 7136 -9891 7192 -9889
rect 7136 -9943 7138 -9891
rect 7138 -9943 7190 -9891
rect 7190 -9943 7192 -9891
rect 7136 -9945 7192 -9943
rect 7217 -9891 7273 -9889
rect 7217 -9943 7219 -9891
rect 7219 -9943 7271 -9891
rect 7271 -9943 7273 -9891
rect 7217 -9945 7273 -9943
rect 7298 -9891 7354 -9889
rect 7298 -9943 7300 -9891
rect 7300 -9943 7352 -9891
rect 7352 -9943 7354 -9891
rect 7298 -9945 7354 -9943
rect 7379 -9891 7435 -9889
rect 7379 -9943 7381 -9891
rect 7381 -9943 7433 -9891
rect 7433 -9943 7435 -9891
rect 7379 -9945 7435 -9943
rect 7461 -9891 7517 -9889
rect 7461 -9943 7463 -9891
rect 7463 -9943 7515 -9891
rect 7515 -9943 7517 -9891
rect 7461 -9945 7517 -9943
rect 7542 -9891 7598 -9889
rect 7542 -9943 7544 -9891
rect 7544 -9943 7596 -9891
rect 7596 -9943 7598 -9891
rect 7542 -9945 7598 -9943
rect 7623 -9891 7679 -9889
rect 7623 -9943 7625 -9891
rect 7625 -9943 7677 -9891
rect 7677 -9943 7679 -9891
rect 7623 -9945 7679 -9943
rect 7704 -9891 7760 -9889
rect 7704 -9943 7706 -9891
rect 7706 -9943 7758 -9891
rect 7758 -9943 7760 -9891
rect 7704 -9945 7760 -9943
rect 7785 -9891 7841 -9889
rect 7785 -9943 7787 -9891
rect 7787 -9943 7839 -9891
rect 7839 -9943 7841 -9891
rect 7785 -9945 7841 -9943
rect 7866 -9891 7922 -9889
rect 7866 -9943 7868 -9891
rect 7868 -9943 7920 -9891
rect 7920 -9943 7922 -9891
rect 7866 -9945 7922 -9943
rect 7947 -9891 8003 -9889
rect 7947 -9943 7949 -9891
rect 7949 -9943 8001 -9891
rect 8001 -9943 8003 -9891
rect 7947 -9945 8003 -9943
rect 8029 -9891 8085 -9889
rect 8029 -9943 8031 -9891
rect 8031 -9943 8083 -9891
rect 8083 -9943 8085 -9891
rect 8029 -9945 8085 -9943
rect 8110 -9891 8166 -9889
rect 8110 -9943 8112 -9891
rect 8112 -9943 8164 -9891
rect 8164 -9943 8166 -9891
rect 8110 -9945 8166 -9943
rect 8191 -9891 8247 -9889
rect 8191 -9943 8193 -9891
rect 8193 -9943 8245 -9891
rect 8245 -9943 8247 -9891
rect 8191 -9945 8247 -9943
rect 8272 -9891 8328 -9889
rect 8272 -9943 8274 -9891
rect 8274 -9943 8326 -9891
rect 8326 -9943 8328 -9891
rect 8272 -9945 8328 -9943
rect 8353 -9891 8409 -9889
rect 8353 -9943 8355 -9891
rect 8355 -9943 8407 -9891
rect 8407 -9943 8409 -9891
rect 8353 -9945 8409 -9943
rect 8434 -9891 8490 -9889
rect 8434 -9943 8436 -9891
rect 8436 -9943 8488 -9891
rect 8488 -9943 8490 -9891
rect 8434 -9945 8490 -9943
rect 8515 -9891 8571 -9889
rect 8515 -9943 8517 -9891
rect 8517 -9943 8569 -9891
rect 8569 -9943 8571 -9891
rect 8515 -9945 8571 -9943
rect 8597 -9891 8653 -9889
rect 8597 -9943 8599 -9891
rect 8599 -9943 8651 -9891
rect 8651 -9943 8653 -9891
rect 8597 -9945 8653 -9943
rect 8678 -9891 8734 -9889
rect 8678 -9943 8680 -9891
rect 8680 -9943 8732 -9891
rect 8732 -9943 8734 -9891
rect 8678 -9945 8734 -9943
rect 8759 -9891 8815 -9889
rect 8759 -9943 8761 -9891
rect 8761 -9943 8813 -9891
rect 8813 -9943 8815 -9891
rect 8759 -9945 8815 -9943
rect 8840 -9891 8896 -9889
rect 8840 -9943 8842 -9891
rect 8842 -9943 8894 -9891
rect 8894 -9943 8896 -9891
rect 8840 -9945 8896 -9943
rect 8921 -9891 8977 -9889
rect 8921 -9943 8923 -9891
rect 8923 -9943 8975 -9891
rect 8975 -9943 8977 -9891
rect 8921 -9945 8977 -9943
rect 9002 -9891 9058 -9889
rect 9002 -9943 9004 -9891
rect 9004 -9943 9056 -9891
rect 9056 -9943 9058 -9891
rect 9002 -9945 9058 -9943
rect 9083 -9891 9139 -9889
rect 9083 -9943 9085 -9891
rect 9085 -9943 9137 -9891
rect 9137 -9943 9139 -9891
rect 9083 -9945 9139 -9943
rect 9165 -9891 9221 -9889
rect 9165 -9943 9167 -9891
rect 9167 -9943 9219 -9891
rect 9219 -9943 9221 -9891
rect 9165 -9945 9221 -9943
rect 9246 -9891 9302 -9889
rect 9246 -9943 9248 -9891
rect 9248 -9943 9300 -9891
rect 9300 -9943 9302 -9891
rect 9246 -9945 9302 -9943
rect 9327 -9891 9383 -9889
rect 9327 -9943 9329 -9891
rect 9329 -9943 9381 -9891
rect 9381 -9943 9383 -9891
rect 9327 -9945 9383 -9943
rect 9408 -9891 9464 -9889
rect 9408 -9943 9410 -9891
rect 9410 -9943 9462 -9891
rect 9462 -9943 9464 -9891
rect 9408 -9945 9464 -9943
rect 9489 -9891 9545 -9889
rect 9489 -9943 9491 -9891
rect 9491 -9943 9543 -9891
rect 9543 -9943 9545 -9891
rect 9489 -9945 9545 -9943
rect 9570 -9891 9626 -9889
rect 9570 -9943 9572 -9891
rect 9572 -9943 9624 -9891
rect 9624 -9943 9626 -9891
rect 9570 -9945 9626 -9943
rect 9651 -9891 9707 -9889
rect 9651 -9943 9653 -9891
rect 9653 -9943 9705 -9891
rect 9705 -9943 9707 -9891
rect 9651 -9945 9707 -9943
rect 9733 -9891 9789 -9889
rect 9733 -9943 9735 -9891
rect 9735 -9943 9787 -9891
rect 9787 -9943 9789 -9891
rect 9733 -9945 9789 -9943
rect 9814 -9891 9870 -9889
rect 9814 -9943 9816 -9891
rect 9816 -9943 9868 -9891
rect 9868 -9943 9870 -9891
rect 9814 -9945 9870 -9943
rect 9895 -9891 9951 -9889
rect 9895 -9943 9897 -9891
rect 9897 -9943 9949 -9891
rect 9949 -9943 9951 -9891
rect 9895 -9945 9951 -9943
rect 9976 -9891 10032 -9889
rect 9976 -9943 9978 -9891
rect 9978 -9943 10030 -9891
rect 10030 -9943 10032 -9891
rect 9976 -9945 10032 -9943
rect 10057 -9891 10113 -9889
rect 10057 -9943 10059 -9891
rect 10059 -9943 10111 -9891
rect 10111 -9943 10113 -9891
rect 10057 -9945 10113 -9943
rect 10138 -9891 10194 -9889
rect 10138 -9943 10140 -9891
rect 10140 -9943 10192 -9891
rect 10192 -9943 10194 -9891
rect 10138 -9945 10194 -9943
rect 10219 -9891 10275 -9889
rect 10219 -9943 10221 -9891
rect 10221 -9943 10273 -9891
rect 10273 -9943 10275 -9891
rect 10219 -9945 10275 -9943
rect 10301 -9891 10357 -9889
rect 10301 -9943 10303 -9891
rect 10303 -9943 10355 -9891
rect 10355 -9943 10357 -9891
rect 10301 -9945 10357 -9943
rect 10382 -9891 10438 -9889
rect 10382 -9943 10384 -9891
rect 10384 -9943 10436 -9891
rect 10436 -9943 10438 -9891
rect 10382 -9945 10438 -9943
rect 10463 -9891 10519 -9889
rect 10463 -9943 10465 -9891
rect 10465 -9943 10517 -9891
rect 10517 -9943 10519 -9891
rect 10463 -9945 10519 -9943
rect 10544 -9891 10600 -9889
rect 10544 -9943 10546 -9891
rect 10546 -9943 10598 -9891
rect 10598 -9943 10600 -9891
rect 10544 -9945 10600 -9943
rect 10625 -9891 10681 -9889
rect 10625 -9943 10627 -9891
rect 10627 -9943 10679 -9891
rect 10679 -9943 10681 -9891
rect 10625 -9945 10681 -9943
rect 10706 -9891 10762 -9889
rect 10706 -9943 10708 -9891
rect 10708 -9943 10760 -9891
rect 10760 -9943 10762 -9891
rect 10706 -9945 10762 -9943
rect 10787 -9891 10843 -9889
rect 10787 -9943 10789 -9891
rect 10789 -9943 10841 -9891
rect 10841 -9943 10843 -9891
rect 10787 -9945 10843 -9943
rect 10869 -9891 10925 -9889
rect 10869 -9943 10871 -9891
rect 10871 -9943 10923 -9891
rect 10923 -9943 10925 -9891
rect 10869 -9945 10925 -9943
rect 10950 -9891 11006 -9889
rect 10950 -9943 10952 -9891
rect 10952 -9943 11004 -9891
rect 11004 -9943 11006 -9891
rect 10950 -9945 11006 -9943
rect 11031 -9891 11087 -9889
rect 11031 -9943 11033 -9891
rect 11033 -9943 11085 -9891
rect 11085 -9943 11087 -9891
rect 11031 -9945 11087 -9943
rect 11112 -9891 11168 -9889
rect 11112 -9943 11114 -9891
rect 11114 -9943 11166 -9891
rect 11166 -9943 11168 -9891
rect 11112 -9945 11168 -9943
rect 11193 -9891 11249 -9889
rect 11193 -9943 11195 -9891
rect 11195 -9943 11247 -9891
rect 11247 -9943 11249 -9891
rect 11193 -9945 11249 -9943
rect 11274 -9891 11330 -9889
rect 11274 -9943 11276 -9891
rect 11276 -9943 11328 -9891
rect 11328 -9943 11330 -9891
rect 11274 -9945 11330 -9943
rect 11355 -9891 11411 -9889
rect 11355 -9943 11357 -9891
rect 11357 -9943 11409 -9891
rect 11409 -9943 11411 -9891
rect 11355 -9945 11411 -9943
rect 11437 -9891 11493 -9889
rect 11437 -9943 11439 -9891
rect 11439 -9943 11491 -9891
rect 11491 -9943 11493 -9891
rect 11437 -9945 11493 -9943
rect 11518 -9891 11574 -9889
rect 11518 -9943 11520 -9891
rect 11520 -9943 11572 -9891
rect 11572 -9943 11574 -9891
rect 11518 -9945 11574 -9943
rect 11599 -9891 11655 -9889
rect 11599 -9943 11601 -9891
rect 11601 -9943 11653 -9891
rect 11653 -9943 11655 -9891
rect 11599 -9945 11655 -9943
rect 11680 -9891 11736 -9889
rect 11680 -9943 11682 -9891
rect 11682 -9943 11734 -9891
rect 11734 -9943 11736 -9891
rect 11680 -9945 11736 -9943
rect 11761 -9891 11817 -9889
rect 11761 -9943 11763 -9891
rect 11763 -9943 11815 -9891
rect 11815 -9943 11817 -9891
rect 11761 -9945 11817 -9943
rect 11842 -9891 11898 -9889
rect 11842 -9943 11844 -9891
rect 11844 -9943 11896 -9891
rect 11896 -9943 11898 -9891
rect 11842 -9945 11898 -9943
rect 11923 -9891 11979 -9889
rect 11923 -9943 11925 -9891
rect 11925 -9943 11977 -9891
rect 11977 -9943 11979 -9891
rect 11923 -9945 11979 -9943
rect 12005 -9891 12061 -9889
rect 12005 -9943 12007 -9891
rect 12007 -9943 12059 -9891
rect 12059 -9943 12061 -9891
rect 12005 -9945 12061 -9943
rect 12086 -9891 12142 -9889
rect 12086 -9943 12088 -9891
rect 12088 -9943 12140 -9891
rect 12140 -9943 12142 -9891
rect 12086 -9945 12142 -9943
rect 12167 -9891 12223 -9889
rect 12167 -9943 12169 -9891
rect 12169 -9943 12221 -9891
rect 12221 -9943 12223 -9891
rect 12167 -9945 12223 -9943
rect 12248 -9891 12304 -9889
rect 12248 -9943 12250 -9891
rect 12250 -9943 12302 -9891
rect 12302 -9943 12304 -9891
rect 12248 -9945 12304 -9943
rect 12329 -9891 12385 -9889
rect 12329 -9943 12331 -9891
rect 12331 -9943 12383 -9891
rect 12383 -9943 12385 -9891
rect 12329 -9945 12385 -9943
rect 12410 -9891 12466 -9889
rect 12410 -9943 12412 -9891
rect 12412 -9943 12464 -9891
rect 12464 -9943 12466 -9891
rect 12410 -9945 12466 -9943
rect 12491 -9891 12547 -9889
rect 12491 -9943 12493 -9891
rect 12493 -9943 12545 -9891
rect 12545 -9943 12547 -9891
rect 12491 -9945 12547 -9943
rect 12573 -9891 12629 -9889
rect 12573 -9943 12575 -9891
rect 12575 -9943 12627 -9891
rect 12627 -9943 12629 -9891
rect 12573 -9945 12629 -9943
rect 12654 -9891 12710 -9889
rect 12654 -9943 12656 -9891
rect 12656 -9943 12708 -9891
rect 12708 -9943 12710 -9891
rect 12654 -9945 12710 -9943
rect 12735 -9891 12791 -9889
rect 12735 -9943 12737 -9891
rect 12737 -9943 12789 -9891
rect 12789 -9943 12791 -9891
rect 12735 -9945 12791 -9943
rect 12816 -9891 12872 -9889
rect 12816 -9943 12818 -9891
rect 12818 -9943 12870 -9891
rect 12870 -9943 12872 -9891
rect 12816 -9945 12872 -9943
rect 12897 -9891 12953 -9889
rect 12897 -9943 12899 -9891
rect 12899 -9943 12951 -9891
rect 12951 -9943 12953 -9891
rect 12897 -9945 12953 -9943
rect 12978 -9891 13034 -9889
rect 12978 -9943 12980 -9891
rect 12980 -9943 13032 -9891
rect 13032 -9943 13034 -9891
rect 12978 -9945 13034 -9943
rect 13059 -9891 13115 -9889
rect 13059 -9943 13061 -9891
rect 13061 -9943 13113 -9891
rect 13113 -9943 13115 -9891
rect 13059 -9945 13115 -9943
rect 13141 -9891 13197 -9889
rect 13141 -9943 13143 -9891
rect 13143 -9943 13195 -9891
rect 13195 -9943 13197 -9891
rect 13141 -9945 13197 -9943
rect 13222 -9891 13278 -9889
rect 13222 -9943 13224 -9891
rect 13224 -9943 13276 -9891
rect 13276 -9943 13278 -9891
rect 13222 -9945 13278 -9943
rect 13303 -9891 13359 -9889
rect 13303 -9943 13305 -9891
rect 13305 -9943 13357 -9891
rect 13357 -9943 13359 -9891
rect 13303 -9945 13359 -9943
rect 13384 -9891 13440 -9889
rect 13384 -9943 13386 -9891
rect 13386 -9943 13438 -9891
rect 13438 -9943 13440 -9891
rect 13384 -9945 13440 -9943
rect 13465 -9891 13521 -9889
rect 13465 -9943 13467 -9891
rect 13467 -9943 13519 -9891
rect 13519 -9943 13521 -9891
rect 13465 -9945 13521 -9943
rect 13546 -9891 13602 -9889
rect 13546 -9943 13548 -9891
rect 13548 -9943 13600 -9891
rect 13600 -9943 13602 -9891
rect 13546 -9945 13602 -9943
rect 13627 -9891 13683 -9889
rect 13627 -9943 13629 -9891
rect 13629 -9943 13681 -9891
rect 13681 -9943 13683 -9891
rect 13627 -9945 13683 -9943
rect 13709 -9891 13765 -9889
rect 13709 -9943 13711 -9891
rect 13711 -9943 13763 -9891
rect 13763 -9943 13765 -9891
rect 13709 -9945 13765 -9943
rect 13790 -9891 13846 -9889
rect 13790 -9943 13792 -9891
rect 13792 -9943 13844 -9891
rect 13844 -9943 13846 -9891
rect 13790 -9945 13846 -9943
rect 13871 -9891 13927 -9889
rect 13871 -9943 13873 -9891
rect 13873 -9943 13925 -9891
rect 13925 -9943 13927 -9891
rect 13871 -9945 13927 -9943
rect 13952 -9891 14008 -9889
rect 13952 -9943 13954 -9891
rect 13954 -9943 14006 -9891
rect 14006 -9943 14008 -9891
rect 13952 -9945 14008 -9943
rect 14033 -9891 14089 -9889
rect 14033 -9943 14035 -9891
rect 14035 -9943 14087 -9891
rect 14087 -9943 14089 -9891
rect 14033 -9945 14089 -9943
rect 14114 -9891 14170 -9889
rect 14114 -9943 14116 -9891
rect 14116 -9943 14168 -9891
rect 14168 -9943 14170 -9891
rect 14114 -9945 14170 -9943
rect 14195 -9891 14251 -9889
rect 14195 -9943 14197 -9891
rect 14197 -9943 14249 -9891
rect 14249 -9943 14251 -9891
rect 14195 -9945 14251 -9943
rect 14277 -9891 14333 -9889
rect 14277 -9943 14279 -9891
rect 14279 -9943 14331 -9891
rect 14331 -9943 14333 -9891
rect 14277 -9945 14333 -9943
rect 14358 -9891 14414 -9889
rect 14358 -9943 14360 -9891
rect 14360 -9943 14412 -9891
rect 14412 -9943 14414 -9891
rect 14358 -9945 14414 -9943
rect 14439 -9891 14495 -9889
rect 14439 -9943 14441 -9891
rect 14441 -9943 14493 -9891
rect 14493 -9943 14495 -9891
rect 14439 -9945 14495 -9943
rect 14520 -9891 14576 -9889
rect 14520 -9943 14522 -9891
rect 14522 -9943 14574 -9891
rect 14574 -9943 14576 -9891
rect 14520 -9945 14576 -9943
rect 14601 -9891 14657 -9889
rect 14601 -9943 14603 -9891
rect 14603 -9943 14655 -9891
rect 14655 -9943 14657 -9891
rect 14601 -9945 14657 -9943
rect 14682 -9891 14738 -9889
rect 14682 -9943 14684 -9891
rect 14684 -9943 14736 -9891
rect 14736 -9943 14738 -9891
rect 14682 -9945 14738 -9943
rect 14763 -9891 14819 -9889
rect 14763 -9943 14765 -9891
rect 14765 -9943 14817 -9891
rect 14817 -9943 14819 -9891
rect 14763 -9945 14819 -9943
rect 14845 -9891 14901 -9889
rect 14845 -9943 14847 -9891
rect 14847 -9943 14899 -9891
rect 14899 -9943 14901 -9891
rect 14845 -9945 14901 -9943
rect 14926 -9891 14982 -9889
rect 14926 -9943 14928 -9891
rect 14928 -9943 14980 -9891
rect 14980 -9943 14982 -9891
rect 14926 -9945 14982 -9943
rect 15007 -9891 15063 -9889
rect 15007 -9943 15009 -9891
rect 15009 -9943 15061 -9891
rect 15061 -9943 15063 -9891
rect 15007 -9945 15063 -9943
rect 15088 -9891 15144 -9889
rect 15088 -9943 15090 -9891
rect 15090 -9943 15142 -9891
rect 15142 -9943 15144 -9891
rect 15088 -9945 15144 -9943
rect 15169 -9891 15225 -9889
rect 15169 -9943 15171 -9891
rect 15171 -9943 15223 -9891
rect 15223 -9943 15225 -9891
rect 15169 -9945 15225 -9943
rect 15250 -9891 15306 -9889
rect 15250 -9943 15252 -9891
rect 15252 -9943 15304 -9891
rect 15304 -9943 15306 -9891
rect 15250 -9945 15306 -9943
rect 15331 -9891 15387 -9889
rect 15331 -9943 15333 -9891
rect 15333 -9943 15385 -9891
rect 15385 -9943 15387 -9891
rect 15331 -9945 15387 -9943
rect 15413 -9891 15469 -9889
rect 15413 -9943 15415 -9891
rect 15415 -9943 15467 -9891
rect 15467 -9943 15469 -9891
rect 15413 -9945 15469 -9943
rect 15494 -9891 15550 -9889
rect 15494 -9943 15496 -9891
rect 15496 -9943 15548 -9891
rect 15548 -9943 15550 -9891
rect 15494 -9945 15550 -9943
rect 15575 -9891 15631 -9889
rect 15575 -9943 15577 -9891
rect 15577 -9943 15629 -9891
rect 15629 -9943 15631 -9891
rect 15575 -9945 15631 -9943
rect 15656 -9891 15712 -9889
rect 15656 -9943 15658 -9891
rect 15658 -9943 15710 -9891
rect 15710 -9943 15712 -9891
rect 15656 -9945 15712 -9943
rect 15737 -9891 15793 -9889
rect 15737 -9943 15739 -9891
rect 15739 -9943 15791 -9891
rect 15791 -9943 15793 -9891
rect 15737 -9945 15793 -9943
rect 15818 -9891 15874 -9889
rect 15818 -9943 15820 -9891
rect 15820 -9943 15872 -9891
rect 15872 -9943 15874 -9891
rect 15818 -9945 15874 -9943
rect 15899 -9891 15955 -9889
rect 15899 -9943 15901 -9891
rect 15901 -9943 15953 -9891
rect 15953 -9943 15955 -9891
rect 15899 -9945 15955 -9943
rect 15981 -9891 16037 -9889
rect 15981 -9943 15983 -9891
rect 15983 -9943 16035 -9891
rect 16035 -9943 16037 -9891
rect 15981 -9945 16037 -9943
rect 16062 -9891 16118 -9889
rect 16062 -9943 16064 -9891
rect 16064 -9943 16116 -9891
rect 16116 -9943 16118 -9891
rect 16062 -9945 16118 -9943
rect 16143 -9891 16199 -9889
rect 16143 -9943 16145 -9891
rect 16145 -9943 16197 -9891
rect 16197 -9943 16199 -9891
rect 16143 -9945 16199 -9943
rect 16224 -9891 16280 -9889
rect 16224 -9943 16226 -9891
rect 16226 -9943 16278 -9891
rect 16278 -9943 16280 -9891
rect 16224 -9945 16280 -9943
rect 16305 -9891 16361 -9889
rect 16305 -9943 16307 -9891
rect 16307 -9943 16359 -9891
rect 16359 -9943 16361 -9891
rect 16305 -9945 16361 -9943
rect 16386 -9891 16442 -9889
rect 16386 -9943 16388 -9891
rect 16388 -9943 16440 -9891
rect 16440 -9943 16442 -9891
rect 16386 -9945 16442 -9943
rect 16467 -9891 16523 -9889
rect 16467 -9943 16469 -9891
rect 16469 -9943 16521 -9891
rect 16521 -9943 16523 -9891
rect 16467 -9945 16523 -9943
rect 16549 -9891 16605 -9889
rect 16549 -9943 16551 -9891
rect 16551 -9943 16603 -9891
rect 16603 -9943 16605 -9891
rect 16549 -9945 16605 -9943
rect 16630 -9891 16686 -9889
rect 16630 -9943 16632 -9891
rect 16632 -9943 16684 -9891
rect 16684 -9943 16686 -9891
rect 16630 -9945 16686 -9943
rect 16711 -9891 16767 -9889
rect 16711 -9943 16713 -9891
rect 16713 -9943 16765 -9891
rect 16765 -9943 16767 -9891
rect 16711 -9945 16767 -9943
rect 16792 -9891 16848 -9889
rect 16792 -9943 16794 -9891
rect 16794 -9943 16846 -9891
rect 16846 -9943 16848 -9891
rect 16792 -9945 16848 -9943
rect 16873 -9891 16929 -9889
rect 16873 -9943 16875 -9891
rect 16875 -9943 16927 -9891
rect 16927 -9943 16929 -9891
rect 16873 -9945 16929 -9943
rect 16954 -9891 17010 -9889
rect 16954 -9943 16956 -9891
rect 16956 -9943 17008 -9891
rect 17008 -9943 17010 -9891
rect 16954 -9945 17010 -9943
rect 17035 -9891 17091 -9889
rect 17035 -9943 17037 -9891
rect 17037 -9943 17089 -9891
rect 17089 -9943 17091 -9891
rect 17035 -9945 17091 -9943
rect 17117 -9891 17173 -9889
rect 17117 -9943 17119 -9891
rect 17119 -9943 17171 -9891
rect 17171 -9943 17173 -9891
rect 17117 -9945 17173 -9943
rect 17198 -9891 17254 -9889
rect 17198 -9943 17200 -9891
rect 17200 -9943 17252 -9891
rect 17252 -9943 17254 -9891
rect 17198 -9945 17254 -9943
rect 17279 -9891 17335 -9889
rect 17279 -9943 17281 -9891
rect 17281 -9943 17333 -9891
rect 17333 -9943 17335 -9891
rect 17279 -9945 17335 -9943
rect 17360 -9891 17416 -9889
rect 17360 -9943 17362 -9891
rect 17362 -9943 17414 -9891
rect 17414 -9943 17416 -9891
rect 17360 -9945 17416 -9943
rect 17441 -9891 17497 -9889
rect 17441 -9943 17443 -9891
rect 17443 -9943 17495 -9891
rect 17495 -9943 17497 -9891
rect 17441 -9945 17497 -9943
rect 17522 -9891 17578 -9889
rect 17522 -9943 17524 -9891
rect 17524 -9943 17576 -9891
rect 17576 -9943 17578 -9891
rect 17522 -9945 17578 -9943
rect 17603 -9891 17659 -9889
rect 17603 -9943 17605 -9891
rect 17605 -9943 17657 -9891
rect 17657 -9943 17659 -9891
rect 17603 -9945 17659 -9943
rect 17684 -9891 17740 -9889
rect 17684 -9943 17686 -9891
rect 17686 -9943 17738 -9891
rect 17738 -9943 17740 -9891
rect 17684 -9945 17740 -9943
rect 17765 -9891 17821 -9889
rect 17765 -9943 17767 -9891
rect 17767 -9943 17819 -9891
rect 17819 -9943 17821 -9891
rect 17765 -9945 17821 -9943
rect 17846 -9891 17902 -9889
rect 17846 -9943 17848 -9891
rect 17848 -9943 17900 -9891
rect 17900 -9943 17902 -9891
rect 17846 -9945 17902 -9943
rect 17927 -9891 17983 -9889
rect 17927 -9943 17929 -9891
rect 17929 -9943 17981 -9891
rect 17981 -9943 17983 -9891
rect 17927 -9945 17983 -9943
rect 18008 -9891 18064 -9889
rect 18008 -9943 18010 -9891
rect 18010 -9943 18062 -9891
rect 18062 -9943 18064 -9891
rect 18008 -9945 18064 -9943
rect 18089 -9891 18145 -9889
rect 18089 -9943 18091 -9891
rect 18091 -9943 18143 -9891
rect 18143 -9943 18145 -9891
rect 18089 -9945 18145 -9943
rect 18171 -9891 18227 -9889
rect 18171 -9943 18173 -9891
rect 18173 -9943 18225 -9891
rect 18225 -9943 18227 -9891
rect 18171 -9945 18227 -9943
rect 18252 -9891 18308 -9889
rect 18252 -9943 18254 -9891
rect 18254 -9943 18306 -9891
rect 18306 -9943 18308 -9891
rect 18252 -9945 18308 -9943
rect 18333 -9891 18389 -9889
rect 18333 -9943 18335 -9891
rect 18335 -9943 18387 -9891
rect 18387 -9943 18389 -9891
rect 18333 -9945 18389 -9943
rect 18414 -9891 18470 -9889
rect 18414 -9943 18416 -9891
rect 18416 -9943 18468 -9891
rect 18468 -9943 18470 -9891
rect 18414 -9945 18470 -9943
rect 18495 -9891 18551 -9889
rect 18495 -9943 18497 -9891
rect 18497 -9943 18549 -9891
rect 18549 -9943 18551 -9891
rect 18495 -9945 18551 -9943
rect 18576 -9891 18632 -9889
rect 18576 -9943 18578 -9891
rect 18578 -9943 18630 -9891
rect 18630 -9943 18632 -9891
rect 18576 -9945 18632 -9943
rect 18657 -9891 18713 -9889
rect 18657 -9943 18659 -9891
rect 18659 -9943 18711 -9891
rect 18711 -9943 18713 -9891
rect 18657 -9945 18713 -9943
rect 18739 -9891 18795 -9889
rect 18739 -9943 18741 -9891
rect 18741 -9943 18793 -9891
rect 18793 -9943 18795 -9891
rect 18739 -9945 18795 -9943
rect 18820 -9891 18876 -9889
rect 18820 -9943 18822 -9891
rect 18822 -9943 18874 -9891
rect 18874 -9943 18876 -9891
rect 18820 -9945 18876 -9943
rect 18901 -9891 18957 -9889
rect 18901 -9943 18903 -9891
rect 18903 -9943 18955 -9891
rect 18955 -9943 18957 -9891
rect 18901 -9945 18957 -9943
rect 18982 -9891 19038 -9889
rect 18982 -9943 18984 -9891
rect 18984 -9943 19036 -9891
rect 19036 -9943 19038 -9891
rect 18982 -9945 19038 -9943
rect 19063 -9891 19119 -9889
rect 19063 -9943 19065 -9891
rect 19065 -9943 19117 -9891
rect 19117 -9943 19119 -9891
rect 19063 -9945 19119 -9943
rect 19144 -9891 19200 -9889
rect 19144 -9943 19146 -9891
rect 19146 -9943 19198 -9891
rect 19198 -9943 19200 -9891
rect 19144 -9945 19200 -9943
rect 19225 -9891 19281 -9889
rect 19225 -9943 19227 -9891
rect 19227 -9943 19279 -9891
rect 19279 -9943 19281 -9891
rect 19225 -9945 19281 -9943
rect 19307 -9891 19363 -9889
rect 19307 -9943 19309 -9891
rect 19309 -9943 19361 -9891
rect 19361 -9943 19363 -9891
rect 19307 -9945 19363 -9943
rect 19388 -9891 19444 -9889
rect 19388 -9943 19390 -9891
rect 19390 -9943 19442 -9891
rect 19442 -9943 19444 -9891
rect 19388 -9945 19444 -9943
rect 19469 -9891 19525 -9889
rect 19469 -9943 19471 -9891
rect 19471 -9943 19523 -9891
rect 19523 -9943 19525 -9891
rect 19469 -9945 19525 -9943
rect 19550 -9891 19606 -9889
rect 19550 -9943 19552 -9891
rect 19552 -9943 19604 -9891
rect 19604 -9943 19606 -9891
rect 19550 -9945 19606 -9943
rect 19631 -9891 19687 -9889
rect 19631 -9943 19633 -9891
rect 19633 -9943 19685 -9891
rect 19685 -9943 19687 -9891
rect 19631 -9945 19687 -9943
rect 19712 -9891 19768 -9889
rect 19712 -9943 19714 -9891
rect 19714 -9943 19766 -9891
rect 19766 -9943 19768 -9891
rect 19712 -9945 19768 -9943
rect 19793 -9891 19849 -9889
rect 19793 -9943 19795 -9891
rect 19795 -9943 19847 -9891
rect 19847 -9943 19849 -9891
rect 19793 -9945 19849 -9943
rect 19875 -9891 19931 -9889
rect 19875 -9943 19877 -9891
rect 19877 -9943 19929 -9891
rect 19929 -9943 19931 -9891
rect 19875 -9945 19931 -9943
rect 19956 -9891 20012 -9889
rect 19956 -9943 19958 -9891
rect 19958 -9943 20010 -9891
rect 20010 -9943 20012 -9891
rect 19956 -9945 20012 -9943
rect 20037 -9891 20093 -9889
rect 20037 -9943 20039 -9891
rect 20039 -9943 20091 -9891
rect 20091 -9943 20093 -9891
rect 20037 -9945 20093 -9943
rect 20118 -9891 20174 -9889
rect 20118 -9943 20120 -9891
rect 20120 -9943 20172 -9891
rect 20172 -9943 20174 -9891
rect 20118 -9945 20174 -9943
rect 20199 -9891 20255 -9889
rect 20199 -9943 20201 -9891
rect 20201 -9943 20253 -9891
rect 20253 -9943 20255 -9891
rect 20199 -9945 20255 -9943
rect 20280 -9891 20336 -9889
rect 20280 -9943 20282 -9891
rect 20282 -9943 20334 -9891
rect 20334 -9943 20336 -9891
rect 20280 -9945 20336 -9943
rect 20361 -9891 20417 -9889
rect 20361 -9943 20363 -9891
rect 20363 -9943 20415 -9891
rect 20415 -9943 20417 -9891
rect 20361 -9945 20417 -9943
rect 20443 -9891 20499 -9889
rect 20443 -9943 20445 -9891
rect 20445 -9943 20497 -9891
rect 20497 -9943 20499 -9891
rect 20443 -9945 20499 -9943
rect 20524 -9891 20580 -9889
rect 20524 -9943 20526 -9891
rect 20526 -9943 20578 -9891
rect 20578 -9943 20580 -9891
rect 20524 -9945 20580 -9943
rect 20605 -9891 20661 -9889
rect 20605 -9943 20607 -9891
rect 20607 -9943 20659 -9891
rect 20659 -9943 20661 -9891
rect 20605 -9945 20661 -9943
rect 20686 -9891 20742 -9889
rect 20686 -9943 20688 -9891
rect 20688 -9943 20740 -9891
rect 20740 -9943 20742 -9891
rect 20686 -9945 20742 -9943
rect 20767 -9891 20823 -9889
rect 20767 -9943 20769 -9891
rect 20769 -9943 20821 -9891
rect 20821 -9943 20823 -9891
rect 20767 -9945 20823 -9943
rect 20848 -9891 20904 -9889
rect 20848 -9943 20850 -9891
rect 20850 -9943 20902 -9891
rect 20902 -9943 20904 -9891
rect 20848 -9945 20904 -9943
rect 20929 -9891 20985 -9889
rect 20929 -9943 20931 -9891
rect 20931 -9943 20983 -9891
rect 20983 -9943 20985 -9891
rect 20929 -9945 20985 -9943
rect 21011 -9891 21067 -9889
rect 21011 -9943 21013 -9891
rect 21013 -9943 21065 -9891
rect 21065 -9943 21067 -9891
rect 21011 -9945 21067 -9943
rect 21092 -9891 21148 -9889
rect 21092 -9943 21094 -9891
rect 21094 -9943 21146 -9891
rect 21146 -9943 21148 -9891
rect 21092 -9945 21148 -9943
rect 21173 -9891 21229 -9889
rect 21173 -9943 21175 -9891
rect 21175 -9943 21227 -9891
rect 21227 -9943 21229 -9891
rect 21173 -9945 21229 -9943
rect 21254 -9891 21310 -9889
rect 21254 -9943 21256 -9891
rect 21256 -9943 21308 -9891
rect 21308 -9943 21310 -9891
rect 21254 -9945 21310 -9943
rect 21335 -9891 21391 -9889
rect 21335 -9943 21337 -9891
rect 21337 -9943 21389 -9891
rect 21389 -9943 21391 -9891
rect 21335 -9945 21391 -9943
rect 21416 -9891 21472 -9889
rect 21416 -9943 21418 -9891
rect 21418 -9943 21470 -9891
rect 21470 -9943 21472 -9891
rect 21416 -9945 21472 -9943
rect 21497 -9891 21553 -9889
rect 21497 -9943 21499 -9891
rect 21499 -9943 21551 -9891
rect 21551 -9943 21553 -9891
rect 21497 -9945 21553 -9943
rect 21579 -9891 21635 -9889
rect 21579 -9943 21581 -9891
rect 21581 -9943 21633 -9891
rect 21633 -9943 21635 -9891
rect 21579 -9945 21635 -9943
rect 21660 -9891 21716 -9889
rect 21660 -9943 21662 -9891
rect 21662 -9943 21714 -9891
rect 21714 -9943 21716 -9891
rect 21660 -9945 21716 -9943
rect 21741 -9891 21797 -9889
rect 21741 -9943 21743 -9891
rect 21743 -9943 21795 -9891
rect 21795 -9943 21797 -9891
rect 21741 -9945 21797 -9943
rect 21822 -9891 21878 -9889
rect 21822 -9943 21824 -9891
rect 21824 -9943 21876 -9891
rect 21876 -9943 21878 -9891
rect 21822 -9945 21878 -9943
rect 21903 -9891 21959 -9889
rect 21903 -9943 21905 -9891
rect 21905 -9943 21957 -9891
rect 21957 -9943 21959 -9891
rect 21903 -9945 21959 -9943
rect 21984 -9891 22040 -9889
rect 21984 -9943 21986 -9891
rect 21986 -9943 22038 -9891
rect 22038 -9943 22040 -9891
rect 21984 -9945 22040 -9943
rect 22065 -9891 22121 -9889
rect 22065 -9943 22067 -9891
rect 22067 -9943 22119 -9891
rect 22119 -9943 22121 -9891
rect 22065 -9945 22121 -9943
rect 22147 -9891 22203 -9889
rect 22147 -9943 22149 -9891
rect 22149 -9943 22201 -9891
rect 22201 -9943 22203 -9891
rect 22147 -9945 22203 -9943
rect 22228 -9891 22284 -9889
rect 22228 -9943 22230 -9891
rect 22230 -9943 22282 -9891
rect 22282 -9943 22284 -9891
rect 22228 -9945 22284 -9943
rect 22309 -9891 22365 -9889
rect 22309 -9943 22311 -9891
rect 22311 -9943 22363 -9891
rect 22363 -9943 22365 -9891
rect 22309 -9945 22365 -9943
rect 22390 -9891 22446 -9889
rect 22390 -9943 22392 -9891
rect 22392 -9943 22444 -9891
rect 22444 -9943 22446 -9891
rect 22390 -9945 22446 -9943
rect 22471 -9891 22527 -9889
rect 22471 -9943 22473 -9891
rect 22473 -9943 22525 -9891
rect 22525 -9943 22527 -9891
rect 22471 -9945 22527 -9943
rect 22552 -9891 22608 -9889
rect 22552 -9943 22554 -9891
rect 22554 -9943 22606 -9891
rect 22606 -9943 22608 -9891
rect 22552 -9945 22608 -9943
rect 22633 -9891 22689 -9889
rect 22633 -9943 22635 -9891
rect 22635 -9943 22687 -9891
rect 22687 -9943 22689 -9891
rect 22633 -9945 22689 -9943
rect 22715 -9891 22771 -9889
rect 22715 -9943 22717 -9891
rect 22717 -9943 22769 -9891
rect 22769 -9943 22771 -9891
rect 22715 -9945 22771 -9943
rect 22796 -9891 22852 -9889
rect 22796 -9943 22798 -9891
rect 22798 -9943 22850 -9891
rect 22850 -9943 22852 -9891
rect 22796 -9945 22852 -9943
rect 22877 -9891 22933 -9889
rect 22877 -9943 22879 -9891
rect 22879 -9943 22931 -9891
rect 22931 -9943 22933 -9891
rect 22877 -9945 22933 -9943
rect 22958 -9891 23014 -9889
rect 22958 -9943 22960 -9891
rect 22960 -9943 23012 -9891
rect 23012 -9943 23014 -9891
rect 22958 -9945 23014 -9943
rect 23039 -9891 23095 -9889
rect 23039 -9943 23041 -9891
rect 23041 -9943 23093 -9891
rect 23093 -9943 23095 -9891
rect 23039 -9945 23095 -9943
rect 23120 -9891 23176 -9889
rect 23120 -9943 23122 -9891
rect 23122 -9943 23174 -9891
rect 23174 -9943 23176 -9891
rect 23120 -9945 23176 -9943
rect 23201 -9891 23257 -9889
rect 23201 -9943 23203 -9891
rect 23203 -9943 23255 -9891
rect 23255 -9943 23257 -9891
rect 23201 -9945 23257 -9943
rect 23283 -9891 23339 -9889
rect 23283 -9943 23285 -9891
rect 23285 -9943 23337 -9891
rect 23337 -9943 23339 -9891
rect 23283 -9945 23339 -9943
rect 23364 -9891 23420 -9889
rect 23364 -9943 23366 -9891
rect 23366 -9943 23418 -9891
rect 23418 -9943 23420 -9891
rect 23364 -9945 23420 -9943
rect 23445 -9891 23501 -9889
rect 23445 -9943 23447 -9891
rect 23447 -9943 23499 -9891
rect 23499 -9943 23501 -9891
rect 23445 -9945 23501 -9943
rect 23526 -9891 23582 -9889
rect 23526 -9943 23528 -9891
rect 23528 -9943 23580 -9891
rect 23580 -9943 23582 -9891
rect 23526 -9945 23582 -9943
rect 23607 -9891 23663 -9889
rect 23607 -9943 23609 -9891
rect 23609 -9943 23661 -9891
rect 23661 -9943 23663 -9891
rect 23607 -9945 23663 -9943
rect 23688 -9891 23744 -9889
rect 23688 -9943 23690 -9891
rect 23690 -9943 23742 -9891
rect 23742 -9943 23744 -9891
rect 23688 -9945 23744 -9943
rect 23769 -9891 23825 -9889
rect 23769 -9943 23771 -9891
rect 23771 -9943 23823 -9891
rect 23823 -9943 23825 -9891
rect 23769 -9945 23825 -9943
rect 23851 -9891 23907 -9889
rect 23851 -9943 23853 -9891
rect 23853 -9943 23905 -9891
rect 23905 -9943 23907 -9891
rect 23851 -9945 23907 -9943
rect 23932 -9891 23988 -9889
rect 23932 -9943 23934 -9891
rect 23934 -9943 23986 -9891
rect 23986 -9943 23988 -9891
rect 23932 -9945 23988 -9943
rect 24013 -9891 24069 -9889
rect 24013 -9943 24015 -9891
rect 24015 -9943 24067 -9891
rect 24067 -9943 24069 -9891
rect 24013 -9945 24069 -9943
rect 24094 -9891 24150 -9889
rect 24094 -9943 24096 -9891
rect 24096 -9943 24148 -9891
rect 24148 -9943 24150 -9891
rect 24094 -9945 24150 -9943
rect 24175 -9891 24231 -9889
rect 24175 -9943 24177 -9891
rect 24177 -9943 24229 -9891
rect 24229 -9943 24231 -9891
rect 24175 -9945 24231 -9943
rect 24256 -9891 24312 -9889
rect 24256 -9943 24258 -9891
rect 24258 -9943 24310 -9891
rect 24310 -9943 24312 -9891
rect 24256 -9945 24312 -9943
rect 24337 -9891 24393 -9889
rect 24337 -9943 24339 -9891
rect 24339 -9943 24391 -9891
rect 24391 -9943 24393 -9891
rect 24337 -9945 24393 -9943
rect 24419 -9891 24475 -9889
rect 24419 -9943 24421 -9891
rect 24421 -9943 24473 -9891
rect 24473 -9943 24475 -9891
rect 24419 -9945 24475 -9943
rect 24500 -9891 24556 -9889
rect 24500 -9943 24502 -9891
rect 24502 -9943 24554 -9891
rect 24554 -9943 24556 -9891
rect 24500 -9945 24556 -9943
rect 24581 -9891 24637 -9889
rect 24581 -9943 24583 -9891
rect 24583 -9943 24635 -9891
rect 24635 -9943 24637 -9891
rect 24581 -9945 24637 -9943
rect 24662 -9891 24718 -9889
rect 24662 -9943 24664 -9891
rect 24664 -9943 24716 -9891
rect 24716 -9943 24718 -9891
rect 24662 -9945 24718 -9943
rect 24743 -9891 24799 -9889
rect 24743 -9943 24745 -9891
rect 24745 -9943 24797 -9891
rect 24797 -9943 24799 -9891
rect 24743 -9945 24799 -9943
rect 24824 -9891 24880 -9889
rect 24824 -9943 24826 -9891
rect 24826 -9943 24878 -9891
rect 24878 -9943 24880 -9891
rect 24824 -9945 24880 -9943
rect 24905 -9891 24961 -9889
rect 24905 -9943 24907 -9891
rect 24907 -9943 24959 -9891
rect 24959 -9943 24961 -9891
rect 24905 -9945 24961 -9943
rect 24987 -9891 25043 -9889
rect 24987 -9943 24989 -9891
rect 24989 -9943 25041 -9891
rect 25041 -9943 25043 -9891
rect 24987 -9945 25043 -9943
rect 25068 -9891 25124 -9889
rect 25068 -9943 25070 -9891
rect 25070 -9943 25122 -9891
rect 25122 -9943 25124 -9891
rect 25068 -9945 25124 -9943
rect 25149 -9891 25205 -9889
rect 25149 -9943 25151 -9891
rect 25151 -9943 25203 -9891
rect 25203 -9943 25205 -9891
rect 25149 -9945 25205 -9943
rect 25230 -9891 25286 -9889
rect 25230 -9943 25232 -9891
rect 25232 -9943 25284 -9891
rect 25284 -9943 25286 -9891
rect 25230 -9945 25286 -9943
rect 25311 -9891 25367 -9889
rect 25311 -9943 25313 -9891
rect 25313 -9943 25365 -9891
rect 25365 -9943 25367 -9891
rect 25311 -9945 25367 -9943
rect 25392 -9891 25448 -9889
rect 25392 -9943 25394 -9891
rect 25394 -9943 25446 -9891
rect 25446 -9943 25448 -9891
rect 25392 -9945 25448 -9943
rect 25473 -9891 25529 -9889
rect 25473 -9943 25475 -9891
rect 25475 -9943 25527 -9891
rect 25527 -9943 25529 -9891
rect 25473 -9945 25529 -9943
rect 25555 -9891 25611 -9889
rect 25555 -9943 25557 -9891
rect 25557 -9943 25609 -9891
rect 25609 -9943 25611 -9891
rect 25555 -9945 25611 -9943
rect 25636 -9891 25692 -9889
rect 25636 -9943 25638 -9891
rect 25638 -9943 25690 -9891
rect 25690 -9943 25692 -9891
rect 25636 -9945 25692 -9943
rect 25717 -9891 25773 -9889
rect 25717 -9943 25719 -9891
rect 25719 -9943 25771 -9891
rect 25771 -9943 25773 -9891
rect 25717 -9945 25773 -9943
rect 25798 -9891 25854 -9889
rect 25798 -9943 25800 -9891
rect 25800 -9943 25852 -9891
rect 25852 -9943 25854 -9891
rect 25798 -9945 25854 -9943
rect 25879 -9891 25935 -9889
rect 25879 -9943 25881 -9891
rect 25881 -9943 25933 -9891
rect 25933 -9943 25935 -9891
rect 25879 -9945 25935 -9943
rect 25960 -9891 26016 -9889
rect 25960 -9943 25962 -9891
rect 25962 -9943 26014 -9891
rect 26014 -9943 26016 -9891
rect 25960 -9945 26016 -9943
rect 26041 -9891 26097 -9889
rect 26041 -9943 26043 -9891
rect 26043 -9943 26095 -9891
rect 26095 -9943 26097 -9891
rect 26041 -9945 26097 -9943
rect 26123 -9891 26179 -9889
rect 26123 -9943 26125 -9891
rect 26125 -9943 26177 -9891
rect 26177 -9943 26179 -9891
rect 26123 -9945 26179 -9943
rect 26204 -9891 26260 -9889
rect 26204 -9943 26206 -9891
rect 26206 -9943 26258 -9891
rect 26258 -9943 26260 -9891
rect 26204 -9945 26260 -9943
<< metal3 >>
rect 3012 3181 11174 3182
rect 11515 3181 24739 3182
rect 3012 3174 24739 3181
rect 3012 3118 3036 3174
rect 3092 3118 3118 3174
rect 3174 3118 3199 3174
rect 3255 3118 3280 3174
rect 3336 3118 3361 3174
rect 3417 3118 3442 3174
rect 3498 3118 3523 3174
rect 3579 3118 3604 3174
rect 3660 3118 3686 3174
rect 3742 3118 3767 3174
rect 3823 3118 3848 3174
rect 3904 3118 3929 3174
rect 3985 3118 4010 3174
rect 4066 3118 4091 3174
rect 4147 3118 4172 3174
rect 4228 3118 4254 3174
rect 4310 3118 4335 3174
rect 4391 3118 4416 3174
rect 4472 3118 4497 3174
rect 4553 3118 4578 3174
rect 4634 3118 4659 3174
rect 4715 3118 4740 3174
rect 4796 3118 4822 3174
rect 4878 3118 4903 3174
rect 4959 3118 4984 3174
rect 5040 3118 5065 3174
rect 5121 3118 5146 3174
rect 5202 3118 5227 3174
rect 5283 3118 5308 3174
rect 5364 3118 5390 3174
rect 5446 3118 5471 3174
rect 5527 3118 5552 3174
rect 5608 3118 5633 3174
rect 5689 3118 5714 3174
rect 5770 3118 5795 3174
rect 5851 3118 5876 3174
rect 5932 3118 5958 3174
rect 6014 3118 6039 3174
rect 6095 3118 6120 3174
rect 6176 3118 6201 3174
rect 6257 3118 6282 3174
rect 6338 3118 6363 3174
rect 6419 3118 6444 3174
rect 6500 3118 6526 3174
rect 6582 3118 6607 3174
rect 6663 3118 6688 3174
rect 6744 3118 6769 3174
rect 6825 3118 6850 3174
rect 6906 3118 6931 3174
rect 6987 3118 7012 3174
rect 7068 3118 7094 3174
rect 7150 3118 7175 3174
rect 7231 3118 7256 3174
rect 7312 3118 7337 3174
rect 7393 3118 7418 3174
rect 7474 3118 7499 3174
rect 7555 3118 7580 3174
rect 7636 3118 7662 3174
rect 7718 3118 7743 3174
rect 7799 3118 7824 3174
rect 7880 3118 7905 3174
rect 7961 3118 7986 3174
rect 8042 3118 8067 3174
rect 8123 3118 8148 3174
rect 8204 3118 8230 3174
rect 8286 3118 8311 3174
rect 8367 3118 8392 3174
rect 8448 3118 8473 3174
rect 8529 3118 8554 3174
rect 8610 3118 8635 3174
rect 8691 3118 8716 3174
rect 8772 3118 8798 3174
rect 8854 3118 8879 3174
rect 8935 3118 8960 3174
rect 9016 3118 9041 3174
rect 9097 3118 9122 3174
rect 9178 3118 9203 3174
rect 9259 3118 9284 3174
rect 9340 3118 9366 3174
rect 9422 3118 9447 3174
rect 9503 3118 9528 3174
rect 9584 3118 9609 3174
rect 9665 3118 9690 3174
rect 9746 3118 9771 3174
rect 9827 3118 9852 3174
rect 9908 3118 9934 3174
rect 9990 3118 10015 3174
rect 10071 3118 10096 3174
rect 10152 3118 10177 3174
rect 10233 3118 10258 3174
rect 10314 3118 10339 3174
rect 10395 3118 10420 3174
rect 10476 3118 10502 3174
rect 10558 3118 10583 3174
rect 10639 3118 10664 3174
rect 10720 3118 10745 3174
rect 10801 3118 10826 3174
rect 10882 3118 10907 3174
rect 10963 3118 10988 3174
rect 11044 3118 11116 3174
rect 11172 3118 11197 3174
rect 11253 3118 11278 3174
rect 11334 3118 11359 3174
rect 11415 3118 11440 3174
rect 11496 3118 11521 3174
rect 11577 3118 11602 3174
rect 11658 3118 11684 3174
rect 11740 3118 11765 3174
rect 11821 3118 11846 3174
rect 11902 3118 11927 3174
rect 11983 3118 12008 3174
rect 12064 3118 12089 3174
rect 12145 3118 12170 3174
rect 12226 3118 12252 3174
rect 12308 3118 12333 3174
rect 12389 3118 12414 3174
rect 12470 3118 12495 3174
rect 12551 3118 12576 3174
rect 12632 3118 12657 3174
rect 12713 3118 12738 3174
rect 12794 3118 12820 3174
rect 12876 3118 12901 3174
rect 12957 3118 12982 3174
rect 13038 3118 13063 3174
rect 13119 3118 13144 3174
rect 13200 3118 13225 3174
rect 13281 3118 13306 3174
rect 13362 3118 13388 3174
rect 13444 3118 13469 3174
rect 13525 3118 13550 3174
rect 13606 3118 13631 3174
rect 13687 3118 13712 3174
rect 13768 3118 13793 3174
rect 13849 3118 13874 3174
rect 13930 3118 13956 3174
rect 14012 3118 14037 3174
rect 14093 3118 14118 3174
rect 14174 3118 14199 3174
rect 14255 3118 14280 3174
rect 14336 3118 14361 3174
rect 14417 3118 14442 3174
rect 14498 3118 14524 3174
rect 14580 3118 14605 3174
rect 14661 3118 14686 3174
rect 14742 3118 14767 3174
rect 14823 3118 14848 3174
rect 14904 3118 14929 3174
rect 14985 3118 15010 3174
rect 15066 3118 15092 3174
rect 15148 3118 15173 3174
rect 15229 3118 15254 3174
rect 15310 3118 15335 3174
rect 15391 3118 15416 3174
rect 15472 3118 15497 3174
rect 15553 3118 15578 3174
rect 15634 3118 15660 3174
rect 15716 3118 15741 3174
rect 15797 3118 15822 3174
rect 15878 3118 15903 3174
rect 15959 3118 15984 3174
rect 16040 3118 16065 3174
rect 16121 3118 16146 3174
rect 16202 3118 16228 3174
rect 16284 3118 16309 3174
rect 16365 3118 16390 3174
rect 16446 3118 16471 3174
rect 16527 3118 16552 3174
rect 16608 3118 16633 3174
rect 16689 3118 16714 3174
rect 16770 3118 16796 3174
rect 16852 3118 16877 3174
rect 16933 3118 16958 3174
rect 17014 3118 17039 3174
rect 17095 3118 17120 3174
rect 17176 3118 17201 3174
rect 17257 3118 17282 3174
rect 17338 3118 17364 3174
rect 17420 3118 17445 3174
rect 17501 3118 17526 3174
rect 17582 3118 17607 3174
rect 17663 3118 17688 3174
rect 17744 3118 17769 3174
rect 17825 3118 17850 3174
rect 17906 3118 17932 3174
rect 17988 3118 18013 3174
rect 18069 3118 18094 3174
rect 18150 3118 18175 3174
rect 18231 3118 18256 3174
rect 18312 3118 18337 3174
rect 18393 3118 18418 3174
rect 18474 3118 18500 3174
rect 18556 3118 18581 3174
rect 18637 3118 18662 3174
rect 18718 3118 18743 3174
rect 18799 3118 18824 3174
rect 18880 3118 18905 3174
rect 18961 3118 18986 3174
rect 19042 3118 19068 3174
rect 19124 3118 19149 3174
rect 19205 3118 19230 3174
rect 19286 3118 19311 3174
rect 19367 3118 19392 3174
rect 19448 3118 19473 3174
rect 19529 3118 19554 3174
rect 19610 3118 19636 3174
rect 19692 3118 19717 3174
rect 19773 3118 19798 3174
rect 19854 3118 19879 3174
rect 19935 3118 19960 3174
rect 20016 3118 20041 3174
rect 20097 3118 20122 3174
rect 20178 3118 20204 3174
rect 20260 3118 20285 3174
rect 20341 3118 20366 3174
rect 20422 3118 20447 3174
rect 20503 3118 20528 3174
rect 20584 3118 20609 3174
rect 20665 3118 20690 3174
rect 20746 3118 20772 3174
rect 20828 3118 20853 3174
rect 20909 3118 20934 3174
rect 20990 3118 21015 3174
rect 21071 3118 21096 3174
rect 21152 3118 21177 3174
rect 21233 3118 21258 3174
rect 21314 3118 21340 3174
rect 21396 3118 21421 3174
rect 21477 3118 21502 3174
rect 21558 3118 21583 3174
rect 21639 3118 21664 3174
rect 21720 3118 21745 3174
rect 21801 3118 21826 3174
rect 21882 3118 21908 3174
rect 21964 3118 21989 3174
rect 22045 3118 22070 3174
rect 22126 3118 22151 3174
rect 22207 3118 22232 3174
rect 22288 3118 22313 3174
rect 22369 3118 22394 3174
rect 22450 3118 22476 3174
rect 22532 3118 22557 3174
rect 22613 3118 22638 3174
rect 22694 3118 22719 3174
rect 22775 3118 22800 3174
rect 22856 3118 22881 3174
rect 22937 3118 22962 3174
rect 23018 3118 23044 3174
rect 23100 3118 23125 3174
rect 23181 3118 23206 3174
rect 23262 3118 23287 3174
rect 23343 3118 23368 3174
rect 23424 3118 23449 3174
rect 23505 3118 23530 3174
rect 23586 3118 23612 3174
rect 23668 3118 23693 3174
rect 23749 3118 23774 3174
rect 23830 3118 23855 3174
rect 23911 3118 23936 3174
rect 23992 3118 24017 3174
rect 24073 3118 24098 3174
rect 24154 3118 24180 3174
rect 24236 3118 24261 3174
rect 24317 3118 24342 3174
rect 24398 3118 24423 3174
rect 24479 3118 24504 3174
rect 24560 3118 24585 3174
rect 24641 3118 24666 3174
rect 24722 3118 24739 3174
rect 3012 3070 24739 3118
rect 3012 3014 3036 3070
rect 3092 3014 3118 3070
rect 3174 3014 3199 3070
rect 3255 3014 3280 3070
rect 3336 3014 3361 3070
rect 3417 3014 3442 3070
rect 3498 3014 3523 3070
rect 3579 3014 3604 3070
rect 3660 3014 3686 3070
rect 3742 3014 3767 3070
rect 3823 3014 3848 3070
rect 3904 3014 3929 3070
rect 3985 3014 4010 3070
rect 4066 3014 4091 3070
rect 4147 3014 4172 3070
rect 4228 3014 4254 3070
rect 4310 3014 4335 3070
rect 4391 3014 4416 3070
rect 4472 3014 4497 3070
rect 4553 3014 4578 3070
rect 4634 3014 4659 3070
rect 4715 3014 4740 3070
rect 4796 3014 4822 3070
rect 4878 3014 4903 3070
rect 4959 3014 4984 3070
rect 5040 3014 5065 3070
rect 5121 3014 5146 3070
rect 5202 3014 5227 3070
rect 5283 3014 5308 3070
rect 5364 3014 5390 3070
rect 5446 3014 5471 3070
rect 5527 3014 5552 3070
rect 5608 3014 5633 3070
rect 5689 3014 5714 3070
rect 5770 3014 5795 3070
rect 5851 3014 5876 3070
rect 5932 3014 5958 3070
rect 6014 3014 6039 3070
rect 6095 3014 6120 3070
rect 6176 3014 6201 3070
rect 6257 3014 6282 3070
rect 6338 3014 6363 3070
rect 6419 3014 6444 3070
rect 6500 3014 6526 3070
rect 6582 3014 6607 3070
rect 6663 3014 6688 3070
rect 6744 3014 6769 3070
rect 6825 3014 6850 3070
rect 6906 3014 6931 3070
rect 6987 3014 7012 3070
rect 7068 3014 7094 3070
rect 7150 3014 7175 3070
rect 7231 3014 7256 3070
rect 7312 3014 7337 3070
rect 7393 3014 7418 3070
rect 7474 3014 7499 3070
rect 7555 3014 7580 3070
rect 7636 3014 7662 3070
rect 7718 3014 7743 3070
rect 7799 3014 7824 3070
rect 7880 3014 7905 3070
rect 7961 3014 7986 3070
rect 8042 3014 8067 3070
rect 8123 3014 8148 3070
rect 8204 3014 8230 3070
rect 8286 3014 8311 3070
rect 8367 3014 8392 3070
rect 8448 3014 8473 3070
rect 8529 3014 8554 3070
rect 8610 3014 8635 3070
rect 8691 3014 8716 3070
rect 8772 3014 8798 3070
rect 8854 3014 8879 3070
rect 8935 3014 8960 3070
rect 9016 3014 9041 3070
rect 9097 3014 9122 3070
rect 9178 3014 9203 3070
rect 9259 3014 9284 3070
rect 9340 3014 9366 3070
rect 9422 3014 9447 3070
rect 9503 3014 9528 3070
rect 9584 3014 9609 3070
rect 9665 3014 9690 3070
rect 9746 3014 9771 3070
rect 9827 3014 9852 3070
rect 9908 3014 9934 3070
rect 9990 3014 10015 3070
rect 10071 3014 10096 3070
rect 10152 3014 10177 3070
rect 10233 3014 10258 3070
rect 10314 3014 10339 3070
rect 10395 3014 10420 3070
rect 10476 3014 10502 3070
rect 10558 3014 10583 3070
rect 10639 3014 10664 3070
rect 10720 3014 10745 3070
rect 10801 3014 10826 3070
rect 10882 3014 10907 3070
rect 10963 3014 10988 3070
rect 11044 3014 11116 3070
rect 11172 3014 11197 3070
rect 11253 3014 11278 3070
rect 11334 3014 11359 3070
rect 11415 3014 11440 3070
rect 11496 3014 11521 3070
rect 11577 3014 11602 3070
rect 11658 3014 11684 3070
rect 11740 3014 11765 3070
rect 11821 3014 11846 3070
rect 11902 3014 11927 3070
rect 11983 3014 12008 3070
rect 12064 3014 12089 3070
rect 12145 3014 12170 3070
rect 12226 3014 12252 3070
rect 12308 3014 12333 3070
rect 12389 3014 12414 3070
rect 12470 3014 12495 3070
rect 12551 3014 12576 3070
rect 12632 3014 12657 3070
rect 12713 3014 12738 3070
rect 12794 3014 12820 3070
rect 12876 3014 12901 3070
rect 12957 3014 12982 3070
rect 13038 3014 13063 3070
rect 13119 3014 13144 3070
rect 13200 3014 13225 3070
rect 13281 3014 13306 3070
rect 13362 3014 13388 3070
rect 13444 3014 13469 3070
rect 13525 3014 13550 3070
rect 13606 3014 13631 3070
rect 13687 3014 13712 3070
rect 13768 3014 13793 3070
rect 13849 3014 13874 3070
rect 13930 3014 13956 3070
rect 14012 3014 14037 3070
rect 14093 3014 14118 3070
rect 14174 3014 14199 3070
rect 14255 3014 14280 3070
rect 14336 3014 14361 3070
rect 14417 3014 14442 3070
rect 14498 3014 14524 3070
rect 14580 3014 14605 3070
rect 14661 3014 14686 3070
rect 14742 3014 14767 3070
rect 14823 3014 14848 3070
rect 14904 3014 14929 3070
rect 14985 3014 15010 3070
rect 15066 3014 15092 3070
rect 15148 3014 15173 3070
rect 15229 3014 15254 3070
rect 15310 3014 15335 3070
rect 15391 3014 15416 3070
rect 15472 3014 15497 3070
rect 15553 3014 15578 3070
rect 15634 3014 15660 3070
rect 15716 3014 15741 3070
rect 15797 3014 15822 3070
rect 15878 3014 15903 3070
rect 15959 3014 15984 3070
rect 16040 3014 16065 3070
rect 16121 3014 16146 3070
rect 16202 3014 16228 3070
rect 16284 3014 16309 3070
rect 16365 3014 16390 3070
rect 16446 3014 16471 3070
rect 16527 3014 16552 3070
rect 16608 3014 16633 3070
rect 16689 3014 16714 3070
rect 16770 3014 16796 3070
rect 16852 3014 16877 3070
rect 16933 3014 16958 3070
rect 17014 3014 17039 3070
rect 17095 3014 17120 3070
rect 17176 3014 17201 3070
rect 17257 3014 17282 3070
rect 17338 3014 17364 3070
rect 17420 3014 17445 3070
rect 17501 3014 17526 3070
rect 17582 3014 17607 3070
rect 17663 3014 17688 3070
rect 17744 3014 17769 3070
rect 17825 3014 17850 3070
rect 17906 3014 17932 3070
rect 17988 3014 18013 3070
rect 18069 3014 18094 3070
rect 18150 3014 18175 3070
rect 18231 3014 18256 3070
rect 18312 3014 18337 3070
rect 18393 3014 18418 3070
rect 18474 3014 18500 3070
rect 18556 3014 18581 3070
rect 18637 3014 18662 3070
rect 18718 3014 18743 3070
rect 18799 3014 18824 3070
rect 18880 3014 18905 3070
rect 18961 3014 18986 3070
rect 19042 3014 19068 3070
rect 19124 3014 19149 3070
rect 19205 3014 19230 3070
rect 19286 3014 19311 3070
rect 19367 3014 19392 3070
rect 19448 3014 19473 3070
rect 19529 3014 19554 3070
rect 19610 3014 19636 3070
rect 19692 3014 19717 3070
rect 19773 3014 19798 3070
rect 19854 3014 19879 3070
rect 19935 3014 19960 3070
rect 20016 3014 20041 3070
rect 20097 3014 20122 3070
rect 20178 3014 20204 3070
rect 20260 3014 20285 3070
rect 20341 3014 20366 3070
rect 20422 3014 20447 3070
rect 20503 3014 20528 3070
rect 20584 3014 20609 3070
rect 20665 3014 20690 3070
rect 20746 3014 20772 3070
rect 20828 3014 20853 3070
rect 20909 3014 20934 3070
rect 20990 3014 21015 3070
rect 21071 3014 21096 3070
rect 21152 3014 21177 3070
rect 21233 3014 21258 3070
rect 21314 3014 21340 3070
rect 21396 3014 21421 3070
rect 21477 3014 21502 3070
rect 21558 3014 21583 3070
rect 21639 3014 21664 3070
rect 21720 3014 21745 3070
rect 21801 3014 21826 3070
rect 21882 3014 21908 3070
rect 21964 3014 21989 3070
rect 22045 3014 22070 3070
rect 22126 3014 22151 3070
rect 22207 3014 22232 3070
rect 22288 3014 22313 3070
rect 22369 3014 22394 3070
rect 22450 3014 22476 3070
rect 22532 3014 22557 3070
rect 22613 3014 22638 3070
rect 22694 3014 22719 3070
rect 22775 3014 22800 3070
rect 22856 3014 22881 3070
rect 22937 3014 22962 3070
rect 23018 3014 23044 3070
rect 23100 3014 23125 3070
rect 23181 3014 23206 3070
rect 23262 3014 23287 3070
rect 23343 3014 23368 3070
rect 23424 3014 23449 3070
rect 23505 3014 23530 3070
rect 23586 3014 23612 3070
rect 23668 3014 23693 3070
rect 23749 3014 23774 3070
rect 23830 3014 23855 3070
rect 23911 3014 23936 3070
rect 23992 3014 24017 3070
rect 24073 3014 24098 3070
rect 24154 3014 24180 3070
rect 24236 3014 24261 3070
rect 24317 3014 24342 3070
rect 24398 3014 24423 3070
rect 24479 3014 24504 3070
rect 24560 3014 24585 3070
rect 24641 3014 24666 3070
rect 24722 3014 24739 3070
rect 3012 2966 24739 3014
rect 3012 2910 3036 2966
rect 3092 2910 3118 2966
rect 3174 2910 3199 2966
rect 3255 2910 3280 2966
rect 3336 2910 3361 2966
rect 3417 2910 3442 2966
rect 3498 2910 3523 2966
rect 3579 2910 3604 2966
rect 3660 2910 3686 2966
rect 3742 2910 3767 2966
rect 3823 2910 3848 2966
rect 3904 2910 3929 2966
rect 3985 2910 4010 2966
rect 4066 2910 4091 2966
rect 4147 2910 4172 2966
rect 4228 2910 4254 2966
rect 4310 2910 4335 2966
rect 4391 2910 4416 2966
rect 4472 2910 4497 2966
rect 4553 2910 4578 2966
rect 4634 2910 4659 2966
rect 4715 2910 4740 2966
rect 4796 2910 4822 2966
rect 4878 2910 4903 2966
rect 4959 2910 4984 2966
rect 5040 2910 5065 2966
rect 5121 2910 5146 2966
rect 5202 2910 5227 2966
rect 5283 2910 5308 2966
rect 5364 2910 5390 2966
rect 5446 2910 5471 2966
rect 5527 2910 5552 2966
rect 5608 2910 5633 2966
rect 5689 2910 5714 2966
rect 5770 2910 5795 2966
rect 5851 2910 5876 2966
rect 5932 2910 5958 2966
rect 6014 2910 6039 2966
rect 6095 2910 6120 2966
rect 6176 2910 6201 2966
rect 6257 2910 6282 2966
rect 6338 2910 6363 2966
rect 6419 2910 6444 2966
rect 6500 2910 6526 2966
rect 6582 2910 6607 2966
rect 6663 2910 6688 2966
rect 6744 2910 6769 2966
rect 6825 2910 6850 2966
rect 6906 2910 6931 2966
rect 6987 2910 7012 2966
rect 7068 2910 7094 2966
rect 7150 2910 7175 2966
rect 7231 2910 7256 2966
rect 7312 2910 7337 2966
rect 7393 2910 7418 2966
rect 7474 2910 7499 2966
rect 7555 2910 7580 2966
rect 7636 2910 7662 2966
rect 7718 2910 7743 2966
rect 7799 2910 7824 2966
rect 7880 2910 7905 2966
rect 7961 2910 7986 2966
rect 8042 2910 8067 2966
rect 8123 2910 8148 2966
rect 8204 2910 8230 2966
rect 8286 2910 8311 2966
rect 8367 2910 8392 2966
rect 8448 2910 8473 2966
rect 8529 2910 8554 2966
rect 8610 2910 8635 2966
rect 8691 2910 8716 2966
rect 8772 2910 8798 2966
rect 8854 2910 8879 2966
rect 8935 2910 8960 2966
rect 9016 2910 9041 2966
rect 9097 2910 9122 2966
rect 9178 2910 9203 2966
rect 9259 2910 9284 2966
rect 9340 2910 9366 2966
rect 9422 2910 9447 2966
rect 9503 2910 9528 2966
rect 9584 2910 9609 2966
rect 9665 2910 9690 2966
rect 9746 2910 9771 2966
rect 9827 2910 9852 2966
rect 9908 2910 9934 2966
rect 9990 2910 10015 2966
rect 10071 2910 10096 2966
rect 10152 2910 10177 2966
rect 10233 2910 10258 2966
rect 10314 2910 10339 2966
rect 10395 2910 10420 2966
rect 10476 2910 10502 2966
rect 10558 2910 10583 2966
rect 10639 2910 10664 2966
rect 10720 2910 10745 2966
rect 10801 2910 10826 2966
rect 10882 2910 10907 2966
rect 10963 2910 10988 2966
rect 11044 2910 11116 2966
rect 11172 2910 11197 2966
rect 11253 2910 11278 2966
rect 11334 2910 11359 2966
rect 11415 2910 11440 2966
rect 11496 2910 11521 2966
rect 11577 2910 11602 2966
rect 11658 2910 11684 2966
rect 11740 2910 11765 2966
rect 11821 2910 11846 2966
rect 11902 2910 11927 2966
rect 11983 2910 12008 2966
rect 12064 2910 12089 2966
rect 12145 2910 12170 2966
rect 12226 2910 12252 2966
rect 12308 2910 12333 2966
rect 12389 2910 12414 2966
rect 12470 2910 12495 2966
rect 12551 2910 12576 2966
rect 12632 2910 12657 2966
rect 12713 2910 12738 2966
rect 12794 2910 12820 2966
rect 12876 2910 12901 2966
rect 12957 2910 12982 2966
rect 13038 2910 13063 2966
rect 13119 2910 13144 2966
rect 13200 2910 13225 2966
rect 13281 2910 13306 2966
rect 13362 2910 13388 2966
rect 13444 2910 13469 2966
rect 13525 2910 13550 2966
rect 13606 2910 13631 2966
rect 13687 2910 13712 2966
rect 13768 2910 13793 2966
rect 13849 2910 13874 2966
rect 13930 2910 13956 2966
rect 14012 2910 14037 2966
rect 14093 2910 14118 2966
rect 14174 2910 14199 2966
rect 14255 2910 14280 2966
rect 14336 2910 14361 2966
rect 14417 2910 14442 2966
rect 14498 2910 14524 2966
rect 14580 2910 14605 2966
rect 14661 2910 14686 2966
rect 14742 2910 14767 2966
rect 14823 2910 14848 2966
rect 14904 2910 14929 2966
rect 14985 2910 15010 2966
rect 15066 2910 15092 2966
rect 15148 2910 15173 2966
rect 15229 2910 15254 2966
rect 15310 2910 15335 2966
rect 15391 2910 15416 2966
rect 15472 2910 15497 2966
rect 15553 2910 15578 2966
rect 15634 2910 15660 2966
rect 15716 2910 15741 2966
rect 15797 2910 15822 2966
rect 15878 2910 15903 2966
rect 15959 2910 15984 2966
rect 16040 2910 16065 2966
rect 16121 2910 16146 2966
rect 16202 2910 16228 2966
rect 16284 2910 16309 2966
rect 16365 2910 16390 2966
rect 16446 2910 16471 2966
rect 16527 2910 16552 2966
rect 16608 2910 16633 2966
rect 16689 2910 16714 2966
rect 16770 2910 16796 2966
rect 16852 2910 16877 2966
rect 16933 2910 16958 2966
rect 17014 2910 17039 2966
rect 17095 2910 17120 2966
rect 17176 2910 17201 2966
rect 17257 2910 17282 2966
rect 17338 2910 17364 2966
rect 17420 2910 17445 2966
rect 17501 2910 17526 2966
rect 17582 2910 17607 2966
rect 17663 2910 17688 2966
rect 17744 2910 17769 2966
rect 17825 2910 17850 2966
rect 17906 2910 17932 2966
rect 17988 2910 18013 2966
rect 18069 2910 18094 2966
rect 18150 2910 18175 2966
rect 18231 2910 18256 2966
rect 18312 2910 18337 2966
rect 18393 2910 18418 2966
rect 18474 2910 18500 2966
rect 18556 2910 18581 2966
rect 18637 2910 18662 2966
rect 18718 2910 18743 2966
rect 18799 2910 18824 2966
rect 18880 2910 18905 2966
rect 18961 2910 18986 2966
rect 19042 2910 19068 2966
rect 19124 2910 19149 2966
rect 19205 2910 19230 2966
rect 19286 2910 19311 2966
rect 19367 2910 19392 2966
rect 19448 2910 19473 2966
rect 19529 2910 19554 2966
rect 19610 2910 19636 2966
rect 19692 2910 19717 2966
rect 19773 2910 19798 2966
rect 19854 2910 19879 2966
rect 19935 2910 19960 2966
rect 20016 2910 20041 2966
rect 20097 2910 20122 2966
rect 20178 2910 20204 2966
rect 20260 2910 20285 2966
rect 20341 2910 20366 2966
rect 20422 2910 20447 2966
rect 20503 2910 20528 2966
rect 20584 2910 20609 2966
rect 20665 2910 20690 2966
rect 20746 2910 20772 2966
rect 20828 2910 20853 2966
rect 20909 2910 20934 2966
rect 20990 2910 21015 2966
rect 21071 2910 21096 2966
rect 21152 2910 21177 2966
rect 21233 2910 21258 2966
rect 21314 2910 21340 2966
rect 21396 2910 21421 2966
rect 21477 2910 21502 2966
rect 21558 2910 21583 2966
rect 21639 2910 21664 2966
rect 21720 2910 21745 2966
rect 21801 2910 21826 2966
rect 21882 2910 21908 2966
rect 21964 2910 21989 2966
rect 22045 2910 22070 2966
rect 22126 2910 22151 2966
rect 22207 2910 22232 2966
rect 22288 2910 22313 2966
rect 22369 2910 22394 2966
rect 22450 2910 22476 2966
rect 22532 2910 22557 2966
rect 22613 2910 22638 2966
rect 22694 2910 22719 2966
rect 22775 2910 22800 2966
rect 22856 2910 22881 2966
rect 22937 2910 22962 2966
rect 23018 2910 23044 2966
rect 23100 2910 23125 2966
rect 23181 2910 23206 2966
rect 23262 2910 23287 2966
rect 23343 2910 23368 2966
rect 23424 2910 23449 2966
rect 23505 2910 23530 2966
rect 23586 2910 23612 2966
rect 23668 2910 23693 2966
rect 23749 2910 23774 2966
rect 23830 2910 23855 2966
rect 23911 2910 23936 2966
rect 23992 2910 24017 2966
rect 24073 2910 24098 2966
rect 24154 2910 24180 2966
rect 24236 2910 24261 2966
rect 24317 2910 24342 2966
rect 24398 2910 24423 2966
rect 24479 2910 24504 2966
rect 24560 2910 24585 2966
rect 24641 2910 24666 2966
rect 24722 2910 24739 2966
rect 3012 2905 24739 2910
rect 6905 2667 6981 2672
rect 6905 2107 6915 2667
rect 6971 2107 6981 2667
rect 6905 1601 6981 2107
rect 7141 2667 7217 2672
rect 7141 2107 7151 2667
rect 7207 2107 7217 2667
rect 7141 1601 7217 2107
rect 7377 2667 7453 2672
rect 7377 2107 7387 2667
rect 7443 2107 7453 2667
rect 7377 1601 7453 2107
rect 7613 2667 7689 2672
rect 7613 2107 7623 2667
rect 7679 2107 7689 2667
rect 7613 1601 7689 2107
rect 7849 2667 7925 2672
rect 7849 2107 7859 2667
rect 7915 2107 7925 2667
rect 7849 1601 7925 2107
rect 8085 2667 8161 2672
rect 8085 2107 8095 2667
rect 8151 2107 8161 2667
rect 8085 1601 8161 2107
rect 8321 2667 8397 2672
rect 8321 2107 8331 2667
rect 8387 2107 8397 2667
rect 8321 1601 8397 2107
rect 8557 2667 8633 2672
rect 8557 2107 8567 2667
rect 8623 2107 8633 2667
rect 8557 1601 8633 2107
rect 8903 2667 8979 2672
rect 8903 2107 8913 2667
rect 8969 2107 8979 2667
rect 8903 1601 8979 2107
rect 9139 2667 9215 2672
rect 9139 2107 9149 2667
rect 9205 2107 9215 2667
rect 9139 1601 9215 2107
rect 9375 2667 9451 2672
rect 9375 2107 9385 2667
rect 9441 2107 9451 2667
rect 9375 1601 9451 2107
rect 9611 2667 9687 2672
rect 9611 2107 9621 2667
rect 9677 2107 9687 2667
rect 9611 1601 9687 2107
rect 9847 2667 9923 2672
rect 9847 2107 9857 2667
rect 9913 2107 9923 2667
rect 9847 1601 9923 2107
rect 10083 2667 10159 2672
rect 10083 2107 10093 2667
rect 10149 2107 10159 2667
rect 10083 1601 10159 2107
rect 10319 2667 10395 2672
rect 10319 2107 10329 2667
rect 10385 2107 10395 2667
rect 10319 1601 10395 2107
rect 10555 2667 10631 2672
rect 10555 2107 10565 2667
rect 10621 2107 10631 2667
rect 12597 2666 12673 2671
rect 12833 2666 12909 2671
rect 13069 2666 13145 2671
rect 13305 2666 13381 2671
rect 13541 2666 13617 2671
rect 13777 2666 13853 2671
rect 14013 2666 14089 2671
rect 14249 2666 14325 2671
rect 14485 2666 14561 2671
rect 14721 2666 14797 2671
rect 14957 2666 15033 2671
rect 15193 2666 15269 2671
rect 15429 2666 15505 2671
rect 16720 2666 16796 2671
rect 16956 2666 17032 2671
rect 17192 2666 17268 2671
rect 17428 2666 17504 2671
rect 17664 2666 17740 2671
rect 17900 2666 17976 2671
rect 18136 2666 18212 2671
rect 18372 2666 18448 2671
rect 18608 2666 18684 2671
rect 18844 2666 18920 2671
rect 19080 2666 19156 2671
rect 19316 2666 19392 2671
rect 19552 2666 19628 2671
rect 20843 2666 20919 2671
rect 21079 2666 21155 2671
rect 21315 2666 21391 2671
rect 21551 2666 21627 2671
rect 21787 2666 21863 2671
rect 22023 2666 22099 2671
rect 22259 2666 22335 2671
rect 22495 2666 22571 2671
rect 22731 2666 22807 2671
rect 22967 2666 23043 2671
rect 23203 2666 23279 2671
rect 23439 2666 23515 2671
rect 23675 2666 23751 2671
rect 10555 1601 10631 2107
rect 12593 2106 12603 2666
rect 12667 2106 12677 2666
rect 12829 2106 12839 2666
rect 12903 2106 12913 2666
rect 13065 2106 13075 2666
rect 13139 2106 13149 2666
rect 13301 2106 13311 2666
rect 13375 2106 13385 2666
rect 13537 2106 13547 2666
rect 13611 2106 13621 2666
rect 13773 2106 13783 2666
rect 13847 2106 13857 2666
rect 14009 2106 14019 2666
rect 14083 2106 14093 2666
rect 14245 2106 14255 2666
rect 14319 2106 14329 2666
rect 14481 2106 14491 2666
rect 14555 2106 14565 2666
rect 14717 2106 14727 2666
rect 14791 2106 14801 2666
rect 14953 2106 14963 2666
rect 15027 2106 15037 2666
rect 15189 2106 15199 2666
rect 15263 2106 15273 2666
rect 15425 2106 15435 2666
rect 15499 2106 15509 2666
rect 16716 2106 16726 2666
rect 16790 2106 16800 2666
rect 16952 2106 16962 2666
rect 17026 2106 17036 2666
rect 17188 2106 17198 2666
rect 17262 2106 17272 2666
rect 17424 2106 17434 2666
rect 17498 2106 17508 2666
rect 17660 2106 17670 2666
rect 17734 2106 17744 2666
rect 17896 2106 17906 2666
rect 17970 2106 17980 2666
rect 18132 2106 18142 2666
rect 18206 2106 18216 2666
rect 18368 2106 18378 2666
rect 18442 2106 18452 2666
rect 18604 2106 18614 2666
rect 18678 2106 18688 2666
rect 18840 2106 18850 2666
rect 18914 2106 18924 2666
rect 19076 2106 19086 2666
rect 19150 2106 19160 2666
rect 19312 2106 19322 2666
rect 19386 2106 19396 2666
rect 19548 2106 19558 2666
rect 19622 2106 19632 2666
rect 20839 2106 20849 2666
rect 20913 2106 20923 2666
rect 21075 2106 21085 2666
rect 21149 2106 21159 2666
rect 21311 2106 21321 2666
rect 21385 2106 21395 2666
rect 21547 2106 21557 2666
rect 21621 2106 21631 2666
rect 21783 2106 21793 2666
rect 21857 2106 21867 2666
rect 22019 2106 22029 2666
rect 22093 2106 22103 2666
rect 22255 2106 22265 2666
rect 22329 2106 22339 2666
rect 22491 2106 22501 2666
rect 22565 2106 22575 2666
rect 22727 2106 22737 2666
rect 22801 2106 22811 2666
rect 22963 2106 22973 2666
rect 23037 2106 23047 2666
rect 23199 2106 23209 2666
rect 23273 2106 23283 2666
rect 23435 2106 23445 2666
rect 23509 2106 23519 2666
rect 23671 2106 23681 2666
rect 23745 2106 23755 2666
rect 12597 2101 12673 2106
rect 12833 2101 12909 2106
rect 13069 2101 13145 2106
rect 13305 2101 13381 2106
rect 13541 2101 13617 2106
rect 13777 2101 13853 2106
rect 14013 2101 14089 2106
rect 14249 2101 14325 2106
rect 14485 2101 14561 2106
rect 14721 2101 14797 2106
rect 14957 2101 15033 2106
rect 15193 2101 15269 2106
rect 15429 2101 15505 2106
rect 16720 2101 16796 2106
rect 16956 2101 17032 2106
rect 17192 2101 17268 2106
rect 17428 2101 17504 2106
rect 17664 2101 17740 2106
rect 17900 2101 17976 2106
rect 18136 2101 18212 2106
rect 18372 2101 18448 2106
rect 18608 2101 18684 2106
rect 18844 2101 18920 2106
rect 19080 2101 19156 2106
rect 19316 2101 19392 2106
rect 19552 2101 19628 2106
rect 20843 2101 20919 2106
rect 21079 2101 21155 2106
rect 21315 2101 21391 2106
rect 21551 2101 21627 2106
rect 21787 2101 21863 2106
rect 22023 2101 22099 2106
rect 22259 2101 22335 2106
rect 22495 2101 22571 2106
rect 22731 2101 22807 2106
rect 22967 2101 23043 2106
rect 23203 2101 23279 2106
rect 23439 2101 23515 2106
rect 23675 2101 23751 2106
rect 12597 1830 12673 1835
rect 12833 1830 12909 1835
rect 13069 1830 13145 1835
rect 13305 1830 13381 1835
rect 13541 1830 13617 1835
rect 13777 1830 13853 1835
rect 14013 1830 14089 1835
rect 14249 1830 14325 1835
rect 14485 1830 14561 1835
rect 14721 1830 14797 1835
rect 14957 1830 15033 1835
rect 15193 1830 15269 1835
rect 15429 1830 15505 1835
rect 16720 1830 16796 1835
rect 16956 1830 17032 1835
rect 17192 1830 17268 1835
rect 17428 1830 17504 1835
rect 17664 1830 17740 1835
rect 17900 1830 17976 1835
rect 18136 1830 18212 1835
rect 18372 1830 18448 1835
rect 18608 1830 18684 1835
rect 18844 1830 18920 1835
rect 19080 1830 19156 1835
rect 19316 1830 19392 1835
rect 19552 1830 19628 1835
rect 20843 1830 20919 1835
rect 21079 1830 21155 1835
rect 21315 1830 21391 1835
rect 21551 1830 21627 1835
rect 21787 1830 21863 1835
rect 22023 1830 22099 1835
rect 22259 1830 22335 1835
rect 22495 1830 22571 1835
rect 22731 1830 22807 1835
rect 22967 1830 23043 1835
rect 23203 1830 23279 1835
rect 23439 1830 23515 1835
rect 23675 1830 23751 1835
rect 4760 1593 11628 1601
rect 4760 1537 4775 1593
rect 4831 1537 4856 1593
rect 4912 1537 4937 1593
rect 4993 1537 5018 1593
rect 5074 1537 5099 1593
rect 5155 1537 5180 1593
rect 5236 1537 5261 1593
rect 5317 1537 5363 1593
rect 5419 1537 5444 1593
rect 5500 1537 5525 1593
rect 5581 1537 5606 1593
rect 5662 1537 5687 1593
rect 5743 1537 5768 1593
rect 5824 1537 5849 1593
rect 5905 1537 5951 1593
rect 6007 1537 6032 1593
rect 6088 1537 6113 1593
rect 6169 1537 6194 1593
rect 6250 1537 6275 1593
rect 6331 1537 6356 1593
rect 6412 1537 6437 1593
rect 6493 1537 6517 1593
rect 6573 1537 6598 1593
rect 6654 1537 6679 1593
rect 6735 1537 6760 1593
rect 6816 1537 6841 1593
rect 6897 1537 6922 1593
rect 6978 1537 7003 1593
rect 7059 1537 7090 1593
rect 7146 1537 7171 1593
rect 7227 1537 7252 1593
rect 7308 1537 7333 1593
rect 7389 1537 7414 1593
rect 7470 1537 7495 1593
rect 7551 1537 7576 1593
rect 7632 1537 7656 1593
rect 7712 1537 7737 1593
rect 7793 1537 7818 1593
rect 7874 1537 7899 1593
rect 7955 1537 7980 1593
rect 8036 1537 8061 1593
rect 8117 1537 8142 1593
rect 8198 1537 8222 1593
rect 8278 1537 8303 1593
rect 8359 1537 8384 1593
rect 8440 1537 8465 1593
rect 8521 1537 8546 1593
rect 8602 1537 8627 1593
rect 8683 1537 8708 1593
rect 8764 1537 8788 1593
rect 8844 1537 8869 1593
rect 8925 1537 8950 1593
rect 9006 1537 9031 1593
rect 9087 1537 9112 1593
rect 9168 1537 9193 1593
rect 9249 1537 9274 1593
rect 9330 1537 9357 1593
rect 9413 1537 9438 1593
rect 9494 1537 9519 1593
rect 9575 1537 9600 1593
rect 9656 1537 9681 1593
rect 9737 1537 9762 1593
rect 9818 1537 9843 1593
rect 9899 1537 9923 1593
rect 9979 1537 10004 1593
rect 10060 1537 10085 1593
rect 10141 1537 10166 1593
rect 10222 1537 10247 1593
rect 10303 1537 10328 1593
rect 10384 1537 10409 1593
rect 10465 1537 10489 1593
rect 10545 1537 10570 1593
rect 10626 1537 10651 1593
rect 10707 1537 10732 1593
rect 10788 1537 10813 1593
rect 10869 1537 10894 1593
rect 10950 1537 10975 1593
rect 11031 1537 11055 1593
rect 11111 1537 11136 1593
rect 11192 1537 11217 1593
rect 11273 1537 11298 1593
rect 11354 1537 11379 1593
rect 11435 1537 11460 1593
rect 11516 1537 11541 1593
rect 11597 1537 11628 1593
rect 4760 1489 11628 1537
rect 4760 1433 4775 1489
rect 4831 1433 4856 1489
rect 4912 1433 4937 1489
rect 4993 1433 5018 1489
rect 5074 1433 5099 1489
rect 5155 1433 5180 1489
rect 5236 1433 5261 1489
rect 5317 1433 5363 1489
rect 5419 1433 5444 1489
rect 5500 1433 5525 1489
rect 5581 1433 5606 1489
rect 5662 1433 5687 1489
rect 5743 1433 5768 1489
rect 5824 1433 5849 1489
rect 5905 1433 5951 1489
rect 6007 1433 6032 1489
rect 6088 1433 6113 1489
rect 6169 1433 6194 1489
rect 6250 1433 6275 1489
rect 6331 1433 6356 1489
rect 6412 1433 6437 1489
rect 6493 1433 6517 1489
rect 6573 1433 6598 1489
rect 6654 1433 6679 1489
rect 6735 1433 6760 1489
rect 6816 1433 6841 1489
rect 6897 1433 6922 1489
rect 6978 1433 7003 1489
rect 7059 1433 7090 1489
rect 7146 1433 7171 1489
rect 7227 1433 7252 1489
rect 7308 1433 7333 1489
rect 7389 1433 7414 1489
rect 7470 1433 7495 1489
rect 7551 1433 7576 1489
rect 7632 1433 7656 1489
rect 7712 1433 7737 1489
rect 7793 1433 7818 1489
rect 7874 1433 7899 1489
rect 7955 1433 7980 1489
rect 8036 1433 8061 1489
rect 8117 1433 8142 1489
rect 8198 1433 8222 1489
rect 8278 1433 8303 1489
rect 8359 1433 8384 1489
rect 8440 1433 8465 1489
rect 8521 1433 8546 1489
rect 8602 1433 8627 1489
rect 8683 1433 8708 1489
rect 8764 1433 8788 1489
rect 8844 1433 8869 1489
rect 8925 1433 8950 1489
rect 9006 1433 9031 1489
rect 9087 1433 9112 1489
rect 9168 1433 9193 1489
rect 9249 1433 9274 1489
rect 9330 1433 9357 1489
rect 9413 1433 9438 1489
rect 9494 1433 9519 1489
rect 9575 1433 9600 1489
rect 9656 1433 9681 1489
rect 9737 1433 9762 1489
rect 9818 1433 9843 1489
rect 9899 1433 9923 1489
rect 9979 1433 10004 1489
rect 10060 1433 10085 1489
rect 10141 1433 10166 1489
rect 10222 1433 10247 1489
rect 10303 1433 10328 1489
rect 10384 1433 10409 1489
rect 10465 1433 10489 1489
rect 10545 1433 10570 1489
rect 10626 1433 10651 1489
rect 10707 1433 10732 1489
rect 10788 1433 10813 1489
rect 10869 1433 10894 1489
rect 10950 1433 10975 1489
rect 11031 1433 11055 1489
rect 11111 1433 11136 1489
rect 11192 1433 11217 1489
rect 11273 1433 11298 1489
rect 11354 1433 11379 1489
rect 11435 1433 11460 1489
rect 11516 1433 11541 1489
rect 11597 1433 11628 1489
rect 4760 1385 11628 1433
rect 4760 1329 4775 1385
rect 4831 1329 4856 1385
rect 4912 1329 4937 1385
rect 4993 1329 5018 1385
rect 5074 1329 5099 1385
rect 5155 1329 5180 1385
rect 5236 1329 5261 1385
rect 5317 1329 5363 1385
rect 5419 1329 5444 1385
rect 5500 1329 5525 1385
rect 5581 1329 5606 1385
rect 5662 1329 5687 1385
rect 5743 1329 5768 1385
rect 5824 1329 5849 1385
rect 5905 1329 5951 1385
rect 6007 1329 6032 1385
rect 6088 1329 6113 1385
rect 6169 1329 6194 1385
rect 6250 1329 6275 1385
rect 6331 1329 6356 1385
rect 6412 1329 6437 1385
rect 6493 1329 6517 1385
rect 6573 1329 6598 1385
rect 6654 1329 6679 1385
rect 6735 1329 6760 1385
rect 6816 1329 6841 1385
rect 6897 1329 6922 1385
rect 6978 1329 7003 1385
rect 7059 1329 7090 1385
rect 7146 1329 7171 1385
rect 7227 1329 7252 1385
rect 7308 1329 7333 1385
rect 7389 1329 7414 1385
rect 7470 1329 7495 1385
rect 7551 1329 7576 1385
rect 7632 1329 7656 1385
rect 7712 1329 7737 1385
rect 7793 1329 7818 1385
rect 7874 1329 7899 1385
rect 7955 1329 7980 1385
rect 8036 1329 8061 1385
rect 8117 1329 8142 1385
rect 8198 1329 8222 1385
rect 8278 1329 8303 1385
rect 8359 1329 8384 1385
rect 8440 1329 8465 1385
rect 8521 1329 8546 1385
rect 8602 1329 8627 1385
rect 8683 1329 8708 1385
rect 8764 1329 8788 1385
rect 8844 1329 8869 1385
rect 8925 1329 8950 1385
rect 9006 1329 9031 1385
rect 9087 1329 9112 1385
rect 9168 1329 9193 1385
rect 9249 1329 9274 1385
rect 9330 1329 9357 1385
rect 9413 1329 9438 1385
rect 9494 1329 9519 1385
rect 9575 1329 9600 1385
rect 9656 1329 9681 1385
rect 9737 1329 9762 1385
rect 9818 1329 9843 1385
rect 9899 1329 9923 1385
rect 9979 1329 10004 1385
rect 10060 1329 10085 1385
rect 10141 1329 10166 1385
rect 10222 1329 10247 1385
rect 10303 1329 10328 1385
rect 10384 1329 10409 1385
rect 10465 1329 10489 1385
rect 10545 1329 10570 1385
rect 10626 1329 10651 1385
rect 10707 1329 10732 1385
rect 10788 1329 10813 1385
rect 10869 1329 10894 1385
rect 10950 1329 10975 1385
rect 11031 1329 11055 1385
rect 11111 1329 11136 1385
rect 11192 1329 11217 1385
rect 11273 1329 11298 1385
rect 11354 1329 11379 1385
rect 11435 1329 11460 1385
rect 11516 1329 11541 1385
rect 11597 1329 11628 1385
rect 4760 1319 11628 1329
rect 12593 1270 12603 1830
rect 12667 1270 12677 1830
rect 12829 1270 12839 1830
rect 12903 1270 12913 1830
rect 13065 1270 13075 1830
rect 13139 1270 13149 1830
rect 13301 1270 13311 1830
rect 13375 1270 13385 1830
rect 13537 1270 13547 1830
rect 13611 1270 13621 1830
rect 13773 1270 13783 1830
rect 13847 1270 13857 1830
rect 14009 1270 14019 1830
rect 14083 1270 14093 1830
rect 14245 1270 14255 1830
rect 14319 1270 14329 1830
rect 14481 1270 14491 1830
rect 14555 1270 14565 1830
rect 14717 1270 14727 1830
rect 14791 1270 14801 1830
rect 14953 1270 14963 1830
rect 15027 1270 15037 1830
rect 15189 1270 15199 1830
rect 15263 1270 15273 1830
rect 15425 1270 15435 1830
rect 15499 1270 15509 1830
rect 16716 1270 16726 1830
rect 16790 1270 16800 1830
rect 16952 1270 16962 1830
rect 17026 1270 17036 1830
rect 17188 1270 17198 1830
rect 17262 1270 17272 1830
rect 17424 1270 17434 1830
rect 17498 1270 17508 1830
rect 17660 1270 17670 1830
rect 17734 1270 17744 1830
rect 17896 1270 17906 1830
rect 17970 1270 17980 1830
rect 18132 1270 18142 1830
rect 18206 1270 18216 1830
rect 18368 1270 18378 1830
rect 18442 1270 18452 1830
rect 18604 1270 18614 1830
rect 18678 1270 18688 1830
rect 18840 1270 18850 1830
rect 18914 1270 18924 1830
rect 19076 1270 19086 1830
rect 19150 1270 19160 1830
rect 19312 1270 19322 1830
rect 19386 1270 19396 1830
rect 19548 1270 19558 1830
rect 19622 1270 19632 1830
rect 20839 1270 20849 1830
rect 20913 1270 20923 1830
rect 21075 1270 21085 1830
rect 21149 1270 21159 1830
rect 21311 1270 21321 1830
rect 21385 1270 21395 1830
rect 21547 1270 21557 1830
rect 21621 1270 21631 1830
rect 21783 1270 21793 1830
rect 21857 1270 21867 1830
rect 22019 1270 22029 1830
rect 22093 1270 22103 1830
rect 22255 1270 22265 1830
rect 22329 1270 22339 1830
rect 22491 1270 22501 1830
rect 22565 1270 22575 1830
rect 22727 1270 22737 1830
rect 22801 1270 22811 1830
rect 22963 1270 22973 1830
rect 23037 1270 23047 1830
rect 23199 1270 23209 1830
rect 23273 1270 23283 1830
rect 23435 1270 23445 1830
rect 23509 1270 23519 1830
rect 23671 1270 23681 1830
rect 23745 1270 23755 1830
rect 12597 1265 12673 1270
rect 12833 1265 12909 1270
rect 13069 1265 13145 1270
rect 13305 1265 13381 1270
rect 13541 1265 13617 1270
rect 13777 1265 13853 1270
rect 14013 1265 14089 1270
rect 14249 1265 14325 1270
rect 14485 1265 14561 1270
rect 14721 1265 14797 1270
rect 14957 1265 15033 1270
rect 15193 1265 15269 1270
rect 15429 1265 15505 1270
rect 16720 1265 16796 1270
rect 16956 1265 17032 1270
rect 17192 1265 17268 1270
rect 17428 1265 17504 1270
rect 17664 1265 17740 1270
rect 17900 1265 17976 1270
rect 18136 1265 18212 1270
rect 18372 1265 18448 1270
rect 18608 1265 18684 1270
rect 18844 1265 18920 1270
rect 19080 1265 19156 1270
rect 19316 1265 19392 1270
rect 19552 1265 19628 1270
rect 20843 1265 20919 1270
rect 21079 1265 21155 1270
rect 21315 1265 21391 1270
rect 21551 1265 21627 1270
rect 21787 1265 21863 1270
rect 22023 1265 22099 1270
rect 22259 1265 22335 1270
rect 22495 1265 22571 1270
rect 22731 1265 22807 1270
rect 22967 1265 23043 1270
rect 23203 1265 23279 1270
rect 23439 1265 23515 1270
rect 23675 1265 23751 1270
rect 4901 1170 10649 1175
rect 4901 610 4911 1170
rect 4975 610 5147 1170
rect 5211 610 5383 1170
rect 5447 610 5619 1170
rect 5683 610 5855 1170
rect 5919 610 6091 1170
rect 6155 610 6327 1170
rect 6391 610 6563 1170
rect 6627 610 6799 1170
rect 6863 610 7035 1170
rect 7099 610 7271 1170
rect 7335 610 7507 1170
rect 7571 610 7747 1170
rect 7803 610 7983 1170
rect 8039 610 8219 1170
rect 8275 610 8455 1170
rect 8511 610 8691 1170
rect 8747 610 8927 1170
rect 8983 610 9163 1170
rect 9219 610 9399 1170
rect 9455 610 9635 1170
rect 9691 610 9871 1170
rect 9927 610 10107 1170
rect 10163 610 10343 1170
rect 10399 610 10579 1170
rect 10635 610 10649 1170
rect 4901 605 10649 610
rect 12374 586 23886 970
rect 8688 339 8753 340
rect 8923 339 8988 340
rect 9157 339 9225 340
rect 10104 339 10169 340
rect 4901 334 10649 339
rect 4901 -226 4911 334
rect 4975 -226 5147 334
rect 5211 -226 5383 334
rect 5447 -226 5619 334
rect 5683 -226 5855 334
rect 5919 -226 6091 334
rect 6155 -226 6327 334
rect 6391 -226 6563 334
rect 6627 -226 6799 334
rect 6863 -226 7035 334
rect 7099 -226 7271 334
rect 7335 -226 7507 334
rect 7571 -226 7747 334
rect 7803 -226 7983 334
rect 8039 -226 8219 334
rect 8275 -226 8455 334
rect 8511 -226 8691 334
rect 8747 -226 8927 334
rect 8983 -226 9163 334
rect 9219 -226 9399 334
rect 9455 -226 9635 334
rect 9691 -226 9871 334
rect 9927 -226 10107 334
rect 10163 -226 10343 334
rect 10399 -226 10579 334
rect 10635 -226 10649 334
rect 4901 -231 10649 -226
rect 4901 -880 10649 -875
rect 4901 -1440 4911 -880
rect 4975 -1440 5147 -880
rect 5211 -1440 5383 -880
rect 5447 -1440 5619 -880
rect 5683 -1440 5855 -880
rect 5919 -1440 6091 -880
rect 6155 -1440 6327 -880
rect 6391 -1440 6563 -880
rect 6627 -1440 6799 -880
rect 6863 -1440 7035 -880
rect 7099 -1440 7271 -880
rect 7335 -1440 7507 -880
rect 7571 -1440 7747 -880
rect 7803 -1440 7983 -880
rect 8039 -1440 8219 -880
rect 8275 -1440 8455 -880
rect 8511 -1440 8691 -880
rect 8747 -1440 8927 -880
rect 8983 -1440 9163 -880
rect 9219 -1440 9399 -880
rect 9455 -1440 9635 -880
rect 9691 -1440 9871 -880
rect 9927 -1440 10107 -880
rect 10163 -1440 10343 -880
rect 10399 -1440 10579 -880
rect 10635 -1440 10649 -880
rect 4901 -1445 10649 -1440
rect 8688 -1711 8753 -1710
rect 8923 -1711 8988 -1710
rect 9157 -1711 9225 -1710
rect 10104 -1711 10169 -1710
rect 4901 -1716 10649 -1711
rect 4901 -2276 4911 -1716
rect 4975 -2276 5147 -1716
rect 5211 -2276 5383 -1716
rect 5447 -2276 5619 -1716
rect 5683 -2276 5855 -1716
rect 5919 -2276 6091 -1716
rect 6155 -2276 6327 -1716
rect 6391 -2276 6563 -1716
rect 6627 -2276 6799 -1716
rect 6863 -2276 7035 -1716
rect 7099 -2276 7271 -1716
rect 7335 -2276 7507 -1716
rect 7571 -2276 7747 -1716
rect 7803 -2276 7983 -1716
rect 8039 -2276 8219 -1716
rect 8275 -2276 8455 -1716
rect 8511 -2276 8691 -1716
rect 8747 -2276 8927 -1716
rect 8983 -2276 9163 -1716
rect 9219 -2276 9399 -1716
rect 9455 -2276 9635 -1716
rect 9691 -2276 9871 -1716
rect 9927 -2276 10107 -1716
rect 10163 -2276 10343 -1716
rect 10399 -2276 10579 -1716
rect 10635 -2276 10649 -1716
rect 4901 -2281 10649 -2276
rect 4905 -2930 10653 -2925
rect 4905 -3490 4919 -2930
rect 4975 -3490 5155 -2930
rect 5211 -3490 5391 -2930
rect 5447 -3490 5627 -2930
rect 5683 -3490 5863 -2930
rect 5919 -3490 6099 -2930
rect 6155 -3490 6335 -2930
rect 6391 -3490 6571 -2930
rect 6627 -3490 6807 -2930
rect 6863 -3490 7043 -2930
rect 7099 -3490 7279 -2930
rect 7335 -3490 7515 -2930
rect 7571 -3490 7751 -2930
rect 7807 -3490 7983 -2930
rect 8047 -3490 8219 -2930
rect 8283 -3490 8455 -2930
rect 8519 -3490 8691 -2930
rect 8755 -3490 8927 -2930
rect 8991 -3490 9163 -2930
rect 9227 -3490 9399 -2930
rect 9463 -3490 9635 -2930
rect 9699 -3490 9871 -2930
rect 9935 -3490 10107 -2930
rect 10171 -3490 10343 -2930
rect 10407 -3490 10579 -2930
rect 10643 -3490 10653 -2930
rect 11697 -3158 20542 -2774
rect 4905 -3495 10653 -3490
rect 5385 -3761 5450 -3760
rect 6329 -3761 6397 -3760
rect 6566 -3761 6631 -3760
rect 6801 -3761 6866 -3760
rect 4905 -3766 10653 -3761
rect 4905 -4326 4919 -3766
rect 4975 -4326 5155 -3766
rect 5211 -4326 5391 -3766
rect 5447 -4326 5627 -3766
rect 5683 -4326 5863 -3766
rect 5919 -4326 6099 -3766
rect 6155 -4326 6335 -3766
rect 6391 -4326 6571 -3766
rect 6627 -4326 6807 -3766
rect 6863 -4326 7043 -3766
rect 7099 -4326 7279 -3766
rect 7335 -4326 7515 -3766
rect 7571 -4326 7751 -3766
rect 7807 -4326 7983 -3766
rect 8047 -4326 8219 -3766
rect 8283 -4326 8455 -3766
rect 8519 -4326 8691 -3766
rect 8755 -4326 8927 -3766
rect 8991 -4326 9163 -3766
rect 9227 -4326 9399 -3766
rect 9463 -4326 9635 -3766
rect 9699 -4326 9871 -3766
rect 9935 -4326 10107 -3766
rect 10171 -4326 10343 -3766
rect 10407 -4326 10579 -3766
rect 10643 -4326 10653 -3766
rect 4905 -4331 10653 -4326
rect 4905 -4980 10653 -4975
rect 4905 -5540 4919 -4980
rect 4975 -5540 5155 -4980
rect 5211 -5540 5391 -4980
rect 5447 -5540 5627 -4980
rect 5683 -5540 5863 -4980
rect 5919 -5540 6099 -4980
rect 6155 -5540 6335 -4980
rect 6391 -5540 6571 -4980
rect 6627 -5540 6807 -4980
rect 6863 -5540 7043 -4980
rect 7099 -5540 7279 -4980
rect 7335 -5540 7515 -4980
rect 7571 -5540 7751 -4980
rect 7807 -5540 7983 -4980
rect 8047 -5540 8219 -4980
rect 8283 -5540 8455 -4980
rect 8519 -5540 8691 -4980
rect 8755 -5540 8927 -4980
rect 8991 -5540 9163 -4980
rect 9227 -5540 9399 -4980
rect 9463 -5540 9635 -4980
rect 9699 -5540 9871 -4980
rect 9935 -5540 10107 -4980
rect 10171 -5540 10343 -4980
rect 10407 -5540 10579 -4980
rect 10643 -5540 10653 -4980
rect 4905 -5545 10653 -5540
rect 5385 -5811 5450 -5810
rect 6329 -5811 6397 -5810
rect 6566 -5811 6631 -5810
rect 6801 -5811 6866 -5810
rect 4905 -5816 10653 -5811
rect 4905 -6376 4919 -5816
rect 4975 -6376 5155 -5816
rect 5211 -6376 5391 -5816
rect 5447 -6376 5627 -5816
rect 5683 -6376 5863 -5816
rect 5919 -6376 6099 -5816
rect 6155 -6376 6335 -5816
rect 6391 -6376 6571 -5816
rect 6627 -6376 6807 -5816
rect 6863 -6376 7043 -5816
rect 7099 -6376 7279 -5816
rect 7335 -6376 7515 -5816
rect 7571 -6376 7751 -5816
rect 7807 -6376 7983 -5816
rect 8047 -6376 8219 -5816
rect 8283 -6376 8455 -5816
rect 8519 -6376 8691 -5816
rect 8755 -6376 8927 -5816
rect 8991 -6376 9163 -5816
rect 9227 -6376 9399 -5816
rect 9463 -6376 9635 -5816
rect 9699 -6376 9871 -5816
rect 9935 -6376 10107 -5816
rect 10171 -6376 10343 -5816
rect 10407 -6376 10579 -5816
rect 10643 -6376 10653 -5816
rect 4905 -6381 10653 -6376
rect 11051 -6698 11639 -6693
rect 11051 -6754 11066 -6698
rect 11122 -6754 11147 -6698
rect 11203 -6754 11228 -6698
rect 11284 -6754 11309 -6698
rect 11365 -6754 11390 -6698
rect 11446 -6754 11471 -6698
rect 11527 -6754 11552 -6698
rect 11608 -6754 11639 -6698
rect 11051 -6802 11639 -6754
rect 11051 -6858 11066 -6802
rect 11122 -6858 11147 -6802
rect 11203 -6858 11228 -6802
rect 11284 -6858 11309 -6802
rect 11365 -6858 11390 -6802
rect 11446 -6858 11471 -6802
rect 11527 -6858 11552 -6802
rect 11608 -6858 11639 -6802
rect 11051 -6906 11639 -6858
rect 12374 -6906 23886 -6522
rect 11051 -6962 11066 -6906
rect 11122 -6962 11147 -6906
rect 11203 -6962 11228 -6906
rect 11284 -6962 11309 -6906
rect 11365 -6962 11390 -6906
rect 11446 -6962 11471 -6906
rect 11527 -6962 11552 -6906
rect 11608 -6962 11639 -6906
rect 11051 -6967 11639 -6962
rect 4083 -7061 5471 -7053
rect 4083 -7117 4092 -7061
rect 4148 -7117 4173 -7061
rect 4229 -7117 4254 -7061
rect 4310 -7117 4335 -7061
rect 4391 -7117 4416 -7061
rect 4472 -7117 4497 -7061
rect 4553 -7117 4578 -7061
rect 4634 -7117 4660 -7061
rect 4716 -7117 4741 -7061
rect 4797 -7117 4822 -7061
rect 4878 -7117 4903 -7061
rect 4959 -7117 4984 -7061
rect 5040 -7117 5065 -7061
rect 5121 -7117 5146 -7061
rect 5202 -7117 5228 -7061
rect 5284 -7117 5309 -7061
rect 5365 -7117 5390 -7061
rect 5446 -7117 5471 -7061
rect 4083 -7165 5471 -7117
rect 4083 -7221 4092 -7165
rect 4148 -7221 4173 -7165
rect 4229 -7221 4254 -7165
rect 4310 -7221 4335 -7165
rect 4391 -7221 4416 -7165
rect 4472 -7221 4497 -7165
rect 4553 -7221 4578 -7165
rect 4634 -7221 4660 -7165
rect 4716 -7221 4741 -7165
rect 4797 -7221 4822 -7165
rect 4878 -7221 4903 -7165
rect 4959 -7221 4984 -7165
rect 5040 -7221 5065 -7165
rect 5121 -7221 5146 -7165
rect 5202 -7221 5228 -7165
rect 5284 -7221 5309 -7165
rect 5365 -7221 5390 -7165
rect 5446 -7221 5471 -7165
rect 4083 -7269 5471 -7221
rect 5973 -7223 6049 -7218
rect 6209 -7223 6285 -7218
rect 6445 -7223 6521 -7218
rect 6681 -7223 6757 -7218
rect 6917 -7223 6993 -7218
rect 7153 -7223 7229 -7218
rect 7389 -7223 7465 -7218
rect 7625 -7223 7701 -7218
rect 7971 -7223 8047 -7218
rect 8207 -7223 8283 -7218
rect 8443 -7223 8519 -7218
rect 8679 -7223 8755 -7218
rect 8915 -7223 8991 -7218
rect 9151 -7223 9227 -7218
rect 9387 -7223 9463 -7218
rect 9623 -7223 9699 -7218
rect 12513 -7219 12589 -7214
rect 4083 -7325 4092 -7269
rect 4148 -7325 4173 -7269
rect 4229 -7325 4254 -7269
rect 4310 -7325 4335 -7269
rect 4391 -7325 4416 -7269
rect 4472 -7325 4497 -7269
rect 4553 -7325 4578 -7269
rect 4634 -7325 4660 -7269
rect 4716 -7325 4741 -7269
rect 4797 -7325 4822 -7269
rect 4878 -7325 4903 -7269
rect 4959 -7325 4984 -7269
rect 5040 -7325 5065 -7269
rect 5121 -7325 5146 -7269
rect 5202 -7325 5228 -7269
rect 5284 -7325 5309 -7269
rect 5365 -7325 5390 -7269
rect 5446 -7325 5471 -7269
rect 4083 -7373 5471 -7325
rect 4083 -7429 4092 -7373
rect 4148 -7429 4173 -7373
rect 4229 -7429 4254 -7373
rect 4310 -7429 4335 -7373
rect 4391 -7429 4416 -7373
rect 4472 -7429 4497 -7373
rect 4553 -7429 4578 -7373
rect 4634 -7429 4660 -7373
rect 4716 -7429 4741 -7373
rect 4797 -7429 4822 -7373
rect 4878 -7429 4903 -7373
rect 4959 -7429 4984 -7373
rect 5040 -7429 5065 -7373
rect 5121 -7429 5146 -7373
rect 5202 -7429 5228 -7373
rect 5284 -7429 5309 -7373
rect 5365 -7429 5390 -7373
rect 5446 -7429 5471 -7373
rect 4083 -7477 5471 -7429
rect 4083 -7533 4092 -7477
rect 4148 -7533 4173 -7477
rect 4229 -7533 4254 -7477
rect 4310 -7533 4335 -7477
rect 4391 -7533 4416 -7477
rect 4472 -7533 4497 -7477
rect 4553 -7533 4578 -7477
rect 4634 -7533 4660 -7477
rect 4716 -7533 4741 -7477
rect 4797 -7533 4822 -7477
rect 4878 -7533 4903 -7477
rect 4959 -7533 4984 -7477
rect 5040 -7533 5065 -7477
rect 5121 -7533 5146 -7477
rect 5202 -7533 5228 -7477
rect 5284 -7533 5309 -7477
rect 5365 -7533 5390 -7477
rect 5446 -7533 5471 -7477
rect 4083 -7581 5471 -7533
rect 4083 -7637 4092 -7581
rect 4148 -7637 4173 -7581
rect 4229 -7637 4254 -7581
rect 4310 -7637 4335 -7581
rect 4391 -7637 4416 -7581
rect 4472 -7637 4497 -7581
rect 4553 -7637 4578 -7581
rect 4634 -7637 4660 -7581
rect 4716 -7637 4741 -7581
rect 4797 -7637 4822 -7581
rect 4878 -7637 4903 -7581
rect 4959 -7637 4984 -7581
rect 5040 -7637 5065 -7581
rect 5121 -7637 5146 -7581
rect 5202 -7637 5228 -7581
rect 5284 -7637 5309 -7581
rect 5365 -7637 5390 -7581
rect 5446 -7637 5471 -7581
rect 4083 -7685 5471 -7637
rect 4083 -7741 4092 -7685
rect 4148 -7741 4173 -7685
rect 4229 -7741 4254 -7685
rect 4310 -7741 4335 -7685
rect 4391 -7741 4416 -7685
rect 4472 -7741 4497 -7685
rect 4553 -7741 4578 -7685
rect 4634 -7741 4660 -7685
rect 4716 -7741 4741 -7685
rect 4797 -7741 4822 -7685
rect 4878 -7741 4903 -7685
rect 4959 -7741 4984 -7685
rect 5040 -7741 5065 -7685
rect 5121 -7741 5146 -7685
rect 5202 -7741 5228 -7685
rect 5284 -7741 5309 -7685
rect 5365 -7741 5390 -7685
rect 5446 -7741 5471 -7685
rect 4083 -7789 5471 -7741
rect 5969 -7783 5979 -7223
rect 6043 -7783 6053 -7223
rect 6205 -7783 6215 -7223
rect 6279 -7783 6289 -7223
rect 6441 -7783 6451 -7223
rect 6515 -7783 6525 -7223
rect 6677 -7783 6687 -7223
rect 6751 -7783 6761 -7223
rect 6913 -7783 6923 -7223
rect 6987 -7783 6997 -7223
rect 7149 -7783 7159 -7223
rect 7223 -7783 7233 -7223
rect 7385 -7783 7395 -7223
rect 7459 -7783 7469 -7223
rect 7621 -7783 7631 -7223
rect 7695 -7783 7705 -7223
rect 7967 -7783 7977 -7223
rect 8041 -7783 8051 -7223
rect 8203 -7783 8213 -7223
rect 8277 -7783 8287 -7223
rect 8439 -7783 8449 -7223
rect 8513 -7783 8523 -7223
rect 8675 -7783 8685 -7223
rect 8749 -7783 8759 -7223
rect 8911 -7783 8921 -7223
rect 8985 -7783 8995 -7223
rect 9147 -7783 9157 -7223
rect 9221 -7783 9231 -7223
rect 9383 -7783 9393 -7223
rect 9457 -7783 9467 -7223
rect 9619 -7783 9629 -7223
rect 9693 -7783 9703 -7223
rect 10620 -7395 12266 -7390
rect 10620 -7515 10625 -7395
rect 10681 -7515 10941 -7395
rect 10997 -7515 11257 -7395
rect 11313 -7515 11573 -7395
rect 11629 -7515 11889 -7395
rect 11945 -7515 12205 -7395
rect 12261 -7515 12266 -7395
rect 10620 -7520 12266 -7515
rect 5973 -7788 6049 -7783
rect 6209 -7788 6285 -7783
rect 6445 -7788 6521 -7783
rect 6681 -7788 6757 -7783
rect 6917 -7788 6993 -7783
rect 7153 -7788 7229 -7783
rect 7389 -7788 7465 -7783
rect 7625 -7788 7701 -7783
rect 7971 -7788 8047 -7783
rect 8207 -7788 8283 -7783
rect 8443 -7788 8519 -7783
rect 8679 -7788 8755 -7783
rect 8915 -7788 8991 -7783
rect 9151 -7788 9227 -7783
rect 9387 -7788 9463 -7783
rect 9623 -7788 9699 -7783
rect 4083 -7845 4092 -7789
rect 4148 -7845 4173 -7789
rect 4229 -7845 4254 -7789
rect 4310 -7845 4335 -7789
rect 4391 -7845 4416 -7789
rect 4472 -7845 4497 -7789
rect 4553 -7845 4578 -7789
rect 4634 -7845 4660 -7789
rect 4716 -7845 4741 -7789
rect 4797 -7845 4822 -7789
rect 4878 -7845 4903 -7789
rect 4959 -7845 4984 -7789
rect 5040 -7845 5065 -7789
rect 5121 -7845 5146 -7789
rect 5202 -7845 5228 -7789
rect 5284 -7845 5309 -7789
rect 5365 -7845 5390 -7789
rect 5446 -7845 5471 -7789
rect 4083 -7893 5471 -7845
rect 4083 -7949 4092 -7893
rect 4148 -7949 4173 -7893
rect 4229 -7949 4254 -7893
rect 4310 -7949 4335 -7893
rect 4391 -7949 4416 -7893
rect 4472 -7949 4497 -7893
rect 4553 -7949 4578 -7893
rect 4634 -7949 4660 -7893
rect 4716 -7949 4741 -7893
rect 4797 -7949 4822 -7893
rect 4878 -7949 4903 -7893
rect 4959 -7949 4984 -7893
rect 5040 -7949 5065 -7893
rect 5121 -7949 5146 -7893
rect 5202 -7949 5228 -7893
rect 5284 -7949 5309 -7893
rect 5365 -7949 5390 -7893
rect 5446 -7949 5471 -7893
rect 4083 -7997 5471 -7949
rect 4083 -8053 4092 -7997
rect 4148 -8053 4173 -7997
rect 4229 -8053 4254 -7997
rect 4310 -8053 4335 -7997
rect 4391 -8053 4416 -7997
rect 4472 -8053 4497 -7997
rect 4553 -8053 4578 -7997
rect 4634 -8053 4660 -7997
rect 4716 -8053 4741 -7997
rect 4797 -8053 4822 -7997
rect 4878 -8053 4903 -7997
rect 4959 -8053 4984 -7997
rect 5040 -8053 5065 -7997
rect 5121 -8053 5146 -7997
rect 5202 -8053 5228 -7997
rect 5284 -8053 5309 -7997
rect 5365 -8053 5390 -7997
rect 5446 -8053 5471 -7997
rect 10825 -8020 11914 -8012
rect 10825 -8036 10834 -8020
rect 5973 -8041 6049 -8036
rect 6209 -8041 6285 -8036
rect 6445 -8041 6521 -8036
rect 6681 -8041 6757 -8036
rect 6917 -8041 6993 -8036
rect 7153 -8041 7229 -8036
rect 7389 -8041 7465 -8036
rect 7625 -8041 7701 -8036
rect 7967 -8041 10834 -8036
rect 4083 -8101 5471 -8053
rect 4083 -8157 4092 -8101
rect 4148 -8157 4173 -8101
rect 4229 -8157 4254 -8101
rect 4310 -8157 4335 -8101
rect 4391 -8157 4416 -8101
rect 4472 -8157 4497 -8101
rect 4553 -8157 4578 -8101
rect 4634 -8157 4660 -8101
rect 4716 -8157 4741 -8101
rect 4797 -8157 4822 -8101
rect 4878 -8157 4903 -8101
rect 4959 -8157 4984 -8101
rect 5040 -8157 5065 -8101
rect 5121 -8157 5146 -8101
rect 5202 -8157 5228 -8101
rect 5284 -8157 5309 -8101
rect 5365 -8157 5390 -8101
rect 5446 -8157 5471 -8101
rect 4083 -8205 5471 -8157
rect 4083 -8261 4092 -8205
rect 4148 -8261 4173 -8205
rect 4229 -8261 4254 -8205
rect 4310 -8261 4335 -8205
rect 4391 -8261 4416 -8205
rect 4472 -8261 4497 -8205
rect 4553 -8261 4578 -8205
rect 4634 -8261 4660 -8205
rect 4716 -8261 4741 -8205
rect 4797 -8261 4822 -8205
rect 4878 -8261 4903 -8205
rect 4959 -8261 4984 -8205
rect 5040 -8261 5065 -8205
rect 5121 -8261 5146 -8205
rect 5202 -8261 5228 -8205
rect 5284 -8261 5309 -8205
rect 5365 -8261 5390 -8205
rect 5446 -8261 5471 -8205
rect 4083 -8309 5471 -8261
rect 4083 -8365 4092 -8309
rect 4148 -8365 4173 -8309
rect 4229 -8365 4254 -8309
rect 4310 -8365 4335 -8309
rect 4391 -8365 4416 -8309
rect 4472 -8365 4497 -8309
rect 4553 -8365 4578 -8309
rect 4634 -8365 4660 -8309
rect 4716 -8365 4741 -8309
rect 4797 -8365 4822 -8309
rect 4878 -8365 4903 -8309
rect 4959 -8365 4984 -8309
rect 5040 -8365 5065 -8309
rect 5121 -8365 5146 -8309
rect 5202 -8365 5228 -8309
rect 5284 -8365 5309 -8309
rect 5365 -8365 5390 -8309
rect 5446 -8365 5471 -8309
rect 4083 -8413 5471 -8365
rect 4083 -8469 4092 -8413
rect 4148 -8469 4173 -8413
rect 4229 -8469 4254 -8413
rect 4310 -8469 4335 -8413
rect 4391 -8469 4416 -8413
rect 4472 -8469 4497 -8413
rect 4553 -8469 4578 -8413
rect 4634 -8469 4660 -8413
rect 4716 -8469 4741 -8413
rect 4797 -8469 4822 -8413
rect 4878 -8469 4903 -8413
rect 4959 -8469 4984 -8413
rect 5040 -8469 5065 -8413
rect 5121 -8469 5146 -8413
rect 5202 -8469 5228 -8413
rect 5284 -8469 5309 -8413
rect 5365 -8469 5390 -8413
rect 5446 -8417 5471 -8413
rect 5446 -8469 5472 -8417
rect 4083 -8517 5472 -8469
rect 4083 -8573 4092 -8517
rect 4148 -8573 4173 -8517
rect 4229 -8573 4254 -8517
rect 4310 -8573 4335 -8517
rect 4391 -8573 4416 -8517
rect 4472 -8573 4497 -8517
rect 4553 -8573 4578 -8517
rect 4634 -8573 4660 -8517
rect 4716 -8573 4741 -8517
rect 4797 -8573 4822 -8517
rect 4878 -8573 4903 -8517
rect 4959 -8573 4984 -8517
rect 5040 -8573 5065 -8517
rect 5121 -8573 5146 -8517
rect 5202 -8573 5228 -8517
rect 5284 -8573 5309 -8517
rect 5365 -8573 5390 -8517
rect 5446 -8573 5472 -8517
rect 4083 -8602 5472 -8573
rect 5969 -8601 5979 -8041
rect 6043 -8601 6053 -8041
rect 6205 -8601 6215 -8041
rect 6279 -8601 6289 -8041
rect 6441 -8601 6451 -8041
rect 6515 -8601 6525 -8041
rect 6677 -8601 6687 -8041
rect 6751 -8601 6761 -8041
rect 6913 -8601 6923 -8041
rect 6987 -8601 6997 -8041
rect 7149 -8601 7159 -8041
rect 7223 -8601 7233 -8041
rect 7385 -8601 7395 -8041
rect 7459 -8601 7469 -8041
rect 7621 -8601 7631 -8041
rect 7695 -8601 7705 -8041
rect 7967 -8601 7977 -8041
rect 8041 -8383 8213 -8041
rect 8041 -8601 8051 -8383
rect 8203 -8601 8213 -8383
rect 8277 -8383 8449 -8041
rect 8277 -8601 8287 -8383
rect 8439 -8601 8449 -8383
rect 8513 -8383 8685 -8041
rect 8513 -8601 8523 -8383
rect 8675 -8601 8685 -8383
rect 8749 -8383 8921 -8041
rect 8749 -8601 8759 -8383
rect 8911 -8601 8921 -8383
rect 8985 -8383 9157 -8041
rect 8985 -8601 8995 -8383
rect 9147 -8601 9157 -8383
rect 9221 -8383 9393 -8041
rect 9221 -8601 9231 -8383
rect 9383 -8601 9393 -8383
rect 9457 -8383 9629 -8041
rect 9457 -8601 9467 -8383
rect 9619 -8601 9629 -8383
rect 9693 -8076 10834 -8041
rect 10890 -8076 10915 -8020
rect 10971 -8076 10996 -8020
rect 11052 -8076 11077 -8020
rect 11133 -8076 11158 -8020
rect 11214 -8076 11239 -8020
rect 11295 -8076 11320 -8020
rect 11376 -8076 11401 -8020
rect 11457 -8076 11482 -8020
rect 11538 -8076 11563 -8020
rect 11619 -8076 11644 -8020
rect 11700 -8076 11725 -8020
rect 11781 -8076 11806 -8020
rect 11862 -8076 11914 -8020
rect 9693 -8124 11914 -8076
rect 9693 -8180 10834 -8124
rect 10890 -8180 10915 -8124
rect 10971 -8180 10996 -8124
rect 11052 -8180 11077 -8124
rect 11133 -8180 11158 -8124
rect 11214 -8180 11239 -8124
rect 11295 -8180 11320 -8124
rect 11376 -8180 11401 -8124
rect 11457 -8180 11482 -8124
rect 11538 -8180 11563 -8124
rect 11619 -8180 11644 -8124
rect 11700 -8180 11725 -8124
rect 11781 -8180 11806 -8124
rect 11862 -8180 11914 -8124
rect 9693 -8228 11914 -8180
rect 9693 -8284 10834 -8228
rect 10890 -8284 10915 -8228
rect 10971 -8284 10996 -8228
rect 11052 -8284 11077 -8228
rect 11133 -8284 11158 -8228
rect 11214 -8284 11239 -8228
rect 11295 -8284 11320 -8228
rect 11376 -8284 11401 -8228
rect 11457 -8284 11482 -8228
rect 11538 -8284 11563 -8228
rect 11619 -8284 11644 -8228
rect 11700 -8284 11725 -8228
rect 11781 -8284 11806 -8228
rect 11862 -8284 11914 -8228
rect 9693 -8332 11914 -8284
rect 9693 -8383 10834 -8332
rect 9693 -8601 9703 -8383
rect 10825 -8388 10834 -8383
rect 10890 -8388 10915 -8332
rect 10971 -8388 10996 -8332
rect 11052 -8388 11077 -8332
rect 11133 -8388 11158 -8332
rect 11214 -8388 11239 -8332
rect 11295 -8388 11320 -8332
rect 11376 -8388 11401 -8332
rect 11457 -8388 11482 -8332
rect 11538 -8388 11563 -8332
rect 11619 -8388 11644 -8332
rect 11700 -8388 11725 -8332
rect 11781 -8388 11806 -8332
rect 11862 -8388 11914 -8332
rect 10825 -8403 11914 -8388
rect 12513 -8059 12523 -7219
rect 12579 -8059 12589 -7219
rect 12513 -8365 12589 -8059
rect 12657 -8054 12667 -7214
rect 12731 -8054 12741 -7214
rect 12657 -8059 12671 -8054
rect 12727 -8059 12741 -8054
rect 12657 -8064 12741 -8059
rect 12809 -7219 12885 -7214
rect 12809 -8059 12819 -7219
rect 12875 -8059 12885 -7219
rect 4044 -9673 5472 -8602
rect 5973 -8606 6049 -8601
rect 6209 -8606 6285 -8601
rect 6445 -8606 6521 -8601
rect 6681 -8606 6757 -8601
rect 6917 -8606 6993 -8601
rect 7153 -8606 7229 -8601
rect 7389 -8606 7465 -8601
rect 7625 -8606 7701 -8601
rect 7971 -8606 8047 -8601
rect 8207 -8606 8283 -8601
rect 8443 -8606 8519 -8601
rect 8679 -8606 8755 -8601
rect 8915 -8606 8991 -8601
rect 9151 -8606 9227 -8601
rect 9387 -8606 9463 -8601
rect 9623 -8606 9699 -8601
rect 12513 -9205 12523 -8365
rect 12579 -9205 12589 -8365
rect 12513 -9673 12589 -9205
rect 12657 -8365 12741 -8360
rect 12657 -8370 12671 -8365
rect 12727 -8370 12741 -8365
rect 12657 -9210 12667 -8370
rect 12731 -9210 12741 -8370
rect 12809 -8365 12885 -8059
rect 12953 -8054 12963 -7214
rect 13027 -8054 13037 -7214
rect 12953 -8059 12967 -8054
rect 13023 -8059 13037 -8054
rect 12953 -8064 13037 -8059
rect 13105 -7219 13181 -7214
rect 13105 -8059 13115 -7219
rect 13171 -8059 13181 -7219
rect 12809 -9205 12819 -8365
rect 12875 -9205 12885 -8365
rect 12809 -9673 12885 -9205
rect 12953 -8365 13037 -8360
rect 12953 -8370 12967 -8365
rect 13023 -8370 13037 -8365
rect 12953 -9210 12963 -8370
rect 13027 -9210 13037 -8370
rect 13105 -8365 13181 -8059
rect 13249 -8054 13259 -7214
rect 13323 -8054 13333 -7214
rect 13249 -8059 13263 -8054
rect 13319 -8059 13333 -8054
rect 13249 -8064 13333 -8059
rect 13401 -7219 13477 -7214
rect 13401 -8059 13411 -7219
rect 13467 -8059 13477 -7219
rect 13105 -9205 13115 -8365
rect 13171 -9205 13181 -8365
rect 13105 -9673 13181 -9205
rect 13249 -8365 13333 -8360
rect 13249 -8370 13263 -8365
rect 13319 -8370 13333 -8365
rect 13249 -9210 13259 -8370
rect 13323 -9210 13333 -8370
rect 13401 -8365 13477 -8059
rect 13545 -8054 13555 -7214
rect 13619 -8054 13629 -7214
rect 13545 -8059 13559 -8054
rect 13615 -8059 13629 -8054
rect 13545 -8064 13629 -8059
rect 13697 -7219 13773 -7214
rect 13697 -8059 13707 -7219
rect 13763 -8059 13773 -7219
rect 13401 -9205 13411 -8365
rect 13467 -9205 13477 -8365
rect 13401 -9673 13477 -9205
rect 13545 -8365 13629 -8360
rect 13545 -8370 13559 -8365
rect 13615 -8370 13629 -8365
rect 13545 -9210 13555 -8370
rect 13619 -9210 13629 -8370
rect 13697 -8365 13773 -8059
rect 13841 -8054 13851 -7214
rect 13915 -8054 13925 -7214
rect 13841 -8059 13855 -8054
rect 13911 -8059 13925 -8054
rect 13841 -8064 13925 -8059
rect 13993 -7219 14069 -7214
rect 13993 -8059 14003 -7219
rect 14059 -8059 14069 -7219
rect 13697 -9205 13707 -8365
rect 13763 -9205 13773 -8365
rect 13697 -9673 13773 -9205
rect 13841 -8365 13925 -8360
rect 13841 -8370 13855 -8365
rect 13911 -8370 13925 -8365
rect 13841 -9210 13851 -8370
rect 13915 -9210 13925 -8370
rect 13993 -8365 14069 -8059
rect 14137 -8054 14147 -7214
rect 14211 -8054 14221 -7214
rect 14137 -8059 14151 -8054
rect 14207 -8059 14221 -8054
rect 14137 -8064 14221 -8059
rect 14289 -7219 14365 -7214
rect 14289 -8059 14299 -7219
rect 14355 -8059 14365 -7219
rect 13993 -9205 14003 -8365
rect 14059 -9205 14069 -8365
rect 13993 -9673 14069 -9205
rect 14137 -8365 14221 -8360
rect 14137 -8370 14151 -8365
rect 14207 -8370 14221 -8365
rect 14137 -9210 14147 -8370
rect 14211 -9210 14221 -8370
rect 14289 -8365 14365 -8059
rect 14433 -8054 14443 -7214
rect 14507 -8054 14517 -7214
rect 14433 -8059 14447 -8054
rect 14503 -8059 14517 -8054
rect 14433 -8064 14517 -8059
rect 14585 -7219 14661 -7214
rect 14585 -8059 14595 -7219
rect 14651 -8059 14661 -7219
rect 14289 -9205 14299 -8365
rect 14355 -9205 14365 -8365
rect 14289 -9673 14365 -9205
rect 14433 -8365 14517 -8360
rect 14433 -8370 14447 -8365
rect 14503 -8370 14517 -8365
rect 14433 -9210 14443 -8370
rect 14507 -9210 14517 -8370
rect 14585 -8365 14661 -8059
rect 14729 -8054 14739 -7214
rect 14803 -8054 14813 -7214
rect 14729 -8059 14743 -8054
rect 14799 -8059 14813 -8054
rect 14729 -8064 14813 -8059
rect 14881 -7219 14957 -7214
rect 14881 -8059 14891 -7219
rect 14947 -8059 14957 -7219
rect 14585 -9205 14595 -8365
rect 14651 -9205 14661 -8365
rect 14585 -9673 14661 -9205
rect 14729 -8365 14813 -8360
rect 14729 -8370 14743 -8365
rect 14799 -8370 14813 -8365
rect 14729 -9210 14739 -8370
rect 14803 -9210 14813 -8370
rect 14881 -8365 14957 -8059
rect 15025 -8054 15035 -7214
rect 15099 -8054 15109 -7214
rect 15025 -8059 15039 -8054
rect 15095 -8059 15109 -8054
rect 15025 -8064 15109 -8059
rect 15177 -7219 15253 -7214
rect 15177 -8059 15187 -7219
rect 15243 -8059 15253 -7219
rect 14881 -9205 14891 -8365
rect 14947 -9205 14957 -8365
rect 14881 -9673 14957 -9205
rect 15025 -8365 15109 -8360
rect 15025 -8370 15039 -8365
rect 15095 -8370 15109 -8365
rect 15025 -9210 15035 -8370
rect 15099 -9210 15109 -8370
rect 15177 -8365 15253 -8059
rect 15321 -8054 15331 -7214
rect 15395 -8054 15405 -7214
rect 15321 -8059 15335 -8054
rect 15391 -8059 15405 -8054
rect 15321 -8064 15405 -8059
rect 15473 -7219 15549 -7214
rect 15473 -8059 15483 -7219
rect 15539 -8059 15549 -7219
rect 15177 -9205 15187 -8365
rect 15243 -9205 15253 -8365
rect 15177 -9673 15253 -9205
rect 15321 -8365 15405 -8360
rect 15321 -8370 15335 -8365
rect 15391 -8370 15405 -8365
rect 15321 -9210 15331 -8370
rect 15395 -9210 15405 -8370
rect 15473 -8365 15549 -8059
rect 15617 -8054 15627 -7214
rect 15691 -8054 15701 -7214
rect 15617 -8059 15631 -8054
rect 15687 -8059 15701 -8054
rect 15617 -8064 15701 -8059
rect 15769 -7219 15845 -7214
rect 15769 -8059 15779 -7219
rect 15835 -8059 15845 -7219
rect 15473 -9205 15483 -8365
rect 15539 -9205 15549 -8365
rect 15473 -9673 15549 -9205
rect 15617 -8365 15701 -8360
rect 15617 -8370 15631 -8365
rect 15687 -8370 15701 -8365
rect 15617 -9210 15627 -8370
rect 15691 -9210 15701 -8370
rect 15769 -8365 15845 -8059
rect 15913 -8054 15923 -7214
rect 15987 -8054 15997 -7214
rect 15913 -8059 15927 -8054
rect 15983 -8059 15997 -8054
rect 15913 -8064 15997 -8059
rect 16065 -7219 16141 -7214
rect 16065 -8059 16075 -7219
rect 16131 -8059 16141 -7219
rect 15769 -9205 15779 -8365
rect 15835 -9205 15845 -8365
rect 15769 -9673 15845 -9205
rect 15913 -8365 15997 -8360
rect 15913 -8370 15927 -8365
rect 15983 -8370 15997 -8365
rect 15913 -9210 15923 -8370
rect 15987 -9210 15997 -8370
rect 16065 -8365 16141 -8059
rect 16209 -8054 16219 -7214
rect 16283 -8054 16293 -7214
rect 16209 -8059 16223 -8054
rect 16279 -8059 16293 -8054
rect 16209 -8064 16293 -8059
rect 16361 -7219 16437 -7214
rect 16361 -8059 16371 -7219
rect 16427 -8059 16437 -7219
rect 16065 -9205 16075 -8365
rect 16131 -9205 16141 -8365
rect 16065 -9673 16141 -9205
rect 16209 -8365 16293 -8360
rect 16209 -8370 16223 -8365
rect 16279 -8370 16293 -8365
rect 16209 -9210 16219 -8370
rect 16283 -9210 16293 -8370
rect 16361 -8365 16437 -8059
rect 16505 -8054 16515 -7214
rect 16579 -8054 16589 -7214
rect 16505 -8059 16519 -8054
rect 16575 -8059 16589 -8054
rect 16505 -8064 16589 -8059
rect 16657 -7219 16733 -7214
rect 16657 -8059 16667 -7219
rect 16723 -8059 16733 -7219
rect 16361 -9205 16371 -8365
rect 16427 -9205 16437 -8365
rect 16361 -9673 16437 -9205
rect 16505 -8365 16589 -8360
rect 16505 -8370 16519 -8365
rect 16575 -8370 16589 -8365
rect 16505 -9210 16515 -8370
rect 16579 -9210 16589 -8370
rect 16657 -8365 16733 -8059
rect 16801 -8054 16811 -7214
rect 16875 -8054 16885 -7214
rect 16801 -8059 16815 -8054
rect 16871 -8059 16885 -8054
rect 16801 -8064 16885 -8059
rect 16953 -7219 17029 -7214
rect 16953 -8059 16963 -7219
rect 17019 -8059 17029 -7219
rect 16657 -9205 16667 -8365
rect 16723 -9205 16733 -8365
rect 16657 -9673 16733 -9205
rect 16801 -8365 16885 -8360
rect 16801 -8370 16815 -8365
rect 16871 -8370 16885 -8365
rect 16801 -9210 16811 -8370
rect 16875 -9210 16885 -8370
rect 16953 -8365 17029 -8059
rect 17097 -8054 17107 -7214
rect 17171 -8054 17181 -7214
rect 17097 -8059 17111 -8054
rect 17167 -8059 17181 -8054
rect 17097 -8064 17181 -8059
rect 17249 -7219 17325 -7214
rect 17249 -8059 17259 -7219
rect 17315 -8059 17325 -7219
rect 16953 -9205 16963 -8365
rect 17019 -9205 17029 -8365
rect 16953 -9673 17029 -9205
rect 17097 -8365 17181 -8360
rect 17097 -8370 17111 -8365
rect 17167 -8370 17181 -8365
rect 17097 -9210 17107 -8370
rect 17171 -9210 17181 -8370
rect 17249 -8365 17325 -8059
rect 17393 -8054 17403 -7214
rect 17467 -8054 17477 -7214
rect 17393 -8059 17407 -8054
rect 17463 -8059 17477 -8054
rect 17393 -8064 17477 -8059
rect 17545 -7219 17621 -7214
rect 17545 -8059 17555 -7219
rect 17611 -8059 17621 -7219
rect 17249 -9205 17259 -8365
rect 17315 -9205 17325 -8365
rect 17249 -9673 17325 -9205
rect 17393 -8365 17477 -8360
rect 17393 -8370 17407 -8365
rect 17463 -8370 17477 -8365
rect 17393 -9210 17403 -8370
rect 17467 -9210 17477 -8370
rect 17545 -8365 17621 -8059
rect 17689 -8054 17699 -7214
rect 17763 -8054 17773 -7214
rect 17689 -8059 17703 -8054
rect 17759 -8059 17773 -8054
rect 17689 -8064 17773 -8059
rect 17841 -7219 17917 -7214
rect 17841 -8059 17851 -7219
rect 17907 -8059 17917 -7219
rect 17545 -9205 17555 -8365
rect 17611 -9205 17621 -8365
rect 17545 -9673 17621 -9205
rect 17689 -8365 17773 -8360
rect 17689 -8370 17703 -8365
rect 17759 -8370 17773 -8365
rect 17689 -9210 17699 -8370
rect 17763 -9210 17773 -8370
rect 17841 -8365 17917 -8059
rect 17985 -8054 17995 -7214
rect 18059 -8054 18069 -7214
rect 17985 -8059 17999 -8054
rect 18055 -8059 18069 -8054
rect 17985 -8064 18069 -8059
rect 18137 -7219 18213 -7214
rect 18137 -8059 18147 -7219
rect 18203 -8059 18213 -7219
rect 17841 -9205 17851 -8365
rect 17907 -9205 17917 -8365
rect 17841 -9673 17917 -9205
rect 17985 -8365 18069 -8360
rect 17985 -8370 17999 -8365
rect 18055 -8370 18069 -8365
rect 17985 -9210 17995 -8370
rect 18059 -9210 18069 -8370
rect 18137 -8365 18213 -8059
rect 18281 -8054 18291 -7214
rect 18355 -8054 18365 -7214
rect 18281 -8059 18295 -8054
rect 18351 -8059 18365 -8054
rect 18281 -8064 18365 -8059
rect 18433 -7219 18509 -7214
rect 18433 -8059 18443 -7219
rect 18499 -8059 18509 -7219
rect 18137 -9205 18147 -8365
rect 18203 -9205 18213 -8365
rect 18137 -9673 18213 -9205
rect 18281 -8365 18365 -8360
rect 18281 -8370 18295 -8365
rect 18351 -8370 18365 -8365
rect 18281 -9210 18291 -8370
rect 18355 -9210 18365 -8370
rect 18433 -8365 18509 -8059
rect 18577 -8054 18587 -7214
rect 18651 -8054 18661 -7214
rect 18577 -8059 18591 -8054
rect 18647 -8059 18661 -8054
rect 18577 -8064 18661 -8059
rect 18729 -7219 18805 -7214
rect 18729 -8059 18739 -7219
rect 18795 -8059 18805 -7219
rect 18433 -9205 18443 -8365
rect 18499 -9205 18509 -8365
rect 18433 -9673 18509 -9205
rect 18577 -8365 18661 -8360
rect 18577 -8370 18591 -8365
rect 18647 -8370 18661 -8365
rect 18577 -9210 18587 -8370
rect 18651 -9210 18661 -8370
rect 18729 -8365 18805 -8059
rect 18873 -8054 18883 -7214
rect 18947 -8054 18957 -7214
rect 18873 -8059 18887 -8054
rect 18943 -8059 18957 -8054
rect 18873 -8064 18957 -8059
rect 19025 -7219 19101 -7214
rect 19025 -8059 19035 -7219
rect 19091 -8059 19101 -7219
rect 18729 -9205 18739 -8365
rect 18795 -9205 18805 -8365
rect 18729 -9673 18805 -9205
rect 18873 -8365 18957 -8360
rect 18873 -8370 18887 -8365
rect 18943 -8370 18957 -8365
rect 18873 -9210 18883 -8370
rect 18947 -9210 18957 -8370
rect 19025 -8365 19101 -8059
rect 19169 -8054 19179 -7214
rect 19243 -8054 19253 -7214
rect 19169 -8059 19183 -8054
rect 19239 -8059 19253 -8054
rect 19169 -8064 19253 -8059
rect 19321 -7219 19397 -7214
rect 19321 -8059 19331 -7219
rect 19387 -8059 19397 -7219
rect 19025 -9205 19035 -8365
rect 19091 -9205 19101 -8365
rect 19025 -9673 19101 -9205
rect 19169 -8365 19253 -8360
rect 19169 -8370 19183 -8365
rect 19239 -8370 19253 -8365
rect 19169 -9210 19179 -8370
rect 19243 -9210 19253 -8370
rect 19321 -8365 19397 -8059
rect 19465 -8054 19475 -7214
rect 19539 -8054 19549 -7214
rect 19465 -8059 19479 -8054
rect 19535 -8059 19549 -8054
rect 19465 -8064 19549 -8059
rect 19617 -7219 19693 -7214
rect 19617 -8059 19627 -7219
rect 19683 -8059 19693 -7219
rect 19321 -9205 19331 -8365
rect 19387 -9205 19397 -8365
rect 19321 -9673 19397 -9205
rect 19465 -8365 19549 -8360
rect 19465 -8370 19479 -8365
rect 19535 -8370 19549 -8365
rect 19465 -9210 19475 -8370
rect 19539 -9210 19549 -8370
rect 19617 -8365 19693 -8059
rect 19761 -8054 19771 -7214
rect 19835 -8054 19845 -7214
rect 19761 -8059 19775 -8054
rect 19831 -8059 19845 -8054
rect 19761 -8064 19845 -8059
rect 19913 -7219 19989 -7214
rect 19913 -8059 19923 -7219
rect 19979 -8059 19989 -7219
rect 19617 -9205 19627 -8365
rect 19683 -9205 19693 -8365
rect 19617 -9673 19693 -9205
rect 19761 -8365 19845 -8360
rect 19761 -8370 19775 -8365
rect 19831 -8370 19845 -8365
rect 19761 -9210 19771 -8370
rect 19835 -9210 19845 -8370
rect 19913 -8365 19989 -8059
rect 20057 -8054 20067 -7214
rect 20131 -8054 20141 -7214
rect 20057 -8059 20071 -8054
rect 20127 -8059 20141 -8054
rect 20057 -8064 20141 -8059
rect 20209 -7219 20285 -7214
rect 20209 -8059 20219 -7219
rect 20275 -8059 20285 -7219
rect 19913 -9205 19923 -8365
rect 19979 -9205 19989 -8365
rect 19913 -9673 19989 -9205
rect 20057 -8365 20141 -8360
rect 20057 -8370 20071 -8365
rect 20127 -8370 20141 -8365
rect 20057 -9210 20067 -8370
rect 20131 -9210 20141 -8370
rect 20209 -8365 20285 -8059
rect 20353 -8054 20363 -7214
rect 20427 -8054 20437 -7214
rect 20353 -8059 20367 -8054
rect 20423 -8059 20437 -8054
rect 20353 -8064 20437 -8059
rect 20505 -7219 20581 -7214
rect 20505 -8059 20515 -7219
rect 20571 -8059 20581 -7219
rect 20209 -9205 20219 -8365
rect 20275 -9205 20285 -8365
rect 20209 -9673 20285 -9205
rect 20353 -8365 20437 -8360
rect 20353 -8370 20367 -8365
rect 20423 -8370 20437 -8365
rect 20353 -9210 20363 -8370
rect 20427 -9210 20437 -8370
rect 20505 -8365 20581 -8059
rect 20649 -8054 20659 -7214
rect 20723 -8054 20733 -7214
rect 20649 -8059 20663 -8054
rect 20719 -8059 20733 -8054
rect 20649 -8064 20733 -8059
rect 20801 -7219 20877 -7214
rect 20801 -8059 20811 -7219
rect 20867 -8059 20877 -7219
rect 20505 -9205 20515 -8365
rect 20571 -9205 20581 -8365
rect 20505 -9673 20581 -9205
rect 20649 -8365 20733 -8360
rect 20649 -8370 20663 -8365
rect 20719 -8370 20733 -8365
rect 20649 -9210 20659 -8370
rect 20723 -9210 20733 -8370
rect 20801 -8365 20877 -8059
rect 20945 -8054 20955 -7214
rect 21019 -8054 21029 -7214
rect 20945 -8059 20959 -8054
rect 21015 -8059 21029 -8054
rect 20945 -8064 21029 -8059
rect 21097 -7219 21173 -7214
rect 21097 -8059 21107 -7219
rect 21163 -8059 21173 -7219
rect 20801 -9205 20811 -8365
rect 20867 -9205 20877 -8365
rect 20801 -9673 20877 -9205
rect 20945 -8365 21029 -8360
rect 20945 -8370 20959 -8365
rect 21015 -8370 21029 -8365
rect 20945 -9210 20955 -8370
rect 21019 -9210 21029 -8370
rect 21097 -8365 21173 -8059
rect 21241 -8054 21251 -7214
rect 21315 -8054 21325 -7214
rect 21241 -8059 21255 -8054
rect 21311 -8059 21325 -8054
rect 21241 -8064 21325 -8059
rect 21393 -7219 21469 -7214
rect 21393 -8059 21403 -7219
rect 21459 -8059 21469 -7219
rect 21097 -9205 21107 -8365
rect 21163 -9205 21173 -8365
rect 21097 -9673 21173 -9205
rect 21241 -8365 21325 -8360
rect 21241 -8370 21255 -8365
rect 21311 -8370 21325 -8365
rect 21241 -9210 21251 -8370
rect 21315 -9210 21325 -8370
rect 21393 -8365 21469 -8059
rect 21537 -8054 21547 -7214
rect 21611 -8054 21621 -7214
rect 21537 -8059 21551 -8054
rect 21607 -8059 21621 -8054
rect 21537 -8064 21621 -8059
rect 21689 -7219 21765 -7214
rect 21689 -8059 21699 -7219
rect 21755 -8059 21765 -7219
rect 21393 -9205 21403 -8365
rect 21459 -9205 21469 -8365
rect 21393 -9673 21469 -9205
rect 21537 -8365 21621 -8360
rect 21537 -8370 21551 -8365
rect 21607 -8370 21621 -8365
rect 21537 -9210 21547 -8370
rect 21611 -9210 21621 -8370
rect 21689 -8365 21765 -8059
rect 21833 -8054 21843 -7214
rect 21907 -8054 21917 -7214
rect 21833 -8059 21847 -8054
rect 21903 -8059 21917 -8054
rect 21833 -8064 21917 -8059
rect 21985 -7219 22061 -7214
rect 21985 -8059 21995 -7219
rect 22051 -8059 22061 -7219
rect 21689 -9205 21699 -8365
rect 21755 -9205 21765 -8365
rect 21689 -9673 21765 -9205
rect 21833 -8365 21917 -8360
rect 21833 -8370 21847 -8365
rect 21903 -8370 21917 -8365
rect 21833 -9210 21843 -8370
rect 21907 -9210 21917 -8370
rect 21985 -8365 22061 -8059
rect 22129 -8054 22139 -7214
rect 22203 -8054 22213 -7214
rect 22129 -8059 22143 -8054
rect 22199 -8059 22213 -8054
rect 22129 -8064 22213 -8059
rect 22281 -7219 22357 -7214
rect 22281 -8059 22291 -7219
rect 22347 -8059 22357 -7219
rect 21985 -9205 21995 -8365
rect 22051 -9205 22061 -8365
rect 21985 -9673 22061 -9205
rect 22129 -8365 22213 -8360
rect 22129 -8370 22143 -8365
rect 22199 -8370 22213 -8365
rect 22129 -9210 22139 -8370
rect 22203 -9210 22213 -8370
rect 22281 -8365 22357 -8059
rect 22425 -8054 22435 -7214
rect 22499 -8054 22509 -7214
rect 22425 -8059 22439 -8054
rect 22495 -8059 22509 -8054
rect 22425 -8064 22509 -8059
rect 22577 -7219 22653 -7214
rect 22577 -8059 22587 -7219
rect 22643 -8059 22653 -7219
rect 22281 -9205 22291 -8365
rect 22347 -9205 22357 -8365
rect 22281 -9673 22357 -9205
rect 22425 -8365 22509 -8360
rect 22425 -8370 22439 -8365
rect 22495 -8370 22509 -8365
rect 22425 -9210 22435 -8370
rect 22499 -9210 22509 -8370
rect 22577 -8365 22653 -8059
rect 22721 -8054 22731 -7214
rect 22795 -8054 22805 -7214
rect 22721 -8059 22735 -8054
rect 22791 -8059 22805 -8054
rect 22721 -8064 22805 -8059
rect 22873 -7219 22949 -7214
rect 22873 -8059 22883 -7219
rect 22939 -8059 22949 -7219
rect 22577 -9205 22587 -8365
rect 22643 -9205 22653 -8365
rect 22577 -9673 22653 -9205
rect 22721 -8365 22805 -8360
rect 22721 -8370 22735 -8365
rect 22791 -8370 22805 -8365
rect 22721 -9210 22731 -8370
rect 22795 -9210 22805 -8370
rect 22873 -8365 22949 -8059
rect 23017 -8054 23027 -7214
rect 23091 -8054 23101 -7214
rect 23017 -8059 23031 -8054
rect 23087 -8059 23101 -8054
rect 23017 -8064 23101 -8059
rect 23169 -7219 23245 -7214
rect 23169 -8059 23179 -7219
rect 23235 -8059 23245 -7219
rect 22873 -9205 22883 -8365
rect 22939 -9205 22949 -8365
rect 22873 -9673 22949 -9205
rect 23017 -8365 23101 -8360
rect 23017 -8370 23031 -8365
rect 23087 -8370 23101 -8365
rect 23017 -9210 23027 -8370
rect 23091 -9210 23101 -8370
rect 23169 -8365 23245 -8059
rect 23313 -8054 23323 -7214
rect 23387 -8054 23397 -7214
rect 23313 -8059 23327 -8054
rect 23383 -8059 23397 -8054
rect 23313 -8064 23397 -8059
rect 23465 -7219 23541 -7214
rect 23465 -8059 23475 -7219
rect 23531 -8059 23541 -7219
rect 23169 -9205 23179 -8365
rect 23235 -9205 23245 -8365
rect 23169 -9673 23245 -9205
rect 23313 -8365 23397 -8360
rect 23313 -8370 23327 -8365
rect 23383 -8370 23397 -8365
rect 23313 -9210 23323 -8370
rect 23387 -9210 23397 -8370
rect 23465 -8365 23541 -8059
rect 23609 -8054 23619 -7214
rect 23683 -8054 23693 -7214
rect 23609 -8059 23623 -8054
rect 23679 -8059 23693 -8054
rect 23609 -8064 23693 -8059
rect 23465 -9205 23475 -8365
rect 23531 -9205 23541 -8365
rect 23465 -9673 23541 -9205
rect 23609 -8365 23693 -8360
rect 23609 -8370 23623 -8365
rect 23679 -8370 23693 -8365
rect 23609 -9210 23619 -8370
rect 23683 -9210 23693 -8370
rect 4044 -9681 26275 -9673
rect 4044 -9737 4053 -9681
rect 4109 -9737 4134 -9681
rect 4190 -9737 4215 -9681
rect 4271 -9737 4296 -9681
rect 4352 -9737 4377 -9681
rect 4433 -9737 4458 -9681
rect 4514 -9737 4539 -9681
rect 4595 -9737 4621 -9681
rect 4677 -9737 4702 -9681
rect 4758 -9737 4783 -9681
rect 4839 -9737 4864 -9681
rect 4920 -9737 4945 -9681
rect 5001 -9737 5026 -9681
rect 5082 -9737 5107 -9681
rect 5163 -9737 5189 -9681
rect 5245 -9737 5270 -9681
rect 5326 -9737 5351 -9681
rect 5407 -9737 5432 -9681
rect 5488 -9737 5513 -9681
rect 5569 -9737 5594 -9681
rect 5650 -9737 5675 -9681
rect 5731 -9737 5757 -9681
rect 5813 -9737 5838 -9681
rect 5894 -9737 5919 -9681
rect 5975 -9737 6000 -9681
rect 6056 -9737 6081 -9681
rect 6137 -9737 6162 -9681
rect 6218 -9737 6243 -9681
rect 6299 -9737 6325 -9681
rect 6381 -9737 6406 -9681
rect 6462 -9737 6487 -9681
rect 6543 -9737 6568 -9681
rect 6624 -9737 6649 -9681
rect 6705 -9737 6730 -9681
rect 6786 -9737 6811 -9681
rect 6867 -9737 6893 -9681
rect 6949 -9737 6974 -9681
rect 7030 -9737 7055 -9681
rect 7111 -9737 7136 -9681
rect 7192 -9737 7217 -9681
rect 7273 -9737 7298 -9681
rect 7354 -9737 7379 -9681
rect 7435 -9737 7461 -9681
rect 7517 -9737 7542 -9681
rect 7598 -9737 7623 -9681
rect 7679 -9737 7704 -9681
rect 7760 -9737 7785 -9681
rect 7841 -9737 7866 -9681
rect 7922 -9737 7947 -9681
rect 8003 -9737 8029 -9681
rect 8085 -9737 8110 -9681
rect 8166 -9737 8191 -9681
rect 8247 -9737 8272 -9681
rect 8328 -9737 8353 -9681
rect 8409 -9737 8434 -9681
rect 8490 -9737 8515 -9681
rect 8571 -9737 8597 -9681
rect 8653 -9737 8678 -9681
rect 8734 -9737 8759 -9681
rect 8815 -9737 8840 -9681
rect 8896 -9737 8921 -9681
rect 8977 -9737 9002 -9681
rect 9058 -9737 9083 -9681
rect 9139 -9737 9165 -9681
rect 9221 -9737 9246 -9681
rect 9302 -9737 9327 -9681
rect 9383 -9737 9408 -9681
rect 9464 -9737 9489 -9681
rect 9545 -9737 9570 -9681
rect 9626 -9737 9651 -9681
rect 9707 -9737 9733 -9681
rect 9789 -9737 9814 -9681
rect 9870 -9737 9895 -9681
rect 9951 -9737 9976 -9681
rect 10032 -9737 10057 -9681
rect 10113 -9737 10138 -9681
rect 10194 -9737 10219 -9681
rect 10275 -9737 10301 -9681
rect 10357 -9737 10382 -9681
rect 10438 -9737 10463 -9681
rect 10519 -9737 10544 -9681
rect 10600 -9737 10625 -9681
rect 10681 -9737 10706 -9681
rect 10762 -9737 10787 -9681
rect 10843 -9737 10869 -9681
rect 10925 -9737 10950 -9681
rect 11006 -9737 11031 -9681
rect 11087 -9737 11112 -9681
rect 11168 -9737 11193 -9681
rect 11249 -9737 11274 -9681
rect 11330 -9737 11355 -9681
rect 11411 -9737 11437 -9681
rect 11493 -9737 11518 -9681
rect 11574 -9737 11599 -9681
rect 11655 -9737 11680 -9681
rect 11736 -9737 11761 -9681
rect 11817 -9737 11842 -9681
rect 11898 -9737 11923 -9681
rect 11979 -9737 12005 -9681
rect 12061 -9737 12086 -9681
rect 12142 -9737 12167 -9681
rect 12223 -9737 12248 -9681
rect 12304 -9737 12329 -9681
rect 12385 -9737 12410 -9681
rect 12466 -9737 12491 -9681
rect 12547 -9737 12573 -9681
rect 12629 -9737 12654 -9681
rect 12710 -9737 12735 -9681
rect 12791 -9737 12816 -9681
rect 12872 -9737 12897 -9681
rect 12953 -9737 12978 -9681
rect 13034 -9737 13059 -9681
rect 13115 -9737 13141 -9681
rect 13197 -9737 13222 -9681
rect 13278 -9737 13303 -9681
rect 13359 -9737 13384 -9681
rect 13440 -9737 13465 -9681
rect 13521 -9737 13546 -9681
rect 13602 -9737 13627 -9681
rect 13683 -9737 13709 -9681
rect 13765 -9737 13790 -9681
rect 13846 -9737 13871 -9681
rect 13927 -9737 13952 -9681
rect 14008 -9737 14033 -9681
rect 14089 -9737 14114 -9681
rect 14170 -9737 14195 -9681
rect 14251 -9737 14277 -9681
rect 14333 -9737 14358 -9681
rect 14414 -9737 14439 -9681
rect 14495 -9737 14520 -9681
rect 14576 -9737 14601 -9681
rect 14657 -9737 14682 -9681
rect 14738 -9737 14763 -9681
rect 14819 -9737 14845 -9681
rect 14901 -9737 14926 -9681
rect 14982 -9737 15007 -9681
rect 15063 -9737 15088 -9681
rect 15144 -9737 15169 -9681
rect 15225 -9737 15250 -9681
rect 15306 -9737 15331 -9681
rect 15387 -9737 15413 -9681
rect 15469 -9737 15494 -9681
rect 15550 -9737 15575 -9681
rect 15631 -9737 15656 -9681
rect 15712 -9737 15737 -9681
rect 15793 -9737 15818 -9681
rect 15874 -9737 15899 -9681
rect 15955 -9737 15981 -9681
rect 16037 -9737 16062 -9681
rect 16118 -9737 16143 -9681
rect 16199 -9737 16224 -9681
rect 16280 -9737 16305 -9681
rect 16361 -9737 16386 -9681
rect 16442 -9737 16467 -9681
rect 16523 -9737 16549 -9681
rect 16605 -9737 16630 -9681
rect 16686 -9737 16711 -9681
rect 16767 -9737 16792 -9681
rect 16848 -9737 16873 -9681
rect 16929 -9737 16954 -9681
rect 17010 -9737 17035 -9681
rect 17091 -9737 17117 -9681
rect 17173 -9737 17198 -9681
rect 17254 -9737 17279 -9681
rect 17335 -9737 17360 -9681
rect 17416 -9737 17441 -9681
rect 17497 -9737 17522 -9681
rect 17578 -9737 17603 -9681
rect 17659 -9737 17684 -9681
rect 17740 -9737 17765 -9681
rect 17821 -9737 17846 -9681
rect 17902 -9737 17927 -9681
rect 17983 -9737 18008 -9681
rect 18064 -9737 18089 -9681
rect 18145 -9737 18171 -9681
rect 18227 -9737 18252 -9681
rect 18308 -9737 18333 -9681
rect 18389 -9737 18414 -9681
rect 18470 -9737 18495 -9681
rect 18551 -9737 18576 -9681
rect 18632 -9737 18657 -9681
rect 18713 -9737 18739 -9681
rect 18795 -9737 18820 -9681
rect 18876 -9737 18901 -9681
rect 18957 -9737 18982 -9681
rect 19038 -9737 19063 -9681
rect 19119 -9737 19144 -9681
rect 19200 -9737 19225 -9681
rect 19281 -9737 19307 -9681
rect 19363 -9737 19388 -9681
rect 19444 -9737 19469 -9681
rect 19525 -9737 19550 -9681
rect 19606 -9737 19631 -9681
rect 19687 -9737 19712 -9681
rect 19768 -9737 19793 -9681
rect 19849 -9737 19875 -9681
rect 19931 -9737 19956 -9681
rect 20012 -9737 20037 -9681
rect 20093 -9737 20118 -9681
rect 20174 -9737 20199 -9681
rect 20255 -9737 20280 -9681
rect 20336 -9737 20361 -9681
rect 20417 -9737 20443 -9681
rect 20499 -9737 20524 -9681
rect 20580 -9737 20605 -9681
rect 20661 -9737 20686 -9681
rect 20742 -9737 20767 -9681
rect 20823 -9737 20848 -9681
rect 20904 -9737 20929 -9681
rect 20985 -9737 21011 -9681
rect 21067 -9737 21092 -9681
rect 21148 -9737 21173 -9681
rect 21229 -9737 21254 -9681
rect 21310 -9737 21335 -9681
rect 21391 -9737 21416 -9681
rect 21472 -9737 21497 -9681
rect 21553 -9737 21579 -9681
rect 21635 -9737 21660 -9681
rect 21716 -9737 21741 -9681
rect 21797 -9737 21822 -9681
rect 21878 -9737 21903 -9681
rect 21959 -9737 21984 -9681
rect 22040 -9737 22065 -9681
rect 22121 -9737 22147 -9681
rect 22203 -9737 22228 -9681
rect 22284 -9737 22309 -9681
rect 22365 -9737 22390 -9681
rect 22446 -9737 22471 -9681
rect 22527 -9737 22552 -9681
rect 22608 -9737 22633 -9681
rect 22689 -9737 22715 -9681
rect 22771 -9737 22796 -9681
rect 22852 -9737 22877 -9681
rect 22933 -9737 22958 -9681
rect 23014 -9737 23039 -9681
rect 23095 -9737 23120 -9681
rect 23176 -9737 23201 -9681
rect 23257 -9737 23283 -9681
rect 23339 -9737 23364 -9681
rect 23420 -9737 23445 -9681
rect 23501 -9737 23526 -9681
rect 23582 -9737 23607 -9681
rect 23663 -9737 23688 -9681
rect 23744 -9737 23769 -9681
rect 23825 -9737 23851 -9681
rect 23907 -9737 23932 -9681
rect 23988 -9737 24013 -9681
rect 24069 -9737 24094 -9681
rect 24150 -9737 24175 -9681
rect 24231 -9737 24256 -9681
rect 24312 -9737 24337 -9681
rect 24393 -9737 24419 -9681
rect 24475 -9737 24500 -9681
rect 24556 -9737 24581 -9681
rect 24637 -9737 24662 -9681
rect 24718 -9737 24743 -9681
rect 24799 -9737 24824 -9681
rect 24880 -9737 24905 -9681
rect 24961 -9737 24987 -9681
rect 25043 -9737 25068 -9681
rect 25124 -9737 25149 -9681
rect 25205 -9737 25230 -9681
rect 25286 -9737 25311 -9681
rect 25367 -9737 25392 -9681
rect 25448 -9737 25473 -9681
rect 25529 -9737 25555 -9681
rect 25611 -9737 25636 -9681
rect 25692 -9737 25717 -9681
rect 25773 -9737 25798 -9681
rect 25854 -9737 25879 -9681
rect 25935 -9737 25960 -9681
rect 26016 -9737 26041 -9681
rect 26097 -9737 26123 -9681
rect 26179 -9737 26204 -9681
rect 26260 -9737 26275 -9681
rect 4044 -9785 26275 -9737
rect 4044 -9841 4053 -9785
rect 4109 -9841 4134 -9785
rect 4190 -9841 4215 -9785
rect 4271 -9841 4296 -9785
rect 4352 -9841 4377 -9785
rect 4433 -9841 4458 -9785
rect 4514 -9841 4539 -9785
rect 4595 -9841 4621 -9785
rect 4677 -9841 4702 -9785
rect 4758 -9841 4783 -9785
rect 4839 -9841 4864 -9785
rect 4920 -9841 4945 -9785
rect 5001 -9841 5026 -9785
rect 5082 -9841 5107 -9785
rect 5163 -9841 5189 -9785
rect 5245 -9841 5270 -9785
rect 5326 -9841 5351 -9785
rect 5407 -9841 5432 -9785
rect 5488 -9841 5513 -9785
rect 5569 -9841 5594 -9785
rect 5650 -9841 5675 -9785
rect 5731 -9841 5757 -9785
rect 5813 -9841 5838 -9785
rect 5894 -9841 5919 -9785
rect 5975 -9841 6000 -9785
rect 6056 -9841 6081 -9785
rect 6137 -9841 6162 -9785
rect 6218 -9841 6243 -9785
rect 6299 -9841 6325 -9785
rect 6381 -9841 6406 -9785
rect 6462 -9841 6487 -9785
rect 6543 -9841 6568 -9785
rect 6624 -9841 6649 -9785
rect 6705 -9841 6730 -9785
rect 6786 -9841 6811 -9785
rect 6867 -9841 6893 -9785
rect 6949 -9841 6974 -9785
rect 7030 -9841 7055 -9785
rect 7111 -9841 7136 -9785
rect 7192 -9841 7217 -9785
rect 7273 -9841 7298 -9785
rect 7354 -9841 7379 -9785
rect 7435 -9841 7461 -9785
rect 7517 -9841 7542 -9785
rect 7598 -9841 7623 -9785
rect 7679 -9841 7704 -9785
rect 7760 -9841 7785 -9785
rect 7841 -9841 7866 -9785
rect 7922 -9841 7947 -9785
rect 8003 -9841 8029 -9785
rect 8085 -9841 8110 -9785
rect 8166 -9841 8191 -9785
rect 8247 -9841 8272 -9785
rect 8328 -9841 8353 -9785
rect 8409 -9841 8434 -9785
rect 8490 -9841 8515 -9785
rect 8571 -9841 8597 -9785
rect 8653 -9841 8678 -9785
rect 8734 -9841 8759 -9785
rect 8815 -9841 8840 -9785
rect 8896 -9841 8921 -9785
rect 8977 -9841 9002 -9785
rect 9058 -9841 9083 -9785
rect 9139 -9841 9165 -9785
rect 9221 -9841 9246 -9785
rect 9302 -9841 9327 -9785
rect 9383 -9841 9408 -9785
rect 9464 -9841 9489 -9785
rect 9545 -9841 9570 -9785
rect 9626 -9841 9651 -9785
rect 9707 -9841 9733 -9785
rect 9789 -9841 9814 -9785
rect 9870 -9841 9895 -9785
rect 9951 -9841 9976 -9785
rect 10032 -9841 10057 -9785
rect 10113 -9841 10138 -9785
rect 10194 -9841 10219 -9785
rect 10275 -9841 10301 -9785
rect 10357 -9841 10382 -9785
rect 10438 -9841 10463 -9785
rect 10519 -9841 10544 -9785
rect 10600 -9841 10625 -9785
rect 10681 -9841 10706 -9785
rect 10762 -9841 10787 -9785
rect 10843 -9841 10869 -9785
rect 10925 -9841 10950 -9785
rect 11006 -9841 11031 -9785
rect 11087 -9841 11112 -9785
rect 11168 -9841 11193 -9785
rect 11249 -9841 11274 -9785
rect 11330 -9841 11355 -9785
rect 11411 -9841 11437 -9785
rect 11493 -9841 11518 -9785
rect 11574 -9841 11599 -9785
rect 11655 -9841 11680 -9785
rect 11736 -9841 11761 -9785
rect 11817 -9841 11842 -9785
rect 11898 -9841 11923 -9785
rect 11979 -9841 12005 -9785
rect 12061 -9841 12086 -9785
rect 12142 -9841 12167 -9785
rect 12223 -9841 12248 -9785
rect 12304 -9841 12329 -9785
rect 12385 -9841 12410 -9785
rect 12466 -9841 12491 -9785
rect 12547 -9841 12573 -9785
rect 12629 -9841 12654 -9785
rect 12710 -9841 12735 -9785
rect 12791 -9841 12816 -9785
rect 12872 -9841 12897 -9785
rect 12953 -9841 12978 -9785
rect 13034 -9841 13059 -9785
rect 13115 -9841 13141 -9785
rect 13197 -9841 13222 -9785
rect 13278 -9841 13303 -9785
rect 13359 -9841 13384 -9785
rect 13440 -9841 13465 -9785
rect 13521 -9841 13546 -9785
rect 13602 -9841 13627 -9785
rect 13683 -9841 13709 -9785
rect 13765 -9841 13790 -9785
rect 13846 -9841 13871 -9785
rect 13927 -9841 13952 -9785
rect 14008 -9841 14033 -9785
rect 14089 -9841 14114 -9785
rect 14170 -9841 14195 -9785
rect 14251 -9841 14277 -9785
rect 14333 -9841 14358 -9785
rect 14414 -9841 14439 -9785
rect 14495 -9841 14520 -9785
rect 14576 -9841 14601 -9785
rect 14657 -9841 14682 -9785
rect 14738 -9841 14763 -9785
rect 14819 -9841 14845 -9785
rect 14901 -9841 14926 -9785
rect 14982 -9841 15007 -9785
rect 15063 -9841 15088 -9785
rect 15144 -9841 15169 -9785
rect 15225 -9841 15250 -9785
rect 15306 -9841 15331 -9785
rect 15387 -9841 15413 -9785
rect 15469 -9841 15494 -9785
rect 15550 -9841 15575 -9785
rect 15631 -9841 15656 -9785
rect 15712 -9841 15737 -9785
rect 15793 -9841 15818 -9785
rect 15874 -9841 15899 -9785
rect 15955 -9841 15981 -9785
rect 16037 -9841 16062 -9785
rect 16118 -9841 16143 -9785
rect 16199 -9841 16224 -9785
rect 16280 -9841 16305 -9785
rect 16361 -9841 16386 -9785
rect 16442 -9841 16467 -9785
rect 16523 -9841 16549 -9785
rect 16605 -9841 16630 -9785
rect 16686 -9841 16711 -9785
rect 16767 -9841 16792 -9785
rect 16848 -9841 16873 -9785
rect 16929 -9841 16954 -9785
rect 17010 -9841 17035 -9785
rect 17091 -9841 17117 -9785
rect 17173 -9841 17198 -9785
rect 17254 -9841 17279 -9785
rect 17335 -9841 17360 -9785
rect 17416 -9841 17441 -9785
rect 17497 -9841 17522 -9785
rect 17578 -9841 17603 -9785
rect 17659 -9841 17684 -9785
rect 17740 -9841 17765 -9785
rect 17821 -9841 17846 -9785
rect 17902 -9841 17927 -9785
rect 17983 -9841 18008 -9785
rect 18064 -9841 18089 -9785
rect 18145 -9841 18171 -9785
rect 18227 -9841 18252 -9785
rect 18308 -9841 18333 -9785
rect 18389 -9841 18414 -9785
rect 18470 -9841 18495 -9785
rect 18551 -9841 18576 -9785
rect 18632 -9841 18657 -9785
rect 18713 -9841 18739 -9785
rect 18795 -9841 18820 -9785
rect 18876 -9841 18901 -9785
rect 18957 -9841 18982 -9785
rect 19038 -9841 19063 -9785
rect 19119 -9841 19144 -9785
rect 19200 -9841 19225 -9785
rect 19281 -9841 19307 -9785
rect 19363 -9841 19388 -9785
rect 19444 -9841 19469 -9785
rect 19525 -9841 19550 -9785
rect 19606 -9841 19631 -9785
rect 19687 -9841 19712 -9785
rect 19768 -9841 19793 -9785
rect 19849 -9841 19875 -9785
rect 19931 -9841 19956 -9785
rect 20012 -9841 20037 -9785
rect 20093 -9841 20118 -9785
rect 20174 -9841 20199 -9785
rect 20255 -9841 20280 -9785
rect 20336 -9841 20361 -9785
rect 20417 -9841 20443 -9785
rect 20499 -9841 20524 -9785
rect 20580 -9841 20605 -9785
rect 20661 -9841 20686 -9785
rect 20742 -9841 20767 -9785
rect 20823 -9841 20848 -9785
rect 20904 -9841 20929 -9785
rect 20985 -9841 21011 -9785
rect 21067 -9841 21092 -9785
rect 21148 -9841 21173 -9785
rect 21229 -9841 21254 -9785
rect 21310 -9841 21335 -9785
rect 21391 -9841 21416 -9785
rect 21472 -9841 21497 -9785
rect 21553 -9841 21579 -9785
rect 21635 -9841 21660 -9785
rect 21716 -9841 21741 -9785
rect 21797 -9841 21822 -9785
rect 21878 -9841 21903 -9785
rect 21959 -9841 21984 -9785
rect 22040 -9841 22065 -9785
rect 22121 -9841 22147 -9785
rect 22203 -9841 22228 -9785
rect 22284 -9841 22309 -9785
rect 22365 -9841 22390 -9785
rect 22446 -9841 22471 -9785
rect 22527 -9841 22552 -9785
rect 22608 -9841 22633 -9785
rect 22689 -9841 22715 -9785
rect 22771 -9841 22796 -9785
rect 22852 -9841 22877 -9785
rect 22933 -9841 22958 -9785
rect 23014 -9841 23039 -9785
rect 23095 -9841 23120 -9785
rect 23176 -9841 23201 -9785
rect 23257 -9841 23283 -9785
rect 23339 -9841 23364 -9785
rect 23420 -9841 23445 -9785
rect 23501 -9841 23526 -9785
rect 23582 -9841 23607 -9785
rect 23663 -9841 23688 -9785
rect 23744 -9841 23769 -9785
rect 23825 -9841 23851 -9785
rect 23907 -9841 23932 -9785
rect 23988 -9841 24013 -9785
rect 24069 -9841 24094 -9785
rect 24150 -9841 24175 -9785
rect 24231 -9841 24256 -9785
rect 24312 -9841 24337 -9785
rect 24393 -9841 24419 -9785
rect 24475 -9841 24500 -9785
rect 24556 -9841 24581 -9785
rect 24637 -9841 24662 -9785
rect 24718 -9841 24743 -9785
rect 24799 -9841 24824 -9785
rect 24880 -9841 24905 -9785
rect 24961 -9841 24987 -9785
rect 25043 -9841 25068 -9785
rect 25124 -9841 25149 -9785
rect 25205 -9841 25230 -9785
rect 25286 -9841 25311 -9785
rect 25367 -9841 25392 -9785
rect 25448 -9841 25473 -9785
rect 25529 -9841 25555 -9785
rect 25611 -9841 25636 -9785
rect 25692 -9841 25717 -9785
rect 25773 -9841 25798 -9785
rect 25854 -9841 25879 -9785
rect 25935 -9841 25960 -9785
rect 26016 -9841 26041 -9785
rect 26097 -9841 26123 -9785
rect 26179 -9841 26204 -9785
rect 26260 -9841 26275 -9785
rect 4044 -9889 26275 -9841
rect 4044 -9945 4053 -9889
rect 4109 -9945 4134 -9889
rect 4190 -9945 4215 -9889
rect 4271 -9945 4296 -9889
rect 4352 -9945 4377 -9889
rect 4433 -9945 4458 -9889
rect 4514 -9945 4539 -9889
rect 4595 -9945 4621 -9889
rect 4677 -9945 4702 -9889
rect 4758 -9945 4783 -9889
rect 4839 -9945 4864 -9889
rect 4920 -9945 4945 -9889
rect 5001 -9945 5026 -9889
rect 5082 -9945 5107 -9889
rect 5163 -9945 5189 -9889
rect 5245 -9945 5270 -9889
rect 5326 -9945 5351 -9889
rect 5407 -9945 5432 -9889
rect 5488 -9945 5513 -9889
rect 5569 -9945 5594 -9889
rect 5650 -9945 5675 -9889
rect 5731 -9945 5757 -9889
rect 5813 -9945 5838 -9889
rect 5894 -9945 5919 -9889
rect 5975 -9945 6000 -9889
rect 6056 -9945 6081 -9889
rect 6137 -9945 6162 -9889
rect 6218 -9945 6243 -9889
rect 6299 -9945 6325 -9889
rect 6381 -9945 6406 -9889
rect 6462 -9945 6487 -9889
rect 6543 -9945 6568 -9889
rect 6624 -9945 6649 -9889
rect 6705 -9945 6730 -9889
rect 6786 -9945 6811 -9889
rect 6867 -9945 6893 -9889
rect 6949 -9945 6974 -9889
rect 7030 -9945 7055 -9889
rect 7111 -9945 7136 -9889
rect 7192 -9945 7217 -9889
rect 7273 -9945 7298 -9889
rect 7354 -9945 7379 -9889
rect 7435 -9945 7461 -9889
rect 7517 -9945 7542 -9889
rect 7598 -9945 7623 -9889
rect 7679 -9945 7704 -9889
rect 7760 -9945 7785 -9889
rect 7841 -9945 7866 -9889
rect 7922 -9945 7947 -9889
rect 8003 -9945 8029 -9889
rect 8085 -9945 8110 -9889
rect 8166 -9945 8191 -9889
rect 8247 -9945 8272 -9889
rect 8328 -9945 8353 -9889
rect 8409 -9945 8434 -9889
rect 8490 -9945 8515 -9889
rect 8571 -9945 8597 -9889
rect 8653 -9945 8678 -9889
rect 8734 -9945 8759 -9889
rect 8815 -9945 8840 -9889
rect 8896 -9945 8921 -9889
rect 8977 -9945 9002 -9889
rect 9058 -9945 9083 -9889
rect 9139 -9945 9165 -9889
rect 9221 -9945 9246 -9889
rect 9302 -9945 9327 -9889
rect 9383 -9945 9408 -9889
rect 9464 -9945 9489 -9889
rect 9545 -9945 9570 -9889
rect 9626 -9945 9651 -9889
rect 9707 -9945 9733 -9889
rect 9789 -9945 9814 -9889
rect 9870 -9945 9895 -9889
rect 9951 -9945 9976 -9889
rect 10032 -9945 10057 -9889
rect 10113 -9945 10138 -9889
rect 10194 -9945 10219 -9889
rect 10275 -9945 10301 -9889
rect 10357 -9945 10382 -9889
rect 10438 -9945 10463 -9889
rect 10519 -9945 10544 -9889
rect 10600 -9945 10625 -9889
rect 10681 -9945 10706 -9889
rect 10762 -9945 10787 -9889
rect 10843 -9945 10869 -9889
rect 10925 -9945 10950 -9889
rect 11006 -9945 11031 -9889
rect 11087 -9945 11112 -9889
rect 11168 -9945 11193 -9889
rect 11249 -9945 11274 -9889
rect 11330 -9945 11355 -9889
rect 11411 -9945 11437 -9889
rect 11493 -9945 11518 -9889
rect 11574 -9945 11599 -9889
rect 11655 -9945 11680 -9889
rect 11736 -9945 11761 -9889
rect 11817 -9945 11842 -9889
rect 11898 -9945 11923 -9889
rect 11979 -9945 12005 -9889
rect 12061 -9945 12086 -9889
rect 12142 -9945 12167 -9889
rect 12223 -9945 12248 -9889
rect 12304 -9945 12329 -9889
rect 12385 -9945 12410 -9889
rect 12466 -9945 12491 -9889
rect 12547 -9945 12573 -9889
rect 12629 -9945 12654 -9889
rect 12710 -9945 12735 -9889
rect 12791 -9945 12816 -9889
rect 12872 -9945 12897 -9889
rect 12953 -9945 12978 -9889
rect 13034 -9945 13059 -9889
rect 13115 -9945 13141 -9889
rect 13197 -9945 13222 -9889
rect 13278 -9945 13303 -9889
rect 13359 -9945 13384 -9889
rect 13440 -9945 13465 -9889
rect 13521 -9945 13546 -9889
rect 13602 -9945 13627 -9889
rect 13683 -9945 13709 -9889
rect 13765 -9945 13790 -9889
rect 13846 -9945 13871 -9889
rect 13927 -9945 13952 -9889
rect 14008 -9945 14033 -9889
rect 14089 -9945 14114 -9889
rect 14170 -9945 14195 -9889
rect 14251 -9945 14277 -9889
rect 14333 -9945 14358 -9889
rect 14414 -9945 14439 -9889
rect 14495 -9945 14520 -9889
rect 14576 -9945 14601 -9889
rect 14657 -9945 14682 -9889
rect 14738 -9945 14763 -9889
rect 14819 -9945 14845 -9889
rect 14901 -9945 14926 -9889
rect 14982 -9945 15007 -9889
rect 15063 -9945 15088 -9889
rect 15144 -9945 15169 -9889
rect 15225 -9945 15250 -9889
rect 15306 -9945 15331 -9889
rect 15387 -9945 15413 -9889
rect 15469 -9945 15494 -9889
rect 15550 -9945 15575 -9889
rect 15631 -9945 15656 -9889
rect 15712 -9945 15737 -9889
rect 15793 -9945 15818 -9889
rect 15874 -9945 15899 -9889
rect 15955 -9945 15981 -9889
rect 16037 -9945 16062 -9889
rect 16118 -9945 16143 -9889
rect 16199 -9945 16224 -9889
rect 16280 -9945 16305 -9889
rect 16361 -9945 16386 -9889
rect 16442 -9945 16467 -9889
rect 16523 -9945 16549 -9889
rect 16605 -9945 16630 -9889
rect 16686 -9945 16711 -9889
rect 16767 -9945 16792 -9889
rect 16848 -9945 16873 -9889
rect 16929 -9945 16954 -9889
rect 17010 -9945 17035 -9889
rect 17091 -9945 17117 -9889
rect 17173 -9945 17198 -9889
rect 17254 -9945 17279 -9889
rect 17335 -9945 17360 -9889
rect 17416 -9945 17441 -9889
rect 17497 -9945 17522 -9889
rect 17578 -9945 17603 -9889
rect 17659 -9945 17684 -9889
rect 17740 -9945 17765 -9889
rect 17821 -9945 17846 -9889
rect 17902 -9945 17927 -9889
rect 17983 -9945 18008 -9889
rect 18064 -9945 18089 -9889
rect 18145 -9945 18171 -9889
rect 18227 -9945 18252 -9889
rect 18308 -9945 18333 -9889
rect 18389 -9945 18414 -9889
rect 18470 -9945 18495 -9889
rect 18551 -9945 18576 -9889
rect 18632 -9945 18657 -9889
rect 18713 -9945 18739 -9889
rect 18795 -9945 18820 -9889
rect 18876 -9945 18901 -9889
rect 18957 -9945 18982 -9889
rect 19038 -9945 19063 -9889
rect 19119 -9945 19144 -9889
rect 19200 -9945 19225 -9889
rect 19281 -9945 19307 -9889
rect 19363 -9945 19388 -9889
rect 19444 -9945 19469 -9889
rect 19525 -9945 19550 -9889
rect 19606 -9945 19631 -9889
rect 19687 -9945 19712 -9889
rect 19768 -9945 19793 -9889
rect 19849 -9945 19875 -9889
rect 19931 -9945 19956 -9889
rect 20012 -9945 20037 -9889
rect 20093 -9945 20118 -9889
rect 20174 -9945 20199 -9889
rect 20255 -9945 20280 -9889
rect 20336 -9945 20361 -9889
rect 20417 -9945 20443 -9889
rect 20499 -9945 20524 -9889
rect 20580 -9945 20605 -9889
rect 20661 -9945 20686 -9889
rect 20742 -9945 20767 -9889
rect 20823 -9945 20848 -9889
rect 20904 -9945 20929 -9889
rect 20985 -9945 21011 -9889
rect 21067 -9945 21092 -9889
rect 21148 -9945 21173 -9889
rect 21229 -9945 21254 -9889
rect 21310 -9945 21335 -9889
rect 21391 -9945 21416 -9889
rect 21472 -9945 21497 -9889
rect 21553 -9945 21579 -9889
rect 21635 -9945 21660 -9889
rect 21716 -9945 21741 -9889
rect 21797 -9945 21822 -9889
rect 21878 -9945 21903 -9889
rect 21959 -9945 21984 -9889
rect 22040 -9945 22065 -9889
rect 22121 -9945 22147 -9889
rect 22203 -9945 22228 -9889
rect 22284 -9945 22309 -9889
rect 22365 -9945 22390 -9889
rect 22446 -9945 22471 -9889
rect 22527 -9945 22552 -9889
rect 22608 -9945 22633 -9889
rect 22689 -9945 22715 -9889
rect 22771 -9945 22796 -9889
rect 22852 -9945 22877 -9889
rect 22933 -9945 22958 -9889
rect 23014 -9945 23039 -9889
rect 23095 -9945 23120 -9889
rect 23176 -9945 23201 -9889
rect 23257 -9945 23283 -9889
rect 23339 -9945 23364 -9889
rect 23420 -9945 23445 -9889
rect 23501 -9945 23526 -9889
rect 23582 -9945 23607 -9889
rect 23663 -9945 23688 -9889
rect 23744 -9945 23769 -9889
rect 23825 -9945 23851 -9889
rect 23907 -9945 23932 -9889
rect 23988 -9945 24013 -9889
rect 24069 -9945 24094 -9889
rect 24150 -9945 24175 -9889
rect 24231 -9945 24256 -9889
rect 24312 -9945 24337 -9889
rect 24393 -9945 24419 -9889
rect 24475 -9945 24500 -9889
rect 24556 -9945 24581 -9889
rect 24637 -9945 24662 -9889
rect 24718 -9945 24743 -9889
rect 24799 -9945 24824 -9889
rect 24880 -9945 24905 -9889
rect 24961 -9945 24987 -9889
rect 25043 -9945 25068 -9889
rect 25124 -9945 25149 -9889
rect 25205 -9945 25230 -9889
rect 25286 -9945 25311 -9889
rect 25367 -9945 25392 -9889
rect 25448 -9945 25473 -9889
rect 25529 -9945 25555 -9889
rect 25611 -9945 25636 -9889
rect 25692 -9945 25717 -9889
rect 25773 -9945 25798 -9889
rect 25854 -9945 25879 -9889
rect 25935 -9945 25960 -9889
rect 26016 -9945 26041 -9889
rect 26097 -9945 26123 -9889
rect 26179 -9945 26204 -9889
rect 26260 -9945 26275 -9889
rect 4044 -9950 26275 -9945
<< via3 >>
rect 12603 2106 12607 2666
rect 12607 2106 12663 2666
rect 12663 2106 12667 2666
rect 12839 2106 12843 2666
rect 12843 2106 12899 2666
rect 12899 2106 12903 2666
rect 13075 2106 13079 2666
rect 13079 2106 13135 2666
rect 13135 2106 13139 2666
rect 13311 2106 13315 2666
rect 13315 2106 13371 2666
rect 13371 2106 13375 2666
rect 13547 2106 13551 2666
rect 13551 2106 13607 2666
rect 13607 2106 13611 2666
rect 13783 2106 13787 2666
rect 13787 2106 13843 2666
rect 13843 2106 13847 2666
rect 14019 2106 14023 2666
rect 14023 2106 14079 2666
rect 14079 2106 14083 2666
rect 14255 2106 14259 2666
rect 14259 2106 14315 2666
rect 14315 2106 14319 2666
rect 14491 2106 14495 2666
rect 14495 2106 14551 2666
rect 14551 2106 14555 2666
rect 14727 2106 14731 2666
rect 14731 2106 14787 2666
rect 14787 2106 14791 2666
rect 14963 2106 14967 2666
rect 14967 2106 15023 2666
rect 15023 2106 15027 2666
rect 15199 2106 15203 2666
rect 15203 2106 15259 2666
rect 15259 2106 15263 2666
rect 15435 2106 15439 2666
rect 15439 2106 15495 2666
rect 15495 2106 15499 2666
rect 16726 2106 16730 2666
rect 16730 2106 16786 2666
rect 16786 2106 16790 2666
rect 16962 2106 16966 2666
rect 16966 2106 17022 2666
rect 17022 2106 17026 2666
rect 17198 2106 17202 2666
rect 17202 2106 17258 2666
rect 17258 2106 17262 2666
rect 17434 2106 17438 2666
rect 17438 2106 17494 2666
rect 17494 2106 17498 2666
rect 17670 2106 17674 2666
rect 17674 2106 17730 2666
rect 17730 2106 17734 2666
rect 17906 2106 17910 2666
rect 17910 2106 17966 2666
rect 17966 2106 17970 2666
rect 18142 2106 18146 2666
rect 18146 2106 18202 2666
rect 18202 2106 18206 2666
rect 18378 2106 18382 2666
rect 18382 2106 18438 2666
rect 18438 2106 18442 2666
rect 18614 2106 18618 2666
rect 18618 2106 18674 2666
rect 18674 2106 18678 2666
rect 18850 2106 18854 2666
rect 18854 2106 18910 2666
rect 18910 2106 18914 2666
rect 19086 2106 19090 2666
rect 19090 2106 19146 2666
rect 19146 2106 19150 2666
rect 19322 2106 19326 2666
rect 19326 2106 19382 2666
rect 19382 2106 19386 2666
rect 19558 2106 19562 2666
rect 19562 2106 19618 2666
rect 19618 2106 19622 2666
rect 20849 2106 20853 2666
rect 20853 2106 20909 2666
rect 20909 2106 20913 2666
rect 21085 2106 21089 2666
rect 21089 2106 21145 2666
rect 21145 2106 21149 2666
rect 21321 2106 21325 2666
rect 21325 2106 21381 2666
rect 21381 2106 21385 2666
rect 21557 2106 21561 2666
rect 21561 2106 21617 2666
rect 21617 2106 21621 2666
rect 21793 2106 21797 2666
rect 21797 2106 21853 2666
rect 21853 2106 21857 2666
rect 22029 2106 22033 2666
rect 22033 2106 22089 2666
rect 22089 2106 22093 2666
rect 22265 2106 22269 2666
rect 22269 2106 22325 2666
rect 22325 2106 22329 2666
rect 22501 2106 22505 2666
rect 22505 2106 22561 2666
rect 22561 2106 22565 2666
rect 22737 2106 22741 2666
rect 22741 2106 22797 2666
rect 22797 2106 22801 2666
rect 22973 2106 22977 2666
rect 22977 2106 23033 2666
rect 23033 2106 23037 2666
rect 23209 2106 23213 2666
rect 23213 2106 23269 2666
rect 23269 2106 23273 2666
rect 23445 2106 23449 2666
rect 23449 2106 23505 2666
rect 23505 2106 23509 2666
rect 23681 2106 23685 2666
rect 23685 2106 23741 2666
rect 23741 2106 23745 2666
rect 12603 1270 12607 1830
rect 12607 1270 12663 1830
rect 12663 1270 12667 1830
rect 12839 1270 12843 1830
rect 12843 1270 12899 1830
rect 12899 1270 12903 1830
rect 13075 1270 13079 1830
rect 13079 1270 13135 1830
rect 13135 1270 13139 1830
rect 13311 1270 13315 1830
rect 13315 1270 13371 1830
rect 13371 1270 13375 1830
rect 13547 1270 13551 1830
rect 13551 1270 13607 1830
rect 13607 1270 13611 1830
rect 13783 1270 13787 1830
rect 13787 1270 13843 1830
rect 13843 1270 13847 1830
rect 14019 1270 14023 1830
rect 14023 1270 14079 1830
rect 14079 1270 14083 1830
rect 14255 1270 14259 1830
rect 14259 1270 14315 1830
rect 14315 1270 14319 1830
rect 14491 1270 14495 1830
rect 14495 1270 14551 1830
rect 14551 1270 14555 1830
rect 14727 1270 14731 1830
rect 14731 1270 14787 1830
rect 14787 1270 14791 1830
rect 14963 1270 14967 1830
rect 14967 1270 15023 1830
rect 15023 1270 15027 1830
rect 15199 1270 15203 1830
rect 15203 1270 15259 1830
rect 15259 1270 15263 1830
rect 15435 1270 15439 1830
rect 15439 1270 15495 1830
rect 15495 1270 15499 1830
rect 16726 1270 16730 1830
rect 16730 1270 16786 1830
rect 16786 1270 16790 1830
rect 16962 1270 16966 1830
rect 16966 1270 17022 1830
rect 17022 1270 17026 1830
rect 17198 1270 17202 1830
rect 17202 1270 17258 1830
rect 17258 1270 17262 1830
rect 17434 1270 17438 1830
rect 17438 1270 17494 1830
rect 17494 1270 17498 1830
rect 17670 1270 17674 1830
rect 17674 1270 17730 1830
rect 17730 1270 17734 1830
rect 17906 1270 17910 1830
rect 17910 1270 17966 1830
rect 17966 1270 17970 1830
rect 18142 1270 18146 1830
rect 18146 1270 18202 1830
rect 18202 1270 18206 1830
rect 18378 1270 18382 1830
rect 18382 1270 18438 1830
rect 18438 1270 18442 1830
rect 18614 1270 18618 1830
rect 18618 1270 18674 1830
rect 18674 1270 18678 1830
rect 18850 1270 18854 1830
rect 18854 1270 18910 1830
rect 18910 1270 18914 1830
rect 19086 1270 19090 1830
rect 19090 1270 19146 1830
rect 19146 1270 19150 1830
rect 19322 1270 19326 1830
rect 19326 1270 19382 1830
rect 19382 1270 19386 1830
rect 19558 1270 19562 1830
rect 19562 1270 19618 1830
rect 19618 1270 19622 1830
rect 20849 1270 20853 1830
rect 20853 1270 20909 1830
rect 20909 1270 20913 1830
rect 21085 1270 21089 1830
rect 21089 1270 21145 1830
rect 21145 1270 21149 1830
rect 21321 1270 21325 1830
rect 21325 1270 21381 1830
rect 21381 1270 21385 1830
rect 21557 1270 21561 1830
rect 21561 1270 21617 1830
rect 21617 1270 21621 1830
rect 21793 1270 21797 1830
rect 21797 1270 21853 1830
rect 21853 1270 21857 1830
rect 22029 1270 22033 1830
rect 22033 1270 22089 1830
rect 22089 1270 22093 1830
rect 22265 1270 22269 1830
rect 22269 1270 22325 1830
rect 22325 1270 22329 1830
rect 22501 1270 22505 1830
rect 22505 1270 22561 1830
rect 22561 1270 22565 1830
rect 22737 1270 22741 1830
rect 22741 1270 22797 1830
rect 22797 1270 22801 1830
rect 22973 1270 22977 1830
rect 22977 1270 23033 1830
rect 23033 1270 23037 1830
rect 23209 1270 23213 1830
rect 23213 1270 23269 1830
rect 23269 1270 23273 1830
rect 23445 1270 23449 1830
rect 23449 1270 23505 1830
rect 23505 1270 23509 1830
rect 23681 1270 23685 1830
rect 23685 1270 23741 1830
rect 23741 1270 23745 1830
rect 4911 610 4915 1170
rect 4915 610 4971 1170
rect 4971 610 4975 1170
rect 5147 610 5151 1170
rect 5151 610 5207 1170
rect 5207 610 5211 1170
rect 5383 610 5387 1170
rect 5387 610 5443 1170
rect 5443 610 5447 1170
rect 5619 610 5623 1170
rect 5623 610 5679 1170
rect 5679 610 5683 1170
rect 5855 610 5859 1170
rect 5859 610 5915 1170
rect 5915 610 5919 1170
rect 6091 610 6095 1170
rect 6095 610 6151 1170
rect 6151 610 6155 1170
rect 6327 610 6331 1170
rect 6331 610 6387 1170
rect 6387 610 6391 1170
rect 6563 610 6567 1170
rect 6567 610 6623 1170
rect 6623 610 6627 1170
rect 6799 610 6803 1170
rect 6803 610 6859 1170
rect 6859 610 6863 1170
rect 7035 610 7039 1170
rect 7039 610 7095 1170
rect 7095 610 7099 1170
rect 7271 610 7275 1170
rect 7275 610 7331 1170
rect 7331 610 7335 1170
rect 7507 610 7511 1170
rect 7511 610 7567 1170
rect 7567 610 7571 1170
rect 4911 -226 4915 334
rect 4915 -226 4971 334
rect 4971 -226 4975 334
rect 5147 -226 5151 334
rect 5151 -226 5207 334
rect 5207 -226 5211 334
rect 5383 -226 5387 334
rect 5387 -226 5443 334
rect 5443 -226 5447 334
rect 5619 -226 5623 334
rect 5623 -226 5679 334
rect 5679 -226 5683 334
rect 5855 -226 5859 334
rect 5859 -226 5915 334
rect 5915 -226 5919 334
rect 6091 -226 6095 334
rect 6095 -226 6151 334
rect 6151 -226 6155 334
rect 6327 -226 6331 334
rect 6331 -226 6387 334
rect 6387 -226 6391 334
rect 6563 -226 6567 334
rect 6567 -226 6623 334
rect 6623 -226 6627 334
rect 6799 -226 6803 334
rect 6803 -226 6859 334
rect 6859 -226 6863 334
rect 7035 -226 7039 334
rect 7039 -226 7095 334
rect 7095 -226 7099 334
rect 7271 -226 7275 334
rect 7275 -226 7331 334
rect 7331 -226 7335 334
rect 7507 -226 7511 334
rect 7511 -226 7567 334
rect 7567 -226 7571 334
rect 4911 -1440 4915 -880
rect 4915 -1440 4971 -880
rect 4971 -1440 4975 -880
rect 5147 -1440 5151 -880
rect 5151 -1440 5207 -880
rect 5207 -1440 5211 -880
rect 5383 -1440 5387 -880
rect 5387 -1440 5443 -880
rect 5443 -1440 5447 -880
rect 5619 -1440 5623 -880
rect 5623 -1440 5679 -880
rect 5679 -1440 5683 -880
rect 5855 -1440 5859 -880
rect 5859 -1440 5915 -880
rect 5915 -1440 5919 -880
rect 6091 -1440 6095 -880
rect 6095 -1440 6151 -880
rect 6151 -1440 6155 -880
rect 6327 -1440 6331 -880
rect 6331 -1440 6387 -880
rect 6387 -1440 6391 -880
rect 6563 -1440 6567 -880
rect 6567 -1440 6623 -880
rect 6623 -1440 6627 -880
rect 6799 -1440 6803 -880
rect 6803 -1440 6859 -880
rect 6859 -1440 6863 -880
rect 7035 -1440 7039 -880
rect 7039 -1440 7095 -880
rect 7095 -1440 7099 -880
rect 7271 -1440 7275 -880
rect 7275 -1440 7331 -880
rect 7331 -1440 7335 -880
rect 7507 -1440 7511 -880
rect 7511 -1440 7567 -880
rect 7567 -1440 7571 -880
rect 4911 -2276 4915 -1716
rect 4915 -2276 4971 -1716
rect 4971 -2276 4975 -1716
rect 5147 -2276 5151 -1716
rect 5151 -2276 5207 -1716
rect 5207 -2276 5211 -1716
rect 5383 -2276 5387 -1716
rect 5387 -2276 5443 -1716
rect 5443 -2276 5447 -1716
rect 5619 -2276 5623 -1716
rect 5623 -2276 5679 -1716
rect 5679 -2276 5683 -1716
rect 5855 -2276 5859 -1716
rect 5859 -2276 5915 -1716
rect 5915 -2276 5919 -1716
rect 6091 -2276 6095 -1716
rect 6095 -2276 6151 -1716
rect 6151 -2276 6155 -1716
rect 6327 -2276 6331 -1716
rect 6331 -2276 6387 -1716
rect 6387 -2276 6391 -1716
rect 6563 -2276 6567 -1716
rect 6567 -2276 6623 -1716
rect 6623 -2276 6627 -1716
rect 6799 -2276 6803 -1716
rect 6803 -2276 6859 -1716
rect 6859 -2276 6863 -1716
rect 7035 -2276 7039 -1716
rect 7039 -2276 7095 -1716
rect 7095 -2276 7099 -1716
rect 7271 -2276 7275 -1716
rect 7275 -2276 7331 -1716
rect 7331 -2276 7335 -1716
rect 7507 -2276 7511 -1716
rect 7511 -2276 7567 -1716
rect 7567 -2276 7571 -1716
rect 7983 -3490 7987 -2930
rect 7987 -3490 8043 -2930
rect 8043 -3490 8047 -2930
rect 8219 -3490 8223 -2930
rect 8223 -3490 8279 -2930
rect 8279 -3490 8283 -2930
rect 8455 -3490 8459 -2930
rect 8459 -3490 8515 -2930
rect 8515 -3490 8519 -2930
rect 8691 -3490 8695 -2930
rect 8695 -3490 8751 -2930
rect 8751 -3490 8755 -2930
rect 8927 -3490 8931 -2930
rect 8931 -3490 8987 -2930
rect 8987 -3490 8991 -2930
rect 9163 -3490 9167 -2930
rect 9167 -3490 9223 -2930
rect 9223 -3490 9227 -2930
rect 9399 -3490 9403 -2930
rect 9403 -3490 9459 -2930
rect 9459 -3490 9463 -2930
rect 9635 -3490 9639 -2930
rect 9639 -3490 9695 -2930
rect 9695 -3490 9699 -2930
rect 9871 -3490 9875 -2930
rect 9875 -3490 9931 -2930
rect 9931 -3490 9935 -2930
rect 10107 -3490 10111 -2930
rect 10111 -3490 10167 -2930
rect 10167 -3490 10171 -2930
rect 10343 -3490 10347 -2930
rect 10347 -3490 10403 -2930
rect 10403 -3490 10407 -2930
rect 10579 -3490 10583 -2930
rect 10583 -3490 10639 -2930
rect 10639 -3490 10643 -2930
rect 7983 -4326 7987 -3766
rect 7987 -4326 8043 -3766
rect 8043 -4326 8047 -3766
rect 8219 -4326 8223 -3766
rect 8223 -4326 8279 -3766
rect 8279 -4326 8283 -3766
rect 8455 -4326 8459 -3766
rect 8459 -4326 8515 -3766
rect 8515 -4326 8519 -3766
rect 8691 -4326 8695 -3766
rect 8695 -4326 8751 -3766
rect 8751 -4326 8755 -3766
rect 8927 -4326 8931 -3766
rect 8931 -4326 8987 -3766
rect 8987 -4326 8991 -3766
rect 9163 -4326 9167 -3766
rect 9167 -4326 9223 -3766
rect 9223 -4326 9227 -3766
rect 9399 -4326 9403 -3766
rect 9403 -4326 9459 -3766
rect 9459 -4326 9463 -3766
rect 9635 -4326 9639 -3766
rect 9639 -4326 9695 -3766
rect 9695 -4326 9699 -3766
rect 9871 -4326 9875 -3766
rect 9875 -4326 9931 -3766
rect 9931 -4326 9935 -3766
rect 10107 -4326 10111 -3766
rect 10111 -4326 10167 -3766
rect 10167 -4326 10171 -3766
rect 10343 -4326 10347 -3766
rect 10347 -4326 10403 -3766
rect 10403 -4326 10407 -3766
rect 10579 -4326 10583 -3766
rect 10583 -4326 10639 -3766
rect 10639 -4326 10643 -3766
rect 7983 -5540 7987 -4980
rect 7987 -5540 8043 -4980
rect 8043 -5540 8047 -4980
rect 8219 -5540 8223 -4980
rect 8223 -5540 8279 -4980
rect 8279 -5540 8283 -4980
rect 8455 -5540 8459 -4980
rect 8459 -5540 8515 -4980
rect 8515 -5540 8519 -4980
rect 8691 -5540 8695 -4980
rect 8695 -5540 8751 -4980
rect 8751 -5540 8755 -4980
rect 8927 -5540 8931 -4980
rect 8931 -5540 8987 -4980
rect 8987 -5540 8991 -4980
rect 9163 -5540 9167 -4980
rect 9167 -5540 9223 -4980
rect 9223 -5540 9227 -4980
rect 9399 -5540 9403 -4980
rect 9403 -5540 9459 -4980
rect 9459 -5540 9463 -4980
rect 9635 -5540 9639 -4980
rect 9639 -5540 9695 -4980
rect 9695 -5540 9699 -4980
rect 9871 -5540 9875 -4980
rect 9875 -5540 9931 -4980
rect 9931 -5540 9935 -4980
rect 10107 -5540 10111 -4980
rect 10111 -5540 10167 -4980
rect 10167 -5540 10171 -4980
rect 10343 -5540 10347 -4980
rect 10347 -5540 10403 -4980
rect 10403 -5540 10407 -4980
rect 10579 -5540 10583 -4980
rect 10583 -5540 10639 -4980
rect 10639 -5540 10643 -4980
rect 7983 -6376 7987 -5816
rect 7987 -6376 8043 -5816
rect 8043 -6376 8047 -5816
rect 8219 -6376 8223 -5816
rect 8223 -6376 8279 -5816
rect 8279 -6376 8283 -5816
rect 8455 -6376 8459 -5816
rect 8459 -6376 8515 -5816
rect 8515 -6376 8519 -5816
rect 8691 -6376 8695 -5816
rect 8695 -6376 8751 -5816
rect 8751 -6376 8755 -5816
rect 8927 -6376 8931 -5816
rect 8931 -6376 8987 -5816
rect 8987 -6376 8991 -5816
rect 9163 -6376 9167 -5816
rect 9167 -6376 9223 -5816
rect 9223 -6376 9227 -5816
rect 9399 -6376 9403 -5816
rect 9403 -6376 9459 -5816
rect 9459 -6376 9463 -5816
rect 9635 -6376 9639 -5816
rect 9639 -6376 9695 -5816
rect 9695 -6376 9699 -5816
rect 9871 -6376 9875 -5816
rect 9875 -6376 9931 -5816
rect 9931 -6376 9935 -5816
rect 10107 -6376 10111 -5816
rect 10111 -6376 10167 -5816
rect 10167 -6376 10171 -5816
rect 10343 -6376 10347 -5816
rect 10347 -6376 10403 -5816
rect 10403 -6376 10407 -5816
rect 10579 -6376 10583 -5816
rect 10583 -6376 10639 -5816
rect 10639 -6376 10643 -5816
rect 5979 -7783 5983 -7223
rect 5983 -7783 6039 -7223
rect 6039 -7783 6043 -7223
rect 6215 -7783 6219 -7223
rect 6219 -7783 6275 -7223
rect 6275 -7783 6279 -7223
rect 6451 -7783 6455 -7223
rect 6455 -7783 6511 -7223
rect 6511 -7783 6515 -7223
rect 6687 -7783 6691 -7223
rect 6691 -7783 6747 -7223
rect 6747 -7783 6751 -7223
rect 6923 -7783 6927 -7223
rect 6927 -7783 6983 -7223
rect 6983 -7783 6987 -7223
rect 7159 -7783 7163 -7223
rect 7163 -7783 7219 -7223
rect 7219 -7783 7223 -7223
rect 7395 -7783 7399 -7223
rect 7399 -7783 7455 -7223
rect 7455 -7783 7459 -7223
rect 7631 -7783 7635 -7223
rect 7635 -7783 7691 -7223
rect 7691 -7783 7695 -7223
rect 7977 -7783 7981 -7223
rect 7981 -7783 8037 -7223
rect 8037 -7783 8041 -7223
rect 8213 -7783 8217 -7223
rect 8217 -7783 8273 -7223
rect 8273 -7783 8277 -7223
rect 8449 -7783 8453 -7223
rect 8453 -7783 8509 -7223
rect 8509 -7783 8513 -7223
rect 8685 -7783 8689 -7223
rect 8689 -7783 8745 -7223
rect 8745 -7783 8749 -7223
rect 8921 -7783 8925 -7223
rect 8925 -7783 8981 -7223
rect 8981 -7783 8985 -7223
rect 9157 -7783 9161 -7223
rect 9161 -7783 9217 -7223
rect 9217 -7783 9221 -7223
rect 9393 -7783 9397 -7223
rect 9397 -7783 9453 -7223
rect 9453 -7783 9457 -7223
rect 9629 -7783 9633 -7223
rect 9633 -7783 9689 -7223
rect 9689 -7783 9693 -7223
rect 5979 -8601 5983 -8041
rect 5983 -8601 6039 -8041
rect 6039 -8601 6043 -8041
rect 6215 -8601 6219 -8041
rect 6219 -8601 6275 -8041
rect 6275 -8601 6279 -8041
rect 6451 -8601 6455 -8041
rect 6455 -8601 6511 -8041
rect 6511 -8601 6515 -8041
rect 6687 -8601 6691 -8041
rect 6691 -8601 6747 -8041
rect 6747 -8601 6751 -8041
rect 6923 -8601 6927 -8041
rect 6927 -8601 6983 -8041
rect 6983 -8601 6987 -8041
rect 7159 -8601 7163 -8041
rect 7163 -8601 7219 -8041
rect 7219 -8601 7223 -8041
rect 7395 -8601 7399 -8041
rect 7399 -8601 7455 -8041
rect 7455 -8601 7459 -8041
rect 7631 -8601 7635 -8041
rect 7635 -8601 7691 -8041
rect 7691 -8601 7695 -8041
rect 7977 -8601 7981 -8041
rect 7981 -8601 8037 -8041
rect 8037 -8601 8041 -8041
rect 8213 -8601 8217 -8041
rect 8217 -8601 8273 -8041
rect 8273 -8601 8277 -8041
rect 8449 -8601 8453 -8041
rect 8453 -8601 8509 -8041
rect 8509 -8601 8513 -8041
rect 8685 -8601 8689 -8041
rect 8689 -8601 8745 -8041
rect 8745 -8601 8749 -8041
rect 8921 -8601 8925 -8041
rect 8925 -8601 8981 -8041
rect 8981 -8601 8985 -8041
rect 9157 -8601 9161 -8041
rect 9161 -8601 9217 -8041
rect 9217 -8601 9221 -8041
rect 9393 -8601 9397 -8041
rect 9397 -8601 9453 -8041
rect 9453 -8601 9457 -8041
rect 9629 -8601 9633 -8041
rect 9633 -8601 9689 -8041
rect 9689 -8601 9693 -8041
rect 12667 -7219 12731 -7214
rect 12667 -8054 12671 -7219
rect 12671 -8054 12727 -7219
rect 12727 -8054 12731 -7219
rect 12667 -9205 12671 -8370
rect 12671 -9205 12727 -8370
rect 12727 -9205 12731 -8370
rect 12667 -9210 12731 -9205
rect 12963 -7219 13027 -7214
rect 12963 -8054 12967 -7219
rect 12967 -8054 13023 -7219
rect 13023 -8054 13027 -7219
rect 12963 -9205 12967 -8370
rect 12967 -9205 13023 -8370
rect 13023 -9205 13027 -8370
rect 12963 -9210 13027 -9205
rect 13259 -7219 13323 -7214
rect 13259 -8054 13263 -7219
rect 13263 -8054 13319 -7219
rect 13319 -8054 13323 -7219
rect 13259 -9205 13263 -8370
rect 13263 -9205 13319 -8370
rect 13319 -9205 13323 -8370
rect 13259 -9210 13323 -9205
rect 13555 -7219 13619 -7214
rect 13555 -8054 13559 -7219
rect 13559 -8054 13615 -7219
rect 13615 -8054 13619 -7219
rect 13555 -9205 13559 -8370
rect 13559 -9205 13615 -8370
rect 13615 -9205 13619 -8370
rect 13555 -9210 13619 -9205
rect 13851 -7219 13915 -7214
rect 13851 -8054 13855 -7219
rect 13855 -8054 13911 -7219
rect 13911 -8054 13915 -7219
rect 13851 -9205 13855 -8370
rect 13855 -9205 13911 -8370
rect 13911 -9205 13915 -8370
rect 13851 -9210 13915 -9205
rect 14147 -7219 14211 -7214
rect 14147 -8054 14151 -7219
rect 14151 -8054 14207 -7219
rect 14207 -8054 14211 -7219
rect 14147 -9205 14151 -8370
rect 14151 -9205 14207 -8370
rect 14207 -9205 14211 -8370
rect 14147 -9210 14211 -9205
rect 14443 -7219 14507 -7214
rect 14443 -8054 14447 -7219
rect 14447 -8054 14503 -7219
rect 14503 -8054 14507 -7219
rect 14443 -9205 14447 -8370
rect 14447 -9205 14503 -8370
rect 14503 -9205 14507 -8370
rect 14443 -9210 14507 -9205
rect 14739 -7219 14803 -7214
rect 14739 -8054 14743 -7219
rect 14743 -8054 14799 -7219
rect 14799 -8054 14803 -7219
rect 14739 -9205 14743 -8370
rect 14743 -9205 14799 -8370
rect 14799 -9205 14803 -8370
rect 14739 -9210 14803 -9205
rect 15035 -7219 15099 -7214
rect 15035 -8054 15039 -7219
rect 15039 -8054 15095 -7219
rect 15095 -8054 15099 -7219
rect 15035 -9205 15039 -8370
rect 15039 -9205 15095 -8370
rect 15095 -9205 15099 -8370
rect 15035 -9210 15099 -9205
rect 15331 -7219 15395 -7214
rect 15331 -8054 15335 -7219
rect 15335 -8054 15391 -7219
rect 15391 -8054 15395 -7219
rect 15331 -9205 15335 -8370
rect 15335 -9205 15391 -8370
rect 15391 -9205 15395 -8370
rect 15331 -9210 15395 -9205
rect 15627 -7219 15691 -7214
rect 15627 -8054 15631 -7219
rect 15631 -8054 15687 -7219
rect 15687 -8054 15691 -7219
rect 15627 -9205 15631 -8370
rect 15631 -9205 15687 -8370
rect 15687 -9205 15691 -8370
rect 15627 -9210 15691 -9205
rect 15923 -7219 15987 -7214
rect 15923 -8054 15927 -7219
rect 15927 -8054 15983 -7219
rect 15983 -8054 15987 -7219
rect 15923 -9205 15927 -8370
rect 15927 -9205 15983 -8370
rect 15983 -9205 15987 -8370
rect 15923 -9210 15987 -9205
rect 16219 -7219 16283 -7214
rect 16219 -8054 16223 -7219
rect 16223 -8054 16279 -7219
rect 16279 -8054 16283 -7219
rect 16219 -9205 16223 -8370
rect 16223 -9205 16279 -8370
rect 16279 -9205 16283 -8370
rect 16219 -9210 16283 -9205
rect 16515 -7219 16579 -7214
rect 16515 -8054 16519 -7219
rect 16519 -8054 16575 -7219
rect 16575 -8054 16579 -7219
rect 16515 -9205 16519 -8370
rect 16519 -9205 16575 -8370
rect 16575 -9205 16579 -8370
rect 16515 -9210 16579 -9205
rect 16811 -7219 16875 -7214
rect 16811 -8054 16815 -7219
rect 16815 -8054 16871 -7219
rect 16871 -8054 16875 -7219
rect 16811 -9205 16815 -8370
rect 16815 -9205 16871 -8370
rect 16871 -9205 16875 -8370
rect 16811 -9210 16875 -9205
rect 17107 -7219 17171 -7214
rect 17107 -8054 17111 -7219
rect 17111 -8054 17167 -7219
rect 17167 -8054 17171 -7219
rect 17107 -9205 17111 -8370
rect 17111 -9205 17167 -8370
rect 17167 -9205 17171 -8370
rect 17107 -9210 17171 -9205
rect 17403 -7219 17467 -7214
rect 17403 -8054 17407 -7219
rect 17407 -8054 17463 -7219
rect 17463 -8054 17467 -7219
rect 17403 -9205 17407 -8370
rect 17407 -9205 17463 -8370
rect 17463 -9205 17467 -8370
rect 17403 -9210 17467 -9205
rect 17699 -7219 17763 -7214
rect 17699 -8054 17703 -7219
rect 17703 -8054 17759 -7219
rect 17759 -8054 17763 -7219
rect 17699 -9205 17703 -8370
rect 17703 -9205 17759 -8370
rect 17759 -9205 17763 -8370
rect 17699 -9210 17763 -9205
rect 17995 -7219 18059 -7214
rect 17995 -8054 17999 -7219
rect 17999 -8054 18055 -7219
rect 18055 -8054 18059 -7219
rect 17995 -9205 17999 -8370
rect 17999 -9205 18055 -8370
rect 18055 -9205 18059 -8370
rect 17995 -9210 18059 -9205
rect 18291 -7219 18355 -7214
rect 18291 -8054 18295 -7219
rect 18295 -8054 18351 -7219
rect 18351 -8054 18355 -7219
rect 18291 -9205 18295 -8370
rect 18295 -9205 18351 -8370
rect 18351 -9205 18355 -8370
rect 18291 -9210 18355 -9205
rect 18587 -7219 18651 -7214
rect 18587 -8054 18591 -7219
rect 18591 -8054 18647 -7219
rect 18647 -8054 18651 -7219
rect 18587 -9205 18591 -8370
rect 18591 -9205 18647 -8370
rect 18647 -9205 18651 -8370
rect 18587 -9210 18651 -9205
rect 18883 -7219 18947 -7214
rect 18883 -8054 18887 -7219
rect 18887 -8054 18943 -7219
rect 18943 -8054 18947 -7219
rect 18883 -9205 18887 -8370
rect 18887 -9205 18943 -8370
rect 18943 -9205 18947 -8370
rect 18883 -9210 18947 -9205
rect 19179 -7219 19243 -7214
rect 19179 -8054 19183 -7219
rect 19183 -8054 19239 -7219
rect 19239 -8054 19243 -7219
rect 19179 -9205 19183 -8370
rect 19183 -9205 19239 -8370
rect 19239 -9205 19243 -8370
rect 19179 -9210 19243 -9205
rect 19475 -7219 19539 -7214
rect 19475 -8054 19479 -7219
rect 19479 -8054 19535 -7219
rect 19535 -8054 19539 -7219
rect 19475 -9205 19479 -8370
rect 19479 -9205 19535 -8370
rect 19535 -9205 19539 -8370
rect 19475 -9210 19539 -9205
rect 19771 -7219 19835 -7214
rect 19771 -8054 19775 -7219
rect 19775 -8054 19831 -7219
rect 19831 -8054 19835 -7219
rect 19771 -9205 19775 -8370
rect 19775 -9205 19831 -8370
rect 19831 -9205 19835 -8370
rect 19771 -9210 19835 -9205
rect 20067 -7219 20131 -7214
rect 20067 -8054 20071 -7219
rect 20071 -8054 20127 -7219
rect 20127 -8054 20131 -7219
rect 20067 -9205 20071 -8370
rect 20071 -9205 20127 -8370
rect 20127 -9205 20131 -8370
rect 20067 -9210 20131 -9205
rect 20363 -7219 20427 -7214
rect 20363 -8054 20367 -7219
rect 20367 -8054 20423 -7219
rect 20423 -8054 20427 -7219
rect 20363 -9205 20367 -8370
rect 20367 -9205 20423 -8370
rect 20423 -9205 20427 -8370
rect 20363 -9210 20427 -9205
rect 20659 -7219 20723 -7214
rect 20659 -8054 20663 -7219
rect 20663 -8054 20719 -7219
rect 20719 -8054 20723 -7219
rect 20659 -9205 20663 -8370
rect 20663 -9205 20719 -8370
rect 20719 -9205 20723 -8370
rect 20659 -9210 20723 -9205
rect 20955 -7219 21019 -7214
rect 20955 -8054 20959 -7219
rect 20959 -8054 21015 -7219
rect 21015 -8054 21019 -7219
rect 20955 -9205 20959 -8370
rect 20959 -9205 21015 -8370
rect 21015 -9205 21019 -8370
rect 20955 -9210 21019 -9205
rect 21251 -7219 21315 -7214
rect 21251 -8054 21255 -7219
rect 21255 -8054 21311 -7219
rect 21311 -8054 21315 -7219
rect 21251 -9205 21255 -8370
rect 21255 -9205 21311 -8370
rect 21311 -9205 21315 -8370
rect 21251 -9210 21315 -9205
rect 21547 -7219 21611 -7214
rect 21547 -8054 21551 -7219
rect 21551 -8054 21607 -7219
rect 21607 -8054 21611 -7219
rect 21547 -9205 21551 -8370
rect 21551 -9205 21607 -8370
rect 21607 -9205 21611 -8370
rect 21547 -9210 21611 -9205
rect 21843 -7219 21907 -7214
rect 21843 -8054 21847 -7219
rect 21847 -8054 21903 -7219
rect 21903 -8054 21907 -7219
rect 21843 -9205 21847 -8370
rect 21847 -9205 21903 -8370
rect 21903 -9205 21907 -8370
rect 21843 -9210 21907 -9205
rect 22139 -7219 22203 -7214
rect 22139 -8054 22143 -7219
rect 22143 -8054 22199 -7219
rect 22199 -8054 22203 -7219
rect 22139 -9205 22143 -8370
rect 22143 -9205 22199 -8370
rect 22199 -9205 22203 -8370
rect 22139 -9210 22203 -9205
rect 22435 -7219 22499 -7214
rect 22435 -8054 22439 -7219
rect 22439 -8054 22495 -7219
rect 22495 -8054 22499 -7219
rect 22435 -9205 22439 -8370
rect 22439 -9205 22495 -8370
rect 22495 -9205 22499 -8370
rect 22435 -9210 22499 -9205
rect 22731 -7219 22795 -7214
rect 22731 -8054 22735 -7219
rect 22735 -8054 22791 -7219
rect 22791 -8054 22795 -7219
rect 22731 -9205 22735 -8370
rect 22735 -9205 22791 -8370
rect 22791 -9205 22795 -8370
rect 22731 -9210 22795 -9205
rect 23027 -7219 23091 -7214
rect 23027 -8054 23031 -7219
rect 23031 -8054 23087 -7219
rect 23087 -8054 23091 -7219
rect 23027 -9205 23031 -8370
rect 23031 -9205 23087 -8370
rect 23087 -9205 23091 -8370
rect 23027 -9210 23091 -9205
rect 23323 -7219 23387 -7214
rect 23323 -8054 23327 -7219
rect 23327 -8054 23383 -7219
rect 23383 -8054 23387 -7219
rect 23323 -9205 23327 -8370
rect 23327 -9205 23383 -8370
rect 23383 -9205 23387 -8370
rect 23323 -9210 23387 -9205
rect 23619 -7219 23683 -7214
rect 23619 -8054 23623 -7219
rect 23623 -8054 23679 -7219
rect 23679 -8054 23683 -7219
rect 23619 -9205 23623 -8370
rect 23623 -9205 23679 -8370
rect 23679 -9205 23683 -8370
rect 23619 -9210 23683 -9205
<< metal4 >>
rect 4910 1170 7743 1171
rect 4910 610 4911 1170
rect 4975 610 5147 1170
rect 5211 610 5383 1170
rect 5447 610 5619 1170
rect 5683 610 5855 1170
rect 5919 610 6091 1170
rect 6155 610 6327 1170
rect 6391 610 6563 1170
rect 6627 610 6799 1170
rect 6863 610 7035 1170
rect 7099 610 7271 1170
rect 7335 610 7507 1170
rect 7571 610 7743 1170
rect 4910 334 7743 610
rect 4910 -226 4911 334
rect 4975 -226 5147 334
rect 5211 -226 5383 334
rect 5447 -226 5619 334
rect 5683 -226 5855 334
rect 5919 -226 6091 334
rect 6155 -226 6327 334
rect 6391 -226 6563 334
rect 6627 -226 6799 334
rect 6863 -226 7035 334
rect 7099 -226 7271 334
rect 7335 -226 7507 334
rect 7571 -226 7743 334
rect 4910 -880 7743 -226
rect 4910 -1440 4911 -880
rect 4975 -1440 5147 -880
rect 5211 -1440 5383 -880
rect 5447 -1440 5619 -880
rect 5683 -1440 5855 -880
rect 5919 -1440 6091 -880
rect 6155 -1440 6327 -880
rect 6391 -1440 6563 -880
rect 6627 -1440 6799 -880
rect 6863 -1440 7035 -880
rect 7099 -1440 7271 -880
rect 7335 -1440 7507 -880
rect 7571 -1440 7743 -880
rect 4910 -1716 7743 -1440
rect 4910 -2276 4911 -1716
rect 4975 -2276 5147 -1716
rect 5211 -2276 5383 -1716
rect 5447 -2276 5619 -1716
rect 5683 -2276 5855 -1716
rect 5919 -2276 6091 -1716
rect 6155 -2276 6327 -1716
rect 6391 -2276 6563 -1716
rect 6627 -2276 6799 -1716
rect 6863 -2276 7035 -1716
rect 7099 -2276 7271 -1716
rect 7335 -2276 7507 -1716
rect 7571 -2276 7743 -1716
rect 4910 -2313 7743 -2276
rect 5925 -2691 7513 -2313
rect 5925 -7222 7507 -2691
rect 7811 -2930 10644 -2929
rect 7811 -3490 7983 -2930
rect 8047 -3490 8219 -2930
rect 8283 -3490 8455 -2930
rect 8519 -3490 8691 -2930
rect 8755 -3490 8927 -2930
rect 8991 -3490 9163 -2930
rect 9227 -3490 9399 -2930
rect 9463 -3490 9635 -2930
rect 9699 -3490 9871 -2930
rect 9935 -3490 10107 -2930
rect 10171 -3490 10343 -2930
rect 10407 -3490 10579 -2930
rect 10643 -3490 10644 -2930
rect 7811 -3766 10644 -3490
rect 7811 -4326 7983 -3766
rect 8047 -4326 8219 -3766
rect 8283 -4326 8455 -3766
rect 8519 -4326 8691 -3766
rect 8755 -4326 8927 -3766
rect 8991 -4326 9163 -3766
rect 9227 -4326 9399 -3766
rect 9463 -4326 9635 -3766
rect 9699 -4326 9871 -3766
rect 9935 -4326 10107 -3766
rect 10171 -4326 10343 -3766
rect 10407 -4326 10579 -3766
rect 10643 -4326 10644 -3766
rect 7811 -4980 10644 -4326
rect 7811 -5540 7983 -4980
rect 8047 -5540 8219 -4980
rect 8283 -5540 8455 -4980
rect 8519 -5540 8691 -4980
rect 8755 -5540 8927 -4980
rect 8991 -5540 9163 -4980
rect 9227 -5540 9399 -4980
rect 9463 -5540 9635 -4980
rect 9699 -5540 9871 -4980
rect 9935 -5540 10107 -4980
rect 10171 -5540 10343 -4980
rect 10407 -5540 10579 -4980
rect 10643 -5540 10644 -4980
rect 7811 -5816 10644 -5540
rect 7811 -6376 7983 -5816
rect 8047 -6376 8219 -5816
rect 8283 -6376 8455 -5816
rect 8519 -6376 8691 -5816
rect 8755 -6376 8927 -5816
rect 8991 -6376 9163 -5816
rect 9227 -6376 9399 -5816
rect 9463 -6376 9635 -5816
rect 9699 -6376 9871 -5816
rect 9935 -6376 10107 -5816
rect 10171 -6376 10343 -5816
rect 10407 -6376 10579 -5816
rect 10643 -6376 10644 -5816
rect 7811 -6413 10644 -6376
rect 8041 -7222 9629 -6413
rect 11185 -6970 11486 3181
rect 12602 2666 12668 2667
rect 12602 2106 12603 2666
rect 12667 2106 12668 2666
rect 12602 1830 12668 2106
rect 12602 1270 12603 1830
rect 12667 1270 12668 1830
rect 12602 771 12668 1270
rect 12838 2666 12904 2667
rect 12838 2106 12839 2666
rect 12903 2106 12904 2666
rect 12838 1830 12904 2106
rect 12838 1270 12839 1830
rect 12903 1270 12904 1830
rect 12838 722 12904 1270
rect 13074 2666 13140 2667
rect 13074 2106 13075 2666
rect 13139 2106 13140 2666
rect 13074 1830 13140 2106
rect 13074 1270 13075 1830
rect 13139 1270 13140 1830
rect 13074 719 13140 1270
rect 13310 2666 13376 2667
rect 13310 2106 13311 2666
rect 13375 2106 13376 2666
rect 13310 1830 13376 2106
rect 13310 1270 13311 1830
rect 13375 1270 13376 1830
rect 13310 707 13376 1270
rect 13546 2666 13612 2667
rect 13546 2106 13547 2666
rect 13611 2106 13612 2666
rect 13546 1830 13612 2106
rect 13546 1270 13547 1830
rect 13611 1270 13612 1830
rect 13546 719 13612 1270
rect 13782 2666 13848 2667
rect 13782 2106 13783 2666
rect 13847 2106 13848 2666
rect 13782 1830 13848 2106
rect 13782 1270 13783 1830
rect 13847 1270 13848 1830
rect 13782 859 13848 1270
rect 14018 2666 14084 2667
rect 14018 2106 14019 2666
rect 14083 2106 14084 2666
rect 14018 1830 14084 2106
rect 14018 1270 14019 1830
rect 14083 1270 14084 1830
rect 14018 859 14084 1270
rect 14254 2666 14320 2667
rect 14254 2106 14255 2666
rect 14319 2106 14320 2666
rect 14254 1830 14320 2106
rect 14254 1270 14255 1830
rect 14319 1270 14320 1830
rect 13782 717 14190 859
rect 14254 729 14320 1270
rect 14490 2666 14556 2667
rect 14490 2106 14491 2666
rect 14555 2106 14556 2666
rect 14490 1830 14556 2106
rect 14490 1270 14491 1830
rect 14555 1270 14556 1830
rect 14490 749 14556 1270
rect 14726 2666 14792 2667
rect 14726 2106 14727 2666
rect 14791 2106 14792 2666
rect 14726 1830 14792 2106
rect 14726 1270 14727 1830
rect 14791 1270 14792 1830
rect 14726 727 14792 1270
rect 14962 2666 15028 2667
rect 14962 2106 14963 2666
rect 15027 2106 15028 2666
rect 14962 1830 15028 2106
rect 14962 1270 14963 1830
rect 15027 1270 15028 1830
rect 14962 734 15028 1270
rect 15198 2666 15264 2667
rect 15198 2106 15199 2666
rect 15263 2106 15264 2666
rect 15198 1830 15264 2106
rect 15198 1270 15199 1830
rect 15263 1270 15264 1830
rect 15198 734 15264 1270
rect 15434 2666 15500 2667
rect 15434 2106 15435 2666
rect 15499 2106 15500 2666
rect 15434 1830 15500 2106
rect 15434 1270 15435 1830
rect 15499 1270 15500 1830
rect 5925 -7223 7696 -7222
rect 5925 -7783 5979 -7223
rect 6043 -7783 6215 -7223
rect 6279 -7783 6451 -7223
rect 6515 -7783 6687 -7223
rect 6751 -7783 6923 -7223
rect 6987 -7783 7159 -7223
rect 7223 -7783 7395 -7223
rect 7459 -7783 7631 -7223
rect 7695 -7783 7696 -7223
rect 5925 -8041 7696 -7783
rect 7976 -7223 9694 -7222
rect 7976 -7783 7977 -7223
rect 8041 -7783 8213 -7223
rect 8277 -7783 8449 -7223
rect 8513 -7783 8685 -7223
rect 8749 -7783 8921 -7223
rect 8985 -7783 9157 -7223
rect 9221 -7783 9393 -7223
rect 9457 -7783 9629 -7223
rect 9693 -7783 9694 -7223
rect 11697 -7412 12081 495
rect 12661 -7214 12737 -6676
rect 11697 -7430 11985 -7412
rect 7976 -7784 9694 -7783
rect 7977 -8040 9694 -7784
rect 5925 -8601 5979 -8041
rect 6043 -8601 6215 -8041
rect 6279 -8601 6451 -8041
rect 6515 -8601 6687 -8041
rect 6751 -8601 6923 -8041
rect 6987 -8601 7159 -8041
rect 7223 -8601 7395 -8041
rect 7459 -8601 7631 -8041
rect 7695 -8601 7696 -8041
rect 5925 -8602 6044 -8601
rect 6214 -8602 6280 -8601
rect 6450 -8602 6516 -8601
rect 6686 -8602 6752 -8601
rect 6922 -8602 6988 -8601
rect 7158 -8602 7224 -8601
rect 7394 -8602 7460 -8601
rect 7630 -8602 7696 -8601
rect 7976 -8041 9694 -8040
rect 7976 -8601 7977 -8041
rect 8041 -8601 8213 -8041
rect 8277 -8601 8449 -8041
rect 8513 -8601 8685 -8041
rect 8749 -8601 8921 -8041
rect 8985 -8601 9157 -8041
rect 9221 -8601 9393 -8041
rect 9457 -8601 9629 -8041
rect 9693 -8601 9694 -8041
rect 7976 -8602 8042 -8601
rect 8212 -8602 8278 -8601
rect 8448 -8602 8514 -8601
rect 8684 -8602 8750 -8601
rect 8920 -8602 8986 -8601
rect 9156 -8602 9222 -8601
rect 9392 -8602 9458 -8601
rect 9628 -8602 9694 -8601
rect 12661 -8054 12667 -7214
rect 12731 -8054 12737 -7214
rect 12661 -8370 12737 -8054
rect 12661 -9210 12667 -8370
rect 12731 -9210 12737 -8370
rect 12661 -9212 12737 -9210
rect 12957 -7214 13033 -6721
rect 12957 -8054 12963 -7214
rect 13027 -8054 13033 -7214
rect 12957 -8370 13033 -8054
rect 12957 -9210 12963 -8370
rect 13027 -9210 13033 -8370
rect 12957 -9212 13033 -9210
rect 13253 -7214 13329 -6712
rect 13253 -8054 13259 -7214
rect 13323 -8054 13329 -7214
rect 13253 -8370 13329 -8054
rect 13253 -9210 13259 -8370
rect 13323 -9210 13329 -8370
rect 13253 -9212 13329 -9210
rect 13549 -7214 13625 -6735
rect 13806 -6744 14190 717
rect 15434 712 15500 1270
rect 16725 2666 16791 2667
rect 16725 2106 16726 2666
rect 16790 2106 16791 2666
rect 16725 1830 16791 2106
rect 16725 1270 16726 1830
rect 16790 1270 16791 1830
rect 16725 749 16791 1270
rect 16961 2666 17027 2667
rect 16961 2106 16962 2666
rect 17026 2106 17027 2666
rect 16961 1830 17027 2106
rect 16961 1270 16962 1830
rect 17026 1270 17027 1830
rect 16961 724 17027 1270
rect 17197 2666 17263 2667
rect 17197 2106 17198 2666
rect 17262 2106 17263 2666
rect 17197 1830 17263 2106
rect 17197 1270 17198 1830
rect 17262 1270 17263 1830
rect 17197 710 17263 1270
rect 17433 2666 17499 2667
rect 17433 2106 17434 2666
rect 17498 2106 17499 2666
rect 17433 1830 17499 2106
rect 17433 1270 17434 1830
rect 17498 1270 17499 1830
rect 17433 729 17499 1270
rect 17669 2666 17735 2667
rect 17669 2106 17670 2666
rect 17734 2106 17735 2666
rect 17669 1830 17735 2106
rect 17669 1270 17670 1830
rect 17734 1270 17735 1830
rect 17669 766 17735 1270
rect 17905 2666 17971 2667
rect 17905 2106 17906 2666
rect 17970 2106 17971 2666
rect 17905 1830 17971 2106
rect 17905 1270 17906 1830
rect 17970 1270 17971 1830
rect 17905 759 17971 1270
rect 18141 2666 18207 2667
rect 18141 2106 18142 2666
rect 18206 2106 18207 2666
rect 18141 1830 18207 2106
rect 18141 1270 18142 1830
rect 18206 1270 18207 1830
rect 18141 862 18207 1270
rect 18377 2666 18443 2667
rect 18377 2106 18378 2666
rect 18442 2106 18443 2666
rect 18377 1830 18443 2106
rect 18377 1270 18378 1830
rect 18442 1270 18443 1830
rect 15863 -6416 16247 494
rect 13806 -6815 14217 -6744
rect 13549 -8054 13555 -7214
rect 13619 -8054 13625 -7214
rect 13549 -8370 13625 -8054
rect 13549 -9210 13555 -8370
rect 13619 -9210 13625 -8370
rect 13549 -9212 13625 -9210
rect 13845 -7214 13921 -6815
rect 13845 -8054 13851 -7214
rect 13915 -8054 13921 -7214
rect 13845 -8370 13921 -8054
rect 13845 -9210 13851 -8370
rect 13915 -9210 13921 -8370
rect 13845 -9212 13921 -9210
rect 14141 -7214 14217 -6815
rect 14141 -8054 14147 -7214
rect 14211 -8054 14217 -7214
rect 14141 -8370 14217 -8054
rect 14141 -9210 14147 -8370
rect 14211 -9210 14217 -8370
rect 14141 -9212 14217 -9210
rect 14437 -7214 14513 -6702
rect 14437 -8054 14443 -7214
rect 14507 -8054 14513 -7214
rect 14437 -8370 14513 -8054
rect 14437 -9210 14443 -8370
rect 14507 -9210 14513 -8370
rect 14437 -9212 14513 -9210
rect 14733 -7214 14809 -6673
rect 14733 -8054 14739 -7214
rect 14803 -8054 14809 -7214
rect 14733 -8370 14809 -8054
rect 14733 -9210 14739 -8370
rect 14803 -9210 14809 -8370
rect 14733 -9212 14809 -9210
rect 15029 -7214 15105 -6699
rect 15029 -8054 15035 -7214
rect 15099 -8054 15105 -7214
rect 15029 -8370 15105 -8054
rect 15029 -9210 15035 -8370
rect 15099 -9210 15105 -8370
rect 15029 -9212 15105 -9210
rect 15325 -6743 15401 -6734
rect 15534 -6743 15697 -6558
rect 16509 -6743 16614 -6558
rect 17972 -6657 18356 862
rect 18377 732 18443 1270
rect 18613 2666 18679 2667
rect 18613 2106 18614 2666
rect 18678 2106 18679 2666
rect 18613 1830 18679 2106
rect 18613 1270 18614 1830
rect 18678 1270 18679 1830
rect 18613 741 18679 1270
rect 18849 2666 18915 2667
rect 18849 2106 18850 2666
rect 18914 2106 18915 2666
rect 18849 1830 18915 2106
rect 18849 1270 18850 1830
rect 18914 1270 18915 1830
rect 18849 727 18915 1270
rect 19085 2666 19151 2667
rect 19085 2106 19086 2666
rect 19150 2106 19151 2666
rect 19085 1830 19151 2106
rect 19085 1270 19086 1830
rect 19150 1270 19151 1830
rect 19085 712 19151 1270
rect 19321 2666 19387 2667
rect 19321 2106 19322 2666
rect 19386 2106 19387 2666
rect 19321 1830 19387 2106
rect 19321 1270 19322 1830
rect 19386 1270 19387 1830
rect 19321 729 19387 1270
rect 19557 2666 19623 2667
rect 19557 2106 19558 2666
rect 19622 2106 19623 2666
rect 19557 1830 19623 2106
rect 19557 1270 19558 1830
rect 19622 1270 19623 1830
rect 19557 736 19623 1270
rect 20848 2666 20914 2667
rect 20848 2106 20849 2666
rect 20913 2106 20914 2666
rect 20848 1830 20914 2106
rect 20848 1270 20849 1830
rect 20913 1270 20914 1830
rect 20848 793 20914 1270
rect 21084 2666 21150 2667
rect 21084 2106 21085 2666
rect 21149 2106 21150 2666
rect 21084 1830 21150 2106
rect 21084 1270 21085 1830
rect 21149 1270 21150 1830
rect 21084 798 21150 1270
rect 21320 2666 21386 2667
rect 21320 2106 21321 2666
rect 21385 2106 21386 2666
rect 21320 1830 21386 2106
rect 21320 1270 21321 1830
rect 21385 1270 21386 1830
rect 21320 812 21386 1270
rect 21556 2666 21622 2667
rect 21556 2106 21557 2666
rect 21621 2106 21622 2666
rect 21556 1830 21622 2106
rect 21556 1270 21557 1830
rect 21621 1270 21622 1830
rect 21556 783 21622 1270
rect 21792 2666 21858 2667
rect 21792 2106 21793 2666
rect 21857 2106 21858 2666
rect 21792 1830 21858 2106
rect 21792 1270 21793 1830
rect 21857 1270 21858 1830
rect 21792 751 21858 1270
rect 22028 2666 22094 2667
rect 22028 2106 22029 2666
rect 22093 2106 22094 2666
rect 22028 1830 22094 2106
rect 22028 1270 22029 1830
rect 22093 1270 22094 1830
rect 22028 756 22094 1270
rect 22264 2666 22330 2667
rect 22264 2106 22265 2666
rect 22329 2106 22330 2666
rect 22264 1830 22330 2106
rect 22264 1270 22265 1830
rect 22329 1270 22330 1830
rect 22264 894 22330 1270
rect 22500 2666 22566 2667
rect 22500 2106 22501 2666
rect 22565 2106 22566 2666
rect 22500 1830 22566 2106
rect 22500 1270 22501 1830
rect 22565 1270 22566 1830
rect 22500 894 22566 1270
rect 22138 741 22566 894
rect 22736 2666 22802 2667
rect 22736 2106 22737 2666
rect 22801 2106 22802 2666
rect 22736 1830 22802 2106
rect 22736 1270 22737 1830
rect 22801 1270 22802 1830
rect 20029 -6416 20413 494
rect 22138 -704 22522 741
rect 22736 722 22802 1270
rect 22972 2666 23038 2667
rect 22972 2106 22973 2666
rect 23037 2106 23038 2666
rect 22972 1830 23038 2106
rect 22972 1270 22973 1830
rect 23037 1270 23038 1830
rect 22972 732 23038 1270
rect 23208 2666 23274 2667
rect 23208 2106 23209 2666
rect 23273 2106 23274 2666
rect 23208 1830 23274 2106
rect 23208 1270 23209 1830
rect 23273 1270 23274 1830
rect 23208 749 23274 1270
rect 23444 2666 23510 2667
rect 23444 2106 23445 2666
rect 23509 2106 23510 2666
rect 23444 1830 23510 2106
rect 23444 1270 23445 1830
rect 23509 1270 23510 1830
rect 23444 697 23510 1270
rect 23680 2666 23746 2667
rect 23680 2106 23681 2666
rect 23745 2106 23746 2666
rect 23680 1830 23746 2106
rect 23680 1270 23681 1830
rect 23745 1270 23746 1830
rect 23680 719 23746 1270
rect 22086 -1104 26971 -704
rect 22138 -4540 22522 -1104
rect 26571 -4540 26971 -1104
rect 22047 -4940 26971 -4540
rect 22138 -6552 22522 -4940
rect 16805 -6743 16881 -6657
rect 15325 -6819 15993 -6743
rect 15325 -7214 15401 -6819
rect 15534 -6870 15697 -6819
rect 15325 -8054 15331 -7214
rect 15395 -8054 15401 -7214
rect 15325 -8370 15401 -8054
rect 15325 -9210 15331 -8370
rect 15395 -9210 15401 -8370
rect 15325 -9212 15401 -9210
rect 15621 -7214 15697 -6870
rect 15621 -8054 15627 -7214
rect 15691 -8054 15697 -7214
rect 15621 -8370 15697 -8054
rect 15621 -9210 15627 -8370
rect 15691 -9210 15697 -8370
rect 15621 -9212 15697 -9210
rect 15917 -7214 15993 -6819
rect 15917 -8054 15923 -7214
rect 15987 -8054 15993 -7214
rect 15917 -8370 15993 -8054
rect 15917 -9210 15923 -8370
rect 15987 -9210 15993 -8370
rect 15917 -9212 15993 -9210
rect 16213 -6819 16881 -6743
rect 16213 -7214 16289 -6819
rect 16213 -8054 16219 -7214
rect 16283 -8054 16289 -7214
rect 16213 -8370 16289 -8054
rect 16213 -9210 16219 -8370
rect 16283 -9210 16289 -8370
rect 16213 -9212 16289 -9210
rect 16509 -6870 16614 -6819
rect 16509 -7214 16585 -6870
rect 16509 -8054 16515 -7214
rect 16579 -8054 16585 -7214
rect 16509 -8370 16585 -8054
rect 16509 -9210 16515 -8370
rect 16579 -9210 16585 -8370
rect 16509 -9212 16585 -9210
rect 16805 -7214 16881 -6819
rect 16805 -8054 16811 -7214
rect 16875 -8054 16881 -7214
rect 16805 -8370 16881 -8054
rect 16805 -9210 16811 -8370
rect 16875 -9210 16881 -8370
rect 16805 -9212 16881 -9210
rect 17101 -7214 17177 -6657
rect 17101 -8054 17107 -7214
rect 17171 -8054 17177 -7214
rect 17101 -8370 17177 -8054
rect 17101 -9210 17107 -8370
rect 17171 -9210 17177 -8370
rect 17101 -9212 17177 -9210
rect 17397 -6743 17433 -6657
rect 17735 -6741 17769 -6657
rect 17397 -7214 17473 -6743
rect 17397 -8054 17403 -7214
rect 17467 -8054 17473 -7214
rect 17397 -8370 17473 -8054
rect 17397 -9210 17403 -8370
rect 17467 -9210 17473 -8370
rect 17397 -9212 17473 -9210
rect 17693 -7214 17769 -6741
rect 17972 -6830 18361 -6657
rect 19701 -6751 19840 -6558
rect 22133 -6661 22522 -6552
rect 20357 -6720 20433 -6719
rect 20949 -6720 21025 -6705
rect 17972 -6870 18065 -6830
rect 17693 -8054 17699 -7214
rect 17763 -8054 17769 -7214
rect 17693 -8370 17769 -8054
rect 17693 -9210 17699 -8370
rect 17763 -9210 17769 -8370
rect 17693 -9212 17769 -9210
rect 17989 -7214 18065 -6870
rect 17989 -8054 17995 -7214
rect 18059 -8054 18065 -7214
rect 17989 -8370 18065 -8054
rect 17989 -9210 17995 -8370
rect 18059 -9210 18065 -8370
rect 17989 -9212 18065 -9210
rect 18285 -7214 18361 -6830
rect 18285 -8054 18291 -7214
rect 18355 -8054 18361 -7214
rect 18285 -8370 18361 -8054
rect 18285 -9210 18291 -8370
rect 18355 -9210 18361 -8370
rect 18285 -9212 18361 -9210
rect 18581 -7214 18657 -6775
rect 18581 -8054 18587 -7214
rect 18651 -8054 18657 -7214
rect 18581 -8370 18657 -8054
rect 18581 -9210 18587 -8370
rect 18651 -9210 18657 -8370
rect 18581 -9212 18657 -9210
rect 18877 -7214 18953 -6775
rect 18877 -8054 18883 -7214
rect 18947 -8054 18953 -7214
rect 18877 -8370 18953 -8054
rect 18877 -9210 18883 -8370
rect 18947 -9210 18953 -8370
rect 18877 -9212 18953 -9210
rect 19173 -7214 19249 -6775
rect 19173 -8054 19179 -7214
rect 19243 -8054 19249 -7214
rect 19173 -8370 19249 -8054
rect 19173 -9210 19179 -8370
rect 19243 -9210 19249 -8370
rect 19173 -9212 19249 -9210
rect 19469 -7214 19545 -6775
rect 19701 -6827 20137 -6751
rect 19701 -6870 19841 -6827
rect 19469 -8054 19475 -7214
rect 19539 -8054 19545 -7214
rect 19469 -8370 19545 -8054
rect 19469 -9210 19475 -8370
rect 19539 -9210 19545 -8370
rect 19469 -9212 19545 -9210
rect 19765 -7214 19841 -6870
rect 19765 -8054 19771 -7214
rect 19835 -8054 19841 -7214
rect 19765 -8370 19841 -8054
rect 19765 -9210 19771 -8370
rect 19835 -9210 19841 -8370
rect 19765 -9212 19841 -9210
rect 20061 -7214 20137 -6827
rect 20061 -8054 20067 -7214
rect 20131 -8054 20137 -7214
rect 20061 -8370 20137 -8054
rect 20061 -9210 20067 -8370
rect 20131 -9210 20137 -8370
rect 20061 -9212 20137 -9210
rect 20357 -6796 21042 -6720
rect 20357 -7214 20433 -6796
rect 20357 -8054 20363 -7214
rect 20427 -8054 20433 -7214
rect 20357 -8370 20433 -8054
rect 20357 -9210 20363 -8370
rect 20427 -9210 20433 -8370
rect 20357 -9212 20433 -9210
rect 20653 -7214 20729 -6796
rect 20653 -8054 20659 -7214
rect 20723 -8054 20729 -7214
rect 20653 -8370 20729 -8054
rect 20653 -9210 20659 -8370
rect 20723 -9210 20729 -8370
rect 20653 -9212 20729 -9210
rect 20949 -7214 21025 -6796
rect 20949 -8054 20955 -7214
rect 21019 -8054 21025 -7214
rect 20949 -8370 21025 -8054
rect 20949 -9210 20955 -8370
rect 21019 -9210 21025 -8370
rect 20949 -9212 21025 -9210
rect 21245 -7214 21321 -6705
rect 21245 -8054 21251 -7214
rect 21315 -8054 21321 -7214
rect 21245 -8370 21321 -8054
rect 21245 -9210 21251 -8370
rect 21315 -9210 21321 -8370
rect 21245 -9212 21321 -9210
rect 21541 -7214 21617 -6705
rect 21541 -8054 21547 -7214
rect 21611 -8054 21617 -7214
rect 21541 -8370 21617 -8054
rect 21541 -9210 21547 -8370
rect 21611 -9210 21617 -8370
rect 21541 -9212 21617 -9210
rect 21837 -7214 21913 -6705
rect 22138 -6771 22522 -6661
rect 21837 -8054 21843 -7214
rect 21907 -8054 21913 -7214
rect 21837 -8370 21913 -8054
rect 21837 -9210 21843 -8370
rect 21907 -9210 21913 -8370
rect 21837 -9212 21913 -9210
rect 22133 -6818 22522 -6771
rect 22133 -7214 22209 -6818
rect 22133 -8054 22139 -7214
rect 22203 -8054 22209 -7214
rect 22133 -8370 22209 -8054
rect 22133 -9210 22139 -8370
rect 22203 -9210 22209 -8370
rect 22133 -9212 22209 -9210
rect 22429 -7214 22505 -6818
rect 22429 -8054 22435 -7214
rect 22499 -8054 22505 -7214
rect 22429 -8370 22505 -8054
rect 22429 -9210 22435 -8370
rect 22499 -9210 22505 -8370
rect 22429 -9212 22505 -9210
rect 22725 -7214 22801 -6619
rect 22725 -8054 22731 -7214
rect 22795 -8054 22801 -7214
rect 22725 -8370 22801 -8054
rect 22725 -9210 22731 -8370
rect 22795 -9210 22801 -8370
rect 22725 -9212 22801 -9210
rect 23021 -7214 23097 -6698
rect 23021 -8054 23027 -7214
rect 23091 -8054 23097 -7214
rect 23021 -8370 23097 -8054
rect 23021 -9210 23027 -8370
rect 23091 -9210 23097 -8370
rect 23021 -9212 23097 -9210
rect 23317 -7214 23393 -6724
rect 23317 -8054 23323 -7214
rect 23387 -8054 23393 -7214
rect 23317 -8370 23393 -8054
rect 23317 -9210 23323 -8370
rect 23387 -9210 23393 -8370
rect 23317 -9212 23393 -9210
rect 23613 -7214 23689 -6724
rect 23613 -8054 23619 -7214
rect 23683 -8054 23689 -7214
rect 23613 -8370 23689 -8054
rect 23613 -9210 23619 -8370
rect 23683 -9210 23689 -8370
rect 23613 -9212 23689 -9210
use sky130_fd_pr__cap_mim_m3_1_BLS9H9  sky130_fd_pr__cap_mim_m3_1_BLS9H9_0
timestamp 1606520558
transform -1 0 13922 0 1 -1094
box -1941 -1600 1941 1600
use sky130_fd_pr__cap_mim_m3_1_BLS9H9  sky130_fd_pr__cap_mim_m3_1_BLS9H9_1
timestamp 1606520558
transform -1 0 18088 0 1 -1094
box -1941 -1600 1941 1600
use sky130_fd_pr__cap_mim_m3_1_BLS9H9  sky130_fd_pr__cap_mim_m3_1_BLS9H9_2
timestamp 1606520558
transform -1 0 18088 0 1 -4838
box -1941 -1600 1941 1600
use sky130_fd_pr__cap_mim_m3_1_BLS9H9  sky130_fd_pr__cap_mim_m3_1_BLS9H9_3
timestamp 1606520558
transform -1 0 13922 0 1 -4838
box -1941 -1600 1941 1600
use sky130_fd_pr__cap_mim_m3_1_BLS9H9  sky130_fd_pr__cap_mim_m3_1_BLS9H9_4
timestamp 1606520558
transform -1 0 22254 0 1 -4838
box -1941 -1600 1941 1600
use sky130_fd_pr__cap_mim_m3_1_BLS9H9  sky130_fd_pr__cap_mim_m3_1_BLS9H9_5
timestamp 1606520558
transform -1 0 22254 0 1 -1094
box -1941 -1600 1941 1600
use sky130_fd_pr__nfet_01v8_8HUREQ  sky130_fd_pr__nfet_01v8_8HUREQ_0
timestamp 1606658823
transform 1 0 6778 0 1 -7912
box -1052 -919 1052 919
use sky130_fd_pr__nfet_01v8_8HUREQ  sky130_fd_pr__nfet_01v8_8HUREQ_1
timestamp 1606658823
transform 1 0 8776 0 1 -7912
box -1052 -919 1052 919
use sky130_fd_pr__nfet_01v8_8JUMX6  sky130_fd_pr__nfet_01v8_8JUMX6_0
timestamp 1606595467
transform 1 0 18101 0 1 -8212
box -5717 -1219 5717 1219
use sky130_fd_pr__nfet_01v8_GQFJAV  sky130_fd_pr__nfet_01v8_GQFJAV_0
timestamp 1606787837
transform 1 0 10596 0 1 -7440
box -211 -285 211 285
use sky130_fd_pr__nfet_01v8_GQFJAV  sky130_fd_pr__nfet_01v8_GQFJAV_1
timestamp 1606787837
transform 1 0 10912 0 1 -7440
box -211 -285 211 285
use sky130_fd_pr__nfet_01v8_GQFJAV  sky130_fd_pr__nfet_01v8_GQFJAV_2
timestamp 1606787837
transform 1 0 11544 0 1 -7440
box -211 -285 211 285
use sky130_fd_pr__nfet_01v8_GQFJAV  sky130_fd_pr__nfet_01v8_GQFJAV_3
timestamp 1606787837
transform 1 0 11228 0 1 -7440
box -211 -285 211 285
use sky130_fd_pr__nfet_01v8_GQFJAV  sky130_fd_pr__nfet_01v8_GQFJAV_4
timestamp 1606787837
transform 1 0 12176 0 1 -7440
box -211 -285 211 285
use sky130_fd_pr__nfet_01v8_GQFJAV  sky130_fd_pr__nfet_01v8_GQFJAV_5
timestamp 1606787837
transform 1 0 11860 0 1 -7440
box -211 -285 211 285
use sky130_fd_pr__pfet_01v8_YC9MKB  sky130_fd_pr__pfet_01v8_YC9MKB_0
timestamp 1606712473
transform 1 0 5712 0 1 2387
box -1052 -519 1052 519
use sky130_fd_pr__pfet_01v8_YC9MKB  sky130_fd_pr__pfet_01v8_YC9MKB_1
timestamp 1606712473
transform 1 0 7710 0 1 2387
box -1052 -519 1052 519
use sky130_fd_pr__pfet_01v8_YC9MKB  sky130_fd_pr__pfet_01v8_YC9MKB_2
timestamp 1606712473
transform 1 0 9708 0 1 2387
box -1052 -519 1052 519
use sky130_fd_pr__pfet_01v8_YCMRKB  sky130_fd_pr__pfet_01v8_YCMRKB_0
timestamp 1606658371
transform 1 0 7777 0 1 -3628
box -3117 -937 3117 937
use sky130_fd_pr__pfet_01v8_YCMRKB  sky130_fd_pr__pfet_01v8_YCMRKB_1
timestamp 1606658371
transform 1 0 7777 0 1 -1578
box -3117 -937 3117 937
use sky130_fd_pr__pfet_01v8_YCMRKB  sky130_fd_pr__pfet_01v8_YCMRKB_2
timestamp 1606658371
transform 1 0 7777 0 1 472
box -3117 -937 3117 937
use sky130_fd_pr__pfet_01v8_YCMRKB  sky130_fd_pr__pfet_01v8_YCMRKB_3
timestamp 1606658371
transform 1 0 7777 0 1 -5678
box -3117 -937 3117 937
use sky130_fd_pr__pfet_01v8_YT7TV5  sky130_fd_pr__pfet_01v8_YT7TV5_0
array 0 2 4123 0 0 1874
timestamp 1606718285
transform 1 0 13992 0 1 1968
box -1642 -937 1642 937
use via_li_m1  via_li_m1_0
array 0 94 72 0 0 74
timestamp 1606675505
transform 1 0 4756 0 1 -6599
box 4 0 76 74
use via_li_m1  via_li_m1_1
array 0 114 -72 0 0 74
timestamp 1606675505
transform 0 1 4675 -1 0 -6434
box 4 0 76 74
use via_li_m1  via_li_m1_2
array 0 83 72 0 0 74
timestamp 1606675505
transform 1 0 4756 0 1 -6775
box 4 0 76 74
use via_li_m1  via_li_m1_3
array 0 83 72 0 0 74
timestamp 1606675505
transform 1 0 4756 0 1 1319
box 4 0 76 74
use via_li_m1  via_li_m1_4
array 0 83 72 0 0 74
timestamp 1606675505
transform 1 0 4756 0 1 1407
box 4 0 76 74
use via_li_m1  via_li_m1_5
array 0 83 72 0 0 74
timestamp 1606675505
transform 1 0 4756 0 1 1495
box 4 0 76 74
use via_li_m1  via_li_m1_6
array 0 83 72 0 0 74
timestamp 1606675505
transform 1 0 4756 0 1 3010
box 4 0 76 74
use via_li_m1  via_li_m1_7
array 0 83 72 0 0 74
timestamp 1606675505
transform 1 0 4756 0 1 2816
box 4 0 76 74
use via_li_m1  via_li_m1_8
array 0 83 72 0 0 74
timestamp 1606675505
transform 1 0 4756 0 1 3098
box 4 0 76 74
use via_li_m1  via_li_m1_9
array 0 83 72 0 0 74
timestamp 1606675505
transform 1 0 12446 0 1 2815
box 4 0 76 74
use via_li_m1  via_li_m1_10
array 0 114 -72 0 0 74
timestamp 1606675505
transform 0 1 4592 -1 0 -6434
box 4 0 76 74
use via_li_m1  via_li_m1_11
array 0 83 72 0 0 74
timestamp 1606675505
transform 1 0 18586 0 1 2815
box 4 0 76 74
use via_li_m1  via_li_m1_12
array 0 83 72 0 0 74
timestamp 1606675505
transform 1 0 12467 0 1 1047
box 4 0 76 74
use via_li_m1  via_li_m1_13
array 0 83 72 0 0 74
timestamp 1606675505
transform 1 0 12446 0 1 3097
box 4 0 76 74
use via_li_m1  via_li_m1_14
array 0 83 72 0 0 74
timestamp 1606675505
transform 1 0 12446 0 1 3009
box 4 0 76 74
use via_li_m1  via_li_m1_15
array 0 83 72 0 0 74
timestamp 1606675505
transform 1 0 18585 0 1 3009
box 4 0 76 74
use via_li_m1  via_li_m1_16
array 0 83 72 0 0 74
timestamp 1606675505
transform 1 0 18585 0 1 3097
box 4 0 76 74
use via_li_m1  via_li_m1_17
array 0 83 72 0 0 74
timestamp 1606675505
transform 1 0 18443 0 1 1047
box 4 0 76 74
use via_li_m1  via_li_m1_18
array 0 299 74 0 3 74
timestamp 1606675505
transform 1 0 4048 0 1 -9954
box 4 0 76 74
use via_li_m1  via_li_m1_19
array 0 66 72 0 2 74
timestamp 1606675505
transform 1 0 5758 0 1 -7082
box 4 0 76 74
use via_li_m1  via_li_m1_20
array 0 114 -72 0 0 74
timestamp 1606675505
transform 0 1 4509 -1 0 -6434
box 4 0 76 74
use via_m3_m4  via_m3_m4_0
array 0 3 104 0 2 104
timestamp 1606691473
transform 1 0 11702 0 1 -7588
box -20 -20 84 84
use via_m3_m4  via_m3_m4_1
array 0 5 104 0 2 104
timestamp 1606691473
transform 1 0 15763 0 1 -3102
box -20 -20 84 84
use via_m3_m4  via_m3_m4_2
array 0 5 104 0 2 104
timestamp 1606691473
transform 1 0 19929 0 1 -3102
box -20 -20 84 84
use via_m3_m4  via_m3_m4_3
array 0 5 104 0 2 104
timestamp 1606691473
transform 1 0 11717 0 1 -3102
box -20 -20 84 84
use via_m3_m4  via_m3_m4_4
array 0 29 -104 0 2 -104
timestamp 1606691473
transform -1 0 12581 0 -1 -6786
box -20 -20 84 84
use via_m3_m4  via_m3_m4_5
array 0 29 104 0 2 104
timestamp 1606691473
transform 1 0 16612 0 1 -6850
box -20 -20 84 84
use via_m3_m4  via_m3_m4_6
array 0 29 104 0 2 104
timestamp 1606691473
transform 1 0 20729 0 1 -6850
box -20 -20 84 84
use via_m3_m4  via_m3_m4_7
array 0 29 -104 0 2 -104
timestamp 1606691473
transform -1 0 12581 0 -1 706
box -20 -20 84 84
use via_m3_m4  via_m3_m4_8
array 0 29 104 0 2 104
timestamp 1606691473
transform 1 0 16612 0 1 642
box -20 -20 84 84
use via_m3_m4  via_m3_m4_9
array 0 29 104 0 2 104
timestamp 1606691473
transform 1 0 20729 0 1 642
box -20 -20 84 84
use via_m3_m4  via_m3_m4_10
array 0 3 104 0 2 104
timestamp 1606691473
transform 1 0 11147 0 1 -6947
box -20 -20 84 84
use via_m3_m4  via_m3_m4_11
array 0 3 104 0 2 104
timestamp 1606691473
transform 1 0 11143 0 1 2907
box -20 -20 84 84
use via_m3_m4  via_m3_m4_12
array 0 7 104 0 2 104
timestamp 1606691473
transform 1 0 11395 0 1 -9977
box -20 -20 84 84
use via_sub_m1  via_sub_m1_0
array 0 51 154 0 0 46
timestamp 1606738885
transform 1 0 4056 0 1 -9577
box 0 0 154 46
use via_sub_m1  via_sub_m1_1
array 0 51 154 0 0 46
timestamp 1606738885
transform 1 0 4056 0 1 -9503
box 0 0 154 46
use via_sub_m1  via_sub_m1_2
array 0 51 154 0 0 46
timestamp 1606738885
transform 1 0 4056 0 1 -9429
box 0 0 154 46
use via_sub_m1  via_sub_m1_3
array 0 51 154 0 0 46
timestamp 1606738885
transform 1 0 4056 0 1 -9355
box 0 0 154 46
use via_sub_m1  via_sub_m1_4
array 0 51 154 0 0 46
timestamp 1606738885
transform 1 0 4056 0 1 -9281
box 0 0 154 46
use via_sub_m1  via_sub_m1_5
array 0 51 154 0 0 46
timestamp 1606738885
transform 1 0 4056 0 1 -9207
box 0 0 154 46
use via_sub_m1  via_sub_m1_6
array 0 51 154 0 0 46
timestamp 1606738885
transform 1 0 4056 0 1 -9133
box 0 0 154 46
use via_sub_m1  via_sub_m1_7
array 0 51 154 0 0 46
timestamp 1606738885
transform 1 0 4056 0 1 -9059
box 0 0 154 46
use via_sub_m1  via_sub_m1_8
array 0 51 154 0 0 46
timestamp 1606738885
transform 1 0 4056 0 1 -8985
box 0 0 154 46
use via_sub_m1  via_sub_m1_9
array 0 10 154 0 0 46
timestamp 1606738885
transform 1 0 4056 0 1 -8911
box 0 0 154 46
use via_sub_m1  via_sub_m1_10
array 0 9 154 0 0 46
timestamp 1606738885
transform 1 0 4056 0 1 -8837
box 0 0 154 46
use via_sub_m1  via_sub_m1_11
array 0 10 154 0 0 46
timestamp 1606738885
transform 1 0 10648 0 1 -7905
box 0 0 154 46
use via_sub_m1  via_sub_m1_12
array 0 10 154 0 0 46
timestamp 1606738885
transform 1 0 10648 0 1 -7817
box 0 0 154 46
<< labels >>
rlabel metal3 11059 2913 11702 3175 1 vdd
port 0 nsew
rlabel metal2 2069 1881 4601 2054 1 iref
port 1 nsew
rlabel metal2 3032 -677 4304 -429 1 vin_n
port 2 nsew
rlabel metal2 3032 -4777 4304 -4529 1 vin_p
port 3 nsew
rlabel metal4 26571 -4940 26971 -704 1 vout
port 4 nsew
rlabel metal3 11535 -9950 11913 -9675 1 vss
port 5 nsew
rlabel metal2 7633 -7999 7921 -7825 1 vbn
rlabel metal2 11970 -8299 12580 -8126 1 voe1
<< end >>

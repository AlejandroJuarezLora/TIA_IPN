* NGSPICE file created from TIA.ext - technology: sky130A

.subckt sky130_fd_pr__res_high_po_2p85_RN83L8 a_n285_n4194# a_n285_3762# a_n415_n4324#
X0 a_n285_3762# a_n285_n4194# a_n415_n4324# sky130_fd_pr__res_high_po w=2.85 l=37.6
.ends

.subckt sky130_fd_pr__nfet_01v8_UPGCN9 G D B S
X0 D G S B sky130_fd_pr__nfet_01v8 ad=3.77 pd=26.6 as=1.88 ps=13.3 w=13 l=0.3
X1 D G S B sky130_fd_pr__nfet_01v8 ad=1.88 pd=13.3 as=1.88 ps=13.3 w=13 l=0.3
X2 S G D B sky130_fd_pr__nfet_01v8 ad=1.88 pd=13.3 as=3.77 ps=26.6 w=13 l=0.3
X3 S G D B sky130_fd_pr__nfet_01v8 ad=1.88 pd=13.3 as=1.88 ps=13.3 w=13 l=0.3
.ends

.subckt sky130_fd_pr__res_high_po_2p85_BNWAAK a_n285_3204# a_n285_n3636# a_n415_n3766#
X0 a_n285_3204# a_n285_n3636# a_n415_n3766# sky130_fd_pr__res_high_po w=2.85 l=32
.ends

.subckt sky130_fd_pr__nfet_01v8_LNQ4EK D S G B
X0 D G S B sky130_fd_pr__nfet_01v8 ad=4.35 pd=30.6 as=2.17 ps=15.3 w=15 l=0.3
X1 S G D B sky130_fd_pr__nfet_01v8 ad=2.17 pd=15.3 as=4.35 ps=30.6 w=15 l=0.3
.ends

.subckt sky130_fd_pr__res_high_po_2p85_ZJW47V a_n285_n1186# a_n285_754# a_n415_n1316#
X0 a_n285_754# a_n285_n1186# a_n415_n1316# sky130_fd_pr__res_high_po w=2.85 l=7.54
.ends

.subckt sky130_fd_pr__res_high_po_2p85_6SZAMJ a_n285_419# a_n285_n851# a_n415_n981#
X0 a_n285_419# a_n285_n851# a_n415_n981# sky130_fd_pr__res_high_po w=2.85 l=4.19
.ends

.subckt sky130_fd_pr__pfet_01v8_YT7TV5 a_n505_21# a_n387_21# a_384_118# w_n1642_n937#
+ a_n623_21# a_620_118# a_n387_n815# a_n1150_118# a_n33_n815# a_n741_21# a_321_n815#
+ a_n560_n718# a_675_n815# a_1092_n718# a_n1331_n815# a_n1449_21# a_n914_n718# a_1446_n718#
+ a_1029_n815# a_n151_21# a_n560_118# a_1092_118# a_n269_n815# a_620_n718# a_1328_118#
+ a_30_118# a_203_n815# a_974_n718# a_n442_n718# a_557_n815# a_n796_n718# a_439_21#
+ a_n1213_n815# a_n1213_21# a_n1095_21# a_557_21# a_1328_n718# a_n1331_21# a_n206_118#
+ a_675_21# a_738_118# a_911_21# a_n1268_118# a_793_21# a_n1504_118# a_502_n718# a_n1095_n815#
+ a_856_n718# a_85_n815# a_n324_n718# a_439_n815# a_203_21# a_n678_n718# a_148_118#
+ a_n1449_n815# a_321_21# a_n678_118# a_n33_21# a_n914_118# a_1446_118# a_384_n718#
+ a_1029_21# a_n741_n815# a_30_n718# a_1147_21# a_738_n718# a_n206_n718# a_n324_118#
+ a_1265_21# a_n1150_n718# a_856_118# a_1383_n815# a_1383_21# a_n1386_118# a_n1504_n718#
+ a_266_n718# a_n88_118# a_266_118# a_n623_n815# a_n977_n815# a_502_118# a_n796_118#
+ a_n88_n718# a_n1032_118# a_911_n815# a_n1032_n718# a_1265_n815# a_n1386_n718# a_n151_n815#
+ a_n859_21# a_148_n718# a_n442_118# a_974_118# a_n505_n815# a_n977_21# a_1210_118#
+ a_793_n815# a_n859_n815# a_85_21# a_1210_n718# a_n269_21# a_1147_n815# a_n1268_n718#
X0 a_1446_118# a_1383_21# a_1328_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X1 a_n1032_n718# a_n1095_n815# a_n1150_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X2 a_n796_118# a_n859_21# a_n914_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X3 a_384_118# a_321_21# a_266_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X4 a_384_n718# a_321_n815# a_266_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X5 a_n88_n718# a_n151_n815# a_n206_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X6 a_1328_118# a_1265_21# a_1210_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X7 a_n1150_n718# a_n1213_n815# a_n1268_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X8 a_n678_118# a_n741_21# a_n796_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X9 a_1210_n718# a_1147_n815# a_1092_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X10 a_266_118# a_203_21# a_148_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X11 a_30_n718# a_n33_n815# a_n88_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X12 a_1210_118# a_1147_21# a_1092_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X13 a_n914_n718# a_n977_n815# a_n1032_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X14 a_n560_n718# a_n623_n815# a_n678_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X15 a_1446_n718# a_1383_n815# a_1328_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X16 a_n560_118# a_n623_21# a_n678_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X17 a_266_n718# a_203_n815# a_148_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X18 a_620_n718# a_557_n815# a_502_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X19 a_n1386_118# a_n1449_21# a_n1504_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X20 a_n324_118# a_n387_21# a_n442_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X21 a_856_118# a_793_21# a_738_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X22 a_1092_118# a_1029_21# a_974_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X23 a_n324_n718# a_n387_n815# a_n442_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X24 a_n442_118# a_n505_21# a_n560_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X25 a_148_118# a_85_21# a_30_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X26 a_n1386_n718# a_n1449_n815# a_n1504_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X27 a_856_n718# a_793_n815# a_738_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X28 a_974_118# a_911_21# a_856_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X29 a_1092_n718# a_1029_n815# a_974_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X30 a_n1268_118# a_n1331_21# a_n1386_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X31 a_n206_118# a_n269_21# a_n324_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X32 a_738_118# a_675_21# a_620_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X33 a_n796_n718# a_n859_n815# a_n914_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X34 a_n1032_118# a_n1095_21# a_n1150_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X35 a_148_n718# a_85_n815# a_30_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X36 a_1328_n718# a_1265_n815# a_1210_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X37 a_n88_118# a_n151_21# a_n206_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X38 a_30_118# a_n33_21# a_n88_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X39 a_620_118# a_557_21# a_502_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X40 a_502_n718# a_439_n815# a_384_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X41 a_n1150_118# a_n1213_21# a_n1268_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X42 a_n206_n718# a_n269_n815# a_n324_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X43 a_738_n718# a_675_n815# a_620_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X44 a_n1268_n718# a_n1331_n815# a_n1386_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X45 a_n914_118# a_n977_21# a_n1032_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X46 a_n442_n718# a_n505_n815# a_n560_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X47 a_502_118# a_439_21# a_384_118# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X48 a_974_n718# a_911_n815# a_856_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X49 a_n678_n718# a_n741_n815# a_n796_n718# w_n1642_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
.ends

.subckt sky130_fd_pr__nfet_01v8_8HUREQ a_384_n709# a_557_n797# a_203_n797# a_n387_21#
+ a_n505_21# a_30_n709# a_n623_21# a_738_n709# a_n206_n709# a_n741_21# a_n324_109#
+ a_856_109# a_85_n797# a_n151_21# a_266_n709# a_439_n797# a_n88_109# a_266_109# a_n88_n709#
+ a_502_109# a_n796_109# a_439_21# a_n741_n797# a_557_21# a_148_n709# a_675_21# a_n442_109#
+ a_793_21# a_203_21# a_n623_n797# a_321_21# a_620_109# a_384_109# a_n33_21# a_n560_n709#
+ a_n151_n797# a_n914_n709# a_n1016_n883# a_793_n797# a_n505_n797# a_n859_n797# a_n560_109#
+ a_620_n709# a_n442_n709# a_30_109# a_n796_n709# a_n387_n797# a_321_n797# a_n33_n797#
+ a_n206_109# a_675_n797# a_738_109# a_502_n709# a_n859_21# a_856_n709# a_n324_n709#
+ a_n678_n709# a_148_109# a_85_21# a_n269_n797# a_n678_109# a_n914_109# a_n269_21#
X0 a_n678_109# a_n741_21# a_n796_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X1 a_266_109# a_203_21# a_148_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X2 a_30_n709# a_n33_n797# a_n88_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X3 a_n560_n709# a_n623_n797# a_n678_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X4 a_n560_109# a_n623_21# a_n678_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X5 a_n324_109# a_n387_21# a_n442_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X6 a_266_n709# a_203_n797# a_148_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X7 a_620_n709# a_557_n797# a_502_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X8 a_856_109# a_793_21# a_738_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X9 a_n324_n709# a_n387_n797# a_n442_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X10 a_n442_109# a_n505_21# a_n560_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X11 a_148_109# a_85_21# a_30_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X12 a_856_n709# a_793_n797# a_738_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X13 a_n206_109# a_n269_21# a_n324_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X14 a_738_109# a_675_21# a_620_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X15 a_n796_n709# a_n859_n797# a_n914_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X16 a_148_n709# a_85_n797# a_30_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X17 a_620_109# a_557_21# a_502_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X18 a_n88_109# a_n151_21# a_n206_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X19 a_30_109# a_n33_21# a_n88_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X20 a_502_n709# a_439_n797# a_384_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X21 a_n206_n709# a_n269_n797# a_n324_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X22 a_738_n709# a_675_n797# a_620_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X23 a_n442_n709# a_n505_n797# a_n560_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X24 a_502_109# a_439_21# a_384_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X25 a_n678_n709# a_n741_n797# a_n796_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X26 a_n796_109# a_n859_21# a_n914_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X27 a_384_109# a_321_21# a_266_109# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X28 a_384_n709# a_321_n797# a_266_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X29 a_n88_n709# a_n151_n797# a_n206_n709# a_n1016_n883# sky130_fd_pr__nfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_BLS9H9 m3_n1941_n1600# c1_n1841_n1500#
X0 c1_n1841_n1500# m3_n1941_n1600# sky130_fd_pr__cap_mim_m3_1 l=15 w=17.5
.ends

.subckt sky130_fd_pr__pfet_01v8_YC9MKB a_856_n300# a_n324_n300# a_n505_n397# a_n678_n300#
+ a_793_n397# a_n859_n397# a_384_n300# a_n387_n397# a_30_n300# a_321_n397# a_n33_n397#
+ a_738_n300# a_n206_n300# a_675_n397# a_266_n300# a_n269_n397# a_n88_n300# a_203_n397#
+ a_557_n397# a_148_n300# a_439_n397# a_85_n397# w_n1052_n519# a_n560_n300# a_n741_n397#
+ a_n914_n300# a_620_n300# a_n442_n300# a_n796_n300# a_n623_n397# a_n151_n397# a_502_n300#
X0 a_n560_n300# a_n623_n397# a_n678_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X1 a_30_n300# a_n33_n397# a_n88_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X2 a_266_n300# a_203_n397# a_148_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X3 a_620_n300# a_557_n397# a_502_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X4 a_n324_n300# a_n387_n397# a_n442_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X5 a_856_n300# a_793_n397# a_738_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X6 a_n796_n300# a_n859_n397# a_n914_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X7 a_148_n300# a_85_n397# a_30_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X8 a_502_n300# a_439_n397# a_384_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X9 a_n206_n300# a_n269_n397# a_n324_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X10 a_738_n300# a_675_n397# a_620_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X11 a_n442_n300# a_n505_n397# a_n560_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X12 a_n678_n300# a_n741_n397# a_n796_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X13 a_384_n300# a_321_n397# a_266_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X14 a_n88_n300# a_n151_n397# a_n206_n300# w_n1052_n519# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
.ends

.subckt sky130_fd_pr__nfet_01v8_GQFJAV a_15_n75# a_n69_97# a_n175_n249# a_n73_n75#
X0 a_15_n75# a_n69_97# a_n73_n75# a_n175_n249# sky130_fd_pr__nfet_01v8 ad=0.218 pd=2.08 as=0.218 ps=2.08 w=0.75 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_YCMRKB a_n1390_n815# a_89_n718# a_1678_21# a_915_118#
+ a_1151_n718# a_1914_21# a_n2216_21# a_734_n815# a_n2153_n718# a_380_21# a_n2098_21#
+ a_2032_n815# a_n973_n718# a_n1445_118# a_1796_21# a_1977_118# a_n92_21# a_2386_n815#
+ a_n1744_n815# a_1088_n815# a_n2334_21# w_n3117_n937# a_2803_n718# a_1206_21# a_1505_n718#
+ a_n2507_n718# a_n1209_n718# a_1088_21# a_1859_n718# a_2213_118# a_n2452_21# a_325_118#
+ a_1324_21# a_262_n815# a_n855_118# a_n2743_118# a_n2570_21# a_n328_n815# a_1387_118#
+ a_1442_21# a_1623_118# a_n2570_n815# a_n1272_n815# a_n501_n718# a_1033_n718# a_2331_n718#
+ a_1560_21# a_616_n815# a_n2035_n718# a_89_118# a_n855_n718# a_2685_n718# a_1387_n718#
+ a_2268_n815# a_n2389_n718# a_n2924_n815# a_n1626_n815# a_2685_118# a_n265_118# a_n2153_118#
+ a_797_118# a_n501_118# a_2921_118# a_1033_118# a_2858_21# a_561_n718# a_144_n815#
+ a_n1563_118# a_n383_n718# a_498_n815# a_n2452_n815# a_n1154_n815# a_915_n718# a_2095_118#
+ a_2213_n718# a_2268_21# a_n918_21# a_2331_118# a_n737_n718# a_2567_n718# a_1269_n718#
+ a_443_118# a_n2806_n815# a_2504_21# a_n1508_n815# a_n1681_n718# a_2386_21# a_26_21#
+ a_1560_n815# a_n973_118# a_n2861_118# a_2622_21# a_1741_118# a_1914_n815# a_443_n718#
+ a_n328_21# a_2740_21# a_797_n718# a_n1209_118# a_n800_n815# a_n265_n718# a_2095_n718#
+ a_n446_21# a_n2334_n815# a_n1036_n815# a_n383_118# a_n2271_118# a_n2688_n815# a_2032_21#
+ a_26_n815# a_1151_118# a_n564_21# a_n619_n718# a_2449_n718# a_2150_21# a_n800_21#
+ a_2740_n815# a_n2861_n718# a_n1563_n718# a_1442_n815# a_n619_118# a_n1681_118# a_n682_21#
+ a_n2507_118# a_1796_n815# a_n1508_21# a_n682_n815# a_n1917_n718# a_325_n718# a_n1626_21#
+ a_679_n718# a_n1917_118# a_n210_21# a_n147_n718# a_561_118# a_n2216_n815# a_970_n815#
+ a_n1744_21# a_n1091_n718# a_n1091_118# a_2449_118# a_n1980_n815# a_n1862_21# a_1741_n718#
+ a_n2979_118# a_n1036_21# a_2622_n815# a_n2743_n718# a_n1445_n718# a_1324_n815# a_1859_118#
+ a_n1327_118# a_n1980_21# a_1678_n815# a_n1799_n718# a_n1154_21# a_n210_n815# a_n564_n815#
+ a_207_n718# a_616_21# a_n2098_n815# a_n1272_21# a_n29_118# a_498_21# a_207_118#
+ a_n2389_118# a_734_21# a_852_n815# a_n2271_n718# a_n1390_21# a_n918_n815# a_2150_n815#
+ a_n737_118# a_n2625_118# a_n29_n718# a_1269_118# a_n1862_n815# a_1505_118# a_852_21#
+ a_2921_n718# a_1623_n718# a_n1799_118# a_2504_n815# a_n2625_n718# a_n1327_n718#
+ a_1206_n815# a_1977_n718# a_970_21# a_n2806_21# a_n2979_n718# a_n2688_21# a_2858_n815#
+ a_144_21# a_n92_n815# a_380_n815# a_n147_118# a_n2035_118# a_n2924_21# a_n446_n815#
+ a_2567_118# a_2803_118# a_679_118# a_262_21#
X0 a_561_n718# a_498_n815# a_443_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X1 a_n383_118# a_n446_21# a_n501_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X2 a_n265_n718# a_n328_n815# a_n383_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X3 a_n1445_118# a_n1508_21# a_n1563_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X4 a_915_118# a_852_21# a_797_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X5 a_n2625_n718# a_n2688_n815# a_n2743_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X6 a_1151_n718# a_1088_n815# a_1033_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X7 a_n2153_118# a_n2216_21# a_n2271_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X8 a_797_n718# a_734_n815# a_679_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X9 a_2803_118# a_2740_21# a_2685_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X10 a_2331_n718# a_2268_n815# a_2213_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X11 a_n29_118# a_n92_21# a_n147_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X12 a_n1681_n718# a_n1744_n815# a_n1799_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X13 a_n1209_118# a_n1272_21# a_n1327_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X14 a_1859_118# a_1796_21# a_1741_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X15 a_n2861_n718# a_n2924_n815# a_n2979_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X16 a_n265_118# a_n328_21# a_n383_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X17 a_n1917_n718# a_n1980_n815# a_n2035_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X18 a_n2035_n718# a_n2098_n815# a_n2153_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X19 a_797_118# a_734_21# a_679_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X20 a_1977_118# a_1914_21# a_1859_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X21 a_1269_n718# a_1206_n815# a_1151_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X22 a_1623_n718# a_1560_n815# a_1505_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X23 a_207_n718# a_144_n815# a_89_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X24 a_89_n718# a_26_n815# a_n29_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X25 a_n1091_118# a_n1154_21# a_n1209_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X26 a_2685_118# a_2622_21# a_2567_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X27 a_1741_118# a_1678_21# a_1623_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X28 a_2803_n718# a_2740_n815# a_2685_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X29 a_n1091_n718# a_n1154_n815# a_n1209_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X30 a_89_118# a_26_21# a_n29_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X31 a_n2271_n718# a_n2334_n815# a_n2389_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X32 a_1859_n718# a_1796_n815# a_1741_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X33 a_2449_118# a_2386_21# a_2331_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X34 a_n1327_n718# a_n1390_n815# a_n1445_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X35 a_n147_118# a_n210_21# a_n265_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X36 a_n147_n718# a_n210_n815# a_n265_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X37 a_n2861_118# a_n2924_21# a_n2979_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.87 ps=6.58 w=3 l=0.3
X38 a_n501_n718# a_n564_n815# a_n619_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X39 a_n2507_n718# a_n2570_n815# a_n2625_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X40 a_679_118# a_616_21# a_561_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X41 a_443_118# a_380_21# a_325_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X42 a_n973_118# a_n1036_21# a_n1091_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X43 a_n1917_118# a_n1980_21# a_n2035_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X44 a_679_n718# a_616_n815# a_561_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X45 a_1623_118# a_1560_21# a_1505_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X46 a_2213_n718# a_2150_n815# a_2095_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X47 a_2567_118# a_2504_21# a_2449_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X48 a_1033_n718# a_970_n815# a_915_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X49 a_n2625_118# a_n2688_21# a_n2743_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X50 a_n1563_n718# a_n1626_n815# a_n1681_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X51 a_n737_n718# a_n800_n815# a_n855_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X52 a_2331_118# a_2268_21# a_2213_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X53 a_n2743_n718# a_n2806_n815# a_n2861_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X54 a_2449_n718# a_2386_n815# a_2331_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X55 a_561_118# a_498_21# a_443_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X56 a_n1799_n718# a_n1862_n815# a_n1917_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X57 a_n2743_118# a_n2806_21# a_n2861_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X58 a_n737_118# a_n800_21# a_n855_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X59 a_1505_n718# a_1442_n815# a_1387_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X60 a_n1799_118# a_n1862_21# a_n1917_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X61 a_325_118# a_262_21# a_207_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X62 a_443_n718# a_380_n815# a_325_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X63 a_1505_118# a_1442_21# a_1387_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X64 a_2685_n718# a_2622_n815# a_2567_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X65 a_n973_n718# a_n1036_n815# a_n1091_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X66 a_n2507_118# a_n2570_21# a_n2625_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X67 a_n2153_n718# a_n2216_n815# a_n2271_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X68 a_2213_118# a_2150_21# a_2095_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X69 a_n855_118# a_n918_21# a_n973_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X70 a_n1209_n718# a_n1272_n815# a_n1327_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X71 a_n383_n718# a_n446_n815# a_n501_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X72 a_n2389_n718# a_n2452_n815# a_n2507_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X73 a_n1681_118# a_n1744_21# a_n1799_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X74 a_n619_118# a_n682_21# a_n737_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X75 a_1977_n718# a_1914_n815# a_1859_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X76 a_207_118# a_144_21# a_89_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X77 a_2095_n718# a_2032_n815# a_1977_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X78 a_1387_118# a_1324_21# a_1269_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X79 a_915_n718# a_852_n815# a_797_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X80 a_n29_n718# a_n92_n815# a_n147_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X81 a_n1445_n718# a_n1508_n815# a_n1563_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X82 a_n619_n718# a_n682_n815# a_n737_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X83 a_n2389_118# a_n2452_21# a_n2507_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X84 a_2095_118# a_2032_21# a_1977_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X85 a_1151_118# a_1088_21# a_1033_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X86 a_n501_118# a_n564_21# a_n619_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X87 a_1033_118# a_970_21# a_915_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X88 a_n1563_118# a_n1626_21# a_n1681_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X89 a_n855_n718# a_n918_n815# a_n973_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X90 a_1387_n718# a_1324_n815# a_1269_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X91 a_n2271_118# a_n2334_21# a_n2389_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X92 a_1741_n718# a_1678_n815# a_1623_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X93 a_325_n718# a_262_n815# a_207_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X94 a_2921_118# a_2858_21# a_2803_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X95 a_1269_118# a_1206_21# a_1151_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X96 a_2567_n718# a_2504_n815# a_2449_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X97 a_2921_n718# a_2858_n815# a_2803_n718# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.435 ps=3.29 w=3 l=0.3
X98 a_n1327_118# a_n1390_21# a_n1445_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
X99 a_n2035_118# a_n2098_21# a_n2153_118# w_n3117_n937# sky130_fd_pr__pfet_01v8 ad=0.435 pd=3.29 as=0.435 ps=3.29 w=3 l=0.3
.ends

.subckt sky130_fd_pr__nfet_01v8_8JUMX6 a_2117_109# a_n399_n1009# a_1879_n1097# a_5225_109#
+ a_3301_109# a_3803_21# a_547_21# a_785_n1009# a_1377_n1009# a_n193_21# a_n2027_109#
+ a_n3301_21# a_n3597_n1097# a_n3211_109# a_n5135_109# a_2767_n1097# a_4189_n1009#
+ a_3893_109# a_4395_21# a_n1673_n1097# a_2265_n1009# a_4691_n1097# a_n103_109# a_637_n1009#
+ a_n4485_n1097# a_4247_21# a_1229_n1009# a_3655_n1097# a_5077_n1009# a_n2561_n1097#
+ a_785_109# a_3655_21# a_399_21# a_n251_n1009# a_1731_n1097# a_n3449_n1097# a_1969_109#
+ a_2619_n1097# a_3153_n1009# a_n1525_n1097# a_n695_109# a_n3153_21# a_2117_n1009#
+ a_n5373_n1097# a_4543_n1097# a_3507_21# a_n2561_21# a_n4929_21# a_n1879_109# a_n4337_n1097#
+ a_5077_109# a_n4987_109# a_2915_21# a_n3005_21# a_3507_n1097# a_4041_n1009# a_3153_109#
+ a_n1583_n1009# a_n103_n1009# a_n2413_n1097# a_4099_21# a_n2413_21# a_3005_n1009#
+ a_n933_n1097# a_5431_n1097# a_n1821_21# a_n5225_n1097# a_n4395_n1009# a_n3063_109#
+ a_1969_n1009# a_399_n1097# a_n3301_n1097# a_n2471_n1009# a_1229_109# a_n3359_n1009#
+ a_n991_n1009# a_4337_109# a_2413_109# a_3359_21# a_3893_n1009# a_5521_109# a_n1435_n1009#
+ a_2767_21# a_n5283_n1009# a_2857_n1009# a_n1139_109# a_n2265_21# a_n4247_n1009#
+ a_n2323_109# a_n4247_109# a_n5431_109# a_2619_21# a_n1673_21# a_n2323_n1009# a_4781_n1009#
+ a_n843_n1009# a_n2117_21# a_3745_n1009# a_n45_n1097# a_n1525_21# a_n5135_n1009#
+ a_1821_n1009# a_251_n1097# a_45_109# a_2709_n1009# a_n193_n1097# a_1081_109# a_n3211_n1009#
+ a_n3507_109# a_n4929_n1097# a_4633_n1009# a_n991_109# a_n5521_21# a_103_n1097# a_4189_109#
+ a_1879_21# a_251_21# a_n4987_n1009# a_2265_109# a_5521_n1009# a_5373_109# a_n1377_21#
+ a_489_n1009# a_103_21# a_n4099_109# a_n2175_109# a_991_n1097# a_n5283_109# a_n45_21#
+ a_n1229_21# a_1583_n1097# a_341_109# a_n3951_n1009# a_n1377_n1097# a_3449_109# a_1525_109#
+ a_n4839_n1009# a_1081_n1009# a_4633_109# a_n933_21# a_n5373_21# a_n251_109# a_4395_n1097#
+ a_n2915_n1009# a_n4781_21# a_n4189_n1097# a_3359_n1097# a_2471_n1097# a_n1435_109#
+ a_n3359_109# a_n5225_21# a_843_n1097# a_n2265_n1097# a_n4543_109# a_1435_n1097#
+ a_n785_n1097# a_3211_21# a_n4633_21# a_5283_n1097# a_n3803_n1009# a_2709_109# a_341_n1009#
+ a_n1229_n1097# a_n5077_n1097# a_4247_n1097# a_n3153_n1097# a_n785_21# a_2323_n1097#
+ a_n2619_109# a_n2117_n1097# a_n1287_n1009# a_n637_n1097# a_n3803_109# a_4987_21#
+ a_n5077_21# a_5135_n1097# a_n637_21# a_n4041_n1097# a_193_109# a_3063_21# a_n4485_21#
+ a_3211_n1097# a_n4099_n1009# a_n3005_n1097# a_1377_109# a_2471_21# a_n3893_21# a_n2175_n1009#
+ a_4485_109# a_2561_109# a_4839_21# a_n695_n1009# a_n1139_n1009# a_45_n1009# a_3597_n1009#
+ a_n4337_21# a_n1969_n1097# a_2323_21# a_1673_n1009# a_n1287_109# a_n3745_21# a_4987_n1097#
+ a_n2471_109# a_n4395_109# a_1731_21# a_n5681_n1183# a_n3063_n1009# a_n3893_n1097#
+ a_n489_21# a_4485_n1009# a_n2027_n1009# a_3745_109# a_n547_n1009# a_2561_n1009#
+ a_n2857_n1097# a_1821_109# a_3449_n1009# a_933_n1009# a_1525_n1009# a_n4781_n1097#
+ a_3951_n1097# a_4839_n1097# a_5373_n1009# a_n3655_109# a_n5579_109# a_n4189_21#
+ a_n3745_n1097# a_637_109# a_n1731_109# a_2175_21# a_2915_n1097# a_n3597_21# a_4337_n1009#
+ a_n1821_n1097# a_4929_109# a_1583_21# a_n1879_n1009# a_n2709_n1097# a_n547_109#
+ a_2413_n1009# a_2027_21# a_n1081_21# a_n3449_21# a_n4633_n1097# a_3803_n1097# a_5225_n1009#
+ a_n4839_109# a_1435_21# a_n2857_21# a_3005_109# a_n2915_109# a_n2767_n1009# a_3301_n1009#
+ a_n4691_n1009# a_n5521_n1097# a_n2709_21# a_n5579_n1009# a_695_n1097# a_1287_n1097#
+ a_3597_109# a_1673_109# a_5431_21# a_n3655_n1009# a_193_n1009# a_4781_109# a_4099_n1097#
+ a_n2619_n1009# a_n1731_n1009# a_1287_21# a_991_21# a_2175_n1097# a_489_109# a_n1583_109#
+ a_n1081_n1097# a_n4691_109# a_n4543_n1009# a_547_n1097# a_1139_n1097# a_n489_n1097#
+ a_2857_109# a_n399_109# a_1139_21# a_843_21# a_n3507_n1009# a_3063_n1097# a_4929_n1009#
+ a_5283_21# a_n1969_21# a_n5431_n1009# a_n2767_109# a_4691_21# a_2027_n1097# a_n341_21#
+ a_4041_109# a_933_109# a_n3951_109# a_5135_21# a_n843_109# a_4543_21# a_695_21#
+ a_3951_21# a_n4041_21# a_n341_n1097#
X0 a_n4099_109# a_n4189_21# a_n4247_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X1 a_489_n1009# a_399_n1097# a_341_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X2 a_n843_n1009# a_n933_n1097# a_n991_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X3 a_n1731_n1009# a_n1821_n1097# a_n1879_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X4 a_3597_109# a_3507_21# a_3449_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X5 a_n1287_109# a_n1377_21# a_n1435_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X6 a_4633_109# a_4543_21# a_4485_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X7 a_4485_n1009# a_4395_n1097# a_4337_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X8 a_489_109# a_399_21# a_341_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X9 a_2709_109# a_2619_21# a_2561_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X10 a_1821_109# a_1731_21# a_1673_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X11 a_n2027_n1009# a_n2117_n1097# a_n2175_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X12 a_n547_n1009# a_n637_n1097# a_n695_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X13 a_n1435_n1009# a_n1525_n1097# a_n1583_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X14 a_3745_109# a_3655_21# a_3597_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X15 a_4781_109# a_4691_21# a_4633_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X16 a_4189_n1009# a_4099_n1097# a_4041_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X17 a_2857_109# a_2767_21# a_2709_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X18 a_n4839_109# a_n4929_21# a_n4987_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X19 a_5077_n1009# a_4987_n1097# a_4929_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X20 a_n1139_n1009# a_n1229_n1097# a_n1287_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X21 a_1969_109# a_1879_21# a_1821_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X22 a_n2619_n1009# a_n2709_n1097# a_n2767_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X23 a_193_n1009# a_103_n1097# a_45_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X24 a_n3951_n1009# a_n4041_n1097# a_n4099_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X25 a_n5431_n1009# a_n5521_n1097# a_n5579_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=1.3 ps=9.58 w=4.5 l=0.45
X26 a_n547_109# a_n637_21# a_n695_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X27 a_45_109# a_n45_21# a_n103_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X28 a_2117_109# a_2027_21# a_1969_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X29 a_3153_109# a_3063_21# a_3005_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X30 a_n3211_109# a_n3301_21# a_n3359_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X31 a_45_n1009# a_n45_n1097# a_n103_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X32 a_n5135_n1009# a_n5225_n1097# a_n5283_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X33 a_n103_n1009# a_n193_n1097# a_n251_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X34 a_n991_n1009# a_n1081_n1097# a_n1139_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X35 a_n3063_n1009# a_n3153_n1097# a_n3211_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X36 a_n5135_109# a_n5225_21# a_n5283_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X37 a_1229_109# a_1139_21# a_1081_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X38 a_n2471_n1009# a_n2561_n1097# a_n2619_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X39 a_n4543_n1009# a_n4633_n1097# a_n4691_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X40 a_n695_109# a_n785_21# a_n843_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X41 a_3301_n1009# a_3211_n1097# a_3153_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X42 a_2265_109# a_2175_21# a_2117_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X43 a_n2323_109# a_n2413_21# a_n2471_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X44 a_4189_109# a_4099_21# a_4041_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X45 a_n4247_109# a_n4337_21# a_n4395_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X46 a_n5283_109# a_n5373_21# a_n5431_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X47 a_1377_109# a_1287_21# a_1229_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X48 a_n4247_n1009# a_n4337_n1097# a_n4395_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X49 a_n1435_109# a_n1525_21# a_n1583_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X50 a_n2175_n1009# a_n2265_n1097# a_n2323_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X51 a_n3359_109# a_n3449_21# a_n3507_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X52 a_n3655_n1009# a_n3745_n1097# a_n3803_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X53 a_n2471_109# a_n2561_21# a_n2619_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X54 a_n695_n1009# a_n785_n1097# a_n843_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X55 a_n1583_n1009# a_n1673_n1097# a_n1731_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X56 a_637_109# a_547_21# a_489_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X57 a_2413_n1009# a_2323_n1097# a_2265_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X58 a_n4395_109# a_n4485_21# a_n4543_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X59 a_3893_n1009# a_3803_n1097# a_3745_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X60 a_1821_n1009# a_1731_n1097# a_1673_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X61 a_3893_109# a_3803_21# a_3745_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X62 a_n1583_109# a_n1673_21# a_n1731_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X63 a_n3507_109# a_n3597_21# a_n3655_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X64 a_785_109# a_695_21# a_637_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X65 a_n3359_n1009# a_n3449_n1097# a_n3507_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X66 a_3005_109# a_2915_21# a_2857_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X67 a_n399_n1009# a_n489_n1097# a_n547_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X68 a_n1287_n1009# a_n1377_n1097# a_n1435_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X69 a_n4839_n1009# a_n4929_n1097# a_n4987_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X70 a_2117_n1009# a_2027_n1097# a_1969_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X71 a_341_n1009# a_251_n1097# a_193_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X72 a_n2767_n1009# a_n2857_n1097# a_n2915_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X73 a_4929_109# a_4839_21# a_4781_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X74 a_4041_109# a_3951_21# a_3893_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X75 a_n103_109# a_n193_21# a_n251_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X76 a_3597_n1009# a_3507_n1097# a_3449_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X77 a_1525_n1009# a_1435_n1097# a_1377_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X78 a_3005_n1009# a_2915_n1097# a_2857_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X79 a_5077_109# a_4987_21# a_4929_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X80 a_1229_n1009# a_1139_n1097# a_1081_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X81 a_n1879_n1009# a_n1969_n1097# a_n2027_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X82 a_2709_n1009# a_2619_n1097# a_2561_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X83 a_n5283_n1009# a_n5373_n1097# a_n5431_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X84 a_933_n1009# a_843_n1097# a_785_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X85 a_n4691_n1009# a_n4781_n1097# a_n4839_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X86 a_5521_n1009# a_5431_n1097# a_5373_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=1.3 pd=9.58 as=0.652 ps=4.79 w=4.5 l=0.45
X87 a_3301_109# a_3211_21# a_3153_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X88 a_5225_109# a_5135_21# a_5077_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X89 a_n991_109# a_n1081_21# a_n1139_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X90 a_n843_109# a_n933_21# a_n991_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X91 a_2413_109# a_2323_21# a_2265_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X92 a_n4987_n1009# a_n5077_n1097# a_n5135_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X93 a_637_n1009# a_547_n1097# a_489_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X94 a_4337_109# a_4247_21# a_4189_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X95 a_n4395_n1009# a_n4485_n1097# a_n4543_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X96 a_5225_n1009# a_5135_n1097# a_5077_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X97 a_3153_n1009# a_3063_n1097# a_3005_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X98 a_n3803_n1009# a_n3893_n1097# a_n3951_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X99 a_5373_109# a_5283_21# a_5225_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X100 a_n5431_109# a_n5521_21# a_n5579_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=1.3 ps=9.58 w=4.5 l=0.45
X101 a_1525_109# a_1435_21# a_1377_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X102 a_4633_n1009# a_4543_n1097# a_4485_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X103 a_2561_n1009# a_2471_n1097# a_2413_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X104 a_4041_n1009# a_3951_n1097# a_3893_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X105 a_3449_109# a_3359_21# a_3301_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X106 a_2561_109# a_2471_21# a_2413_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X107 a_4485_109# a_4395_21# a_4337_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X108 a_n4543_109# a_n4633_21# a_n4691_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X109 a_n4099_n1009# a_n4189_n1097# a_n4247_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X110 a_1673_109# a_1583_21# a_1525_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X111 a_n3507_n1009# a_n3597_n1097# a_n3655_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X112 a_n2619_109# a_n2709_21# a_n2767_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X113 a_n1731_109# a_n1821_21# a_n1879_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X114 a_4337_n1009# a_4247_n1097# a_4189_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X115 a_2265_n1009# a_2175_n1097# a_2117_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X116 a_n3655_109# a_n3745_21# a_n3803_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X117 a_3745_n1009# a_3655_n1097# a_3597_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X118 a_933_109# a_843_21# a_785_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X119 a_1673_n1009# a_1583_n1097# a_1525_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X120 a_n4691_109# a_n4781_21# a_n4839_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X121 a_n251_109# a_n341_21# a_n399_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X122 a_n2767_109# a_n2857_21# a_n2915_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X123 a_n3803_109# a_n3893_21# a_n3951_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X124 a_1081_109# a_991_21# a_933_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X125 a_3449_n1009# a_3359_n1097# a_3301_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X126 a_4929_n1009# a_4839_n1097# a_4781_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X127 a_1377_n1009# a_1287_n1097# a_1229_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X128 a_n1879_109# a_n1969_21# a_n2027_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X129 a_2857_n1009# a_2767_n1097# a_2709_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X130 a_1081_n1009# a_991_n1097# a_933_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X131 a_n2915_109# a_n3005_21# a_n3063_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X132 a_193_109# a_103_21# a_45_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X133 a_n3951_109# a_n4041_21# a_n4099_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X134 a_n399_109# a_n489_21# a_n547_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X135 a_n3211_n1009# a_n3301_n1097# a_n3359_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X136 a_n251_n1009# a_n341_n1097# a_n399_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X137 a_n2027_109# a_n2117_21# a_n2175_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X138 a_785_n1009# a_695_n1097# a_637_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X139 a_1969_n1009# a_1879_n1097# a_1821_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X140 a_n3063_109# a_n3153_21# a_n3211_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X141 a_5373_n1009# a_5283_n1097# a_5225_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X142 a_341_109# a_251_21# a_193_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X143 a_n4987_109# a_n5077_21# a_n5135_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X144 a_4781_n1009# a_4691_n1097# a_4633_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X145 a_n1139_109# a_n1229_21# a_n1287_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X146 a_n2915_n1009# a_n3005_n1097# a_n3063_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X147 a_n2175_109# a_n2265_21# a_n2323_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
X148 a_5521_109# a_5431_21# a_5373_109# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=1.3 pd=9.58 as=0.652 ps=4.79 w=4.5 l=0.45
X149 a_n2323_n1009# a_n2413_n1097# a_n2471_n1009# a_n5681_n1183# sky130_fd_pr__nfet_01v8 ad=0.652 pd=4.79 as=0.652 ps=4.79 w=4.5 l=0.45
.ends

.subckt opamp_v1 vdd iref vin_n vin_p vout vss a_4019_n9933#
Xsky130_fd_pr__pfet_01v8_YT7TV5_0[0] iref iref vdd vdd iref vdd iref vout iref iref
+ iref vdd iref vdd iref iref vout vout iref iref vdd vdd iref vdd vdd vout iref vout
+ vout iref vdd iref iref iref iref iref vdd iref vout iref vout iref vdd iref vdd
+ vout iref vdd iref vdd iref iref vout vdd iref iref vout iref vout vout vdd iref
+ iref vout iref vout vout vdd iref vout vdd iref iref vout vdd vout vdd vout iref
+ iref vout vdd vdd vdd iref vdd iref vout iref iref vdd vout vout iref iref vout
+ iref iref iref vout iref iref vdd sky130_fd_pr__pfet_01v8_YT7TV5
Xsky130_fd_pr__pfet_01v8_YT7TV5_0[1] iref iref vdd vdd iref vdd iref vout iref iref
+ iref vdd iref vdd iref iref vout vout iref iref vdd vdd iref vdd vdd vout iref vout
+ vout iref vdd iref iref iref iref iref vdd iref vout iref vout iref vdd iref vdd
+ vout iref vdd iref vdd iref iref vout vdd iref iref vout iref vout vout vdd iref
+ iref vout iref vout vout vdd iref vout vdd iref iref vout vdd vout vdd vout iref
+ iref vout vdd vdd vdd iref vdd iref vout iref iref vdd vout vout iref iref vout
+ iref iref iref vout iref iref vdd sky130_fd_pr__pfet_01v8_YT7TV5
Xsky130_fd_pr__pfet_01v8_YT7TV5_0[2] iref iref vdd vdd iref vdd iref vout iref iref
+ iref vdd iref vdd iref iref vout vout iref iref vdd vdd iref vdd vdd vout iref vout
+ vout iref vdd iref iref iref iref iref vdd iref vout iref vout iref vdd iref vdd
+ vout iref vdd iref vdd iref iref vout vdd iref iref vout iref vout vout vdd iref
+ iref vout iref vout vout vdd iref vout vdd iref iref vout vdd vout vdd vout iref
+ iref vout vdd vdd vdd iref vdd iref vout iref iref vdd vout vout iref iref vout
+ iref iref iref vout iref iref vdd sky130_fd_pr__pfet_01v8_YT7TV5
Xsky130_fd_pr__nfet_01v8_8HUREQ_0 vbn vbn vbn vbn vbn vss vbn vss vss vbn vbn vbn
+ vbn vbn vss vbn vbn vss vbn vss vbn vbn vbn vbn vbn vbn vss vbn vbn vbn vbn vbn
+ vbn vbn vbn vbn vss vss vbn vbn vbn vbn vbn vss vss vbn vbn vbn vbn vss vbn vss
+ vss vbn vbn vbn vss vbn vbn vbn vss vss vbn sky130_fd_pr__nfet_01v8_8HUREQ
Xsky130_fd_pr__nfet_01v8_8HUREQ_1 voe1 vbn vbn vbn vbn vss vbn vss vss vbn voe1 voe1
+ vbn vbn vss vbn voe1 vss voe1 vss voe1 vbn vbn vbn voe1 vbn vss vbn vbn vbn vbn
+ voe1 voe1 vbn voe1 vbn vss vss vbn vbn vbn voe1 voe1 vss vss voe1 vbn vbn vbn vss
+ vbn vss vss vbn voe1 voe1 vss voe1 vbn vbn vss vss vbn sky130_fd_pr__nfet_01v8_8HUREQ
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_0 a_10927_n7515# vout sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_1 a_10927_n7515# vout sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_2 a_10927_n7515# vout sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__pfet_01v8_YC9MKB_1 w_4660_n6791# w_4660_n6791# iref vdd iref iref w_4660_n6791#
+ iref vdd iref iref vdd vdd iref vdd iref w_4660_n6791# iref iref w_4660_n6791# iref
+ iref vdd w_4660_n6791# iref vdd w_4660_n6791# vdd w_4660_n6791# iref iref vdd sky130_fd_pr__pfet_01v8_YC9MKB
Xsky130_fd_pr__pfet_01v8_YC9MKB_0 iref iref iref vdd iref iref iref iref vdd iref
+ iref vdd vdd iref vdd iref iref iref iref iref iref iref vdd iref iref vdd iref
+ vdd iref iref iref vdd sky130_fd_pr__pfet_01v8_YC9MKB
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_3 a_10927_n7515# vout sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__pfet_01v8_YC9MKB_2 w_4660_n6791# w_4660_n6791# iref vdd iref iref w_4660_n6791#
+ iref vdd iref iref vdd vdd iref vdd iref w_4660_n6791# iref iref w_4660_n6791# iref
+ iref vdd w_4660_n6791# iref vdd w_4660_n6791# vdd w_4660_n6791# iref iref vdd sky130_fd_pr__pfet_01v8_YC9MKB
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_4 a_10927_n7515# vout sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__cap_mim_m3_1_BLS9H9_5 a_10927_n7515# vout sky130_fd_pr__cap_mim_m3_1_BLS9H9
Xsky130_fd_pr__nfet_01v8_GQFJAV_0 a_10927_n7515# vdd vss voe1 sky130_fd_pr__nfet_01v8_GQFJAV
Xsky130_fd_pr__nfet_01v8_GQFJAV_1 a_10927_n7515# vdd vss voe1 sky130_fd_pr__nfet_01v8_GQFJAV
Xsky130_fd_pr__nfet_01v8_GQFJAV_2 a_10927_n7515# vdd vss voe1 sky130_fd_pr__nfet_01v8_GQFJAV
Xsky130_fd_pr__nfet_01v8_GQFJAV_3 a_10927_n7515# vdd vss voe1 sky130_fd_pr__nfet_01v8_GQFJAV
Xsky130_fd_pr__nfet_01v8_GQFJAV_4 a_10927_n7515# vdd vss voe1 sky130_fd_pr__nfet_01v8_GQFJAV
Xsky130_fd_pr__nfet_01v8_GQFJAV_5 a_10927_n7515# vdd vss voe1 sky130_fd_pr__nfet_01v8_GQFJAV
Xsky130_fd_pr__pfet_01v8_YCMRKB_0 vin_p w_4660_n6791# vin_p voe1 voe1 vin_p vin_p
+ vin_p voe1 vin_p vin_p vin_p voe1 voe1 vin_p w_4660_n6791# vin_p vin_p vin_p vin_p
+ vin_p w_4660_n6791# voe1 vin_p w_4660_n6791# w_4660_n6791# voe1 vin_p voe1 w_4660_n6791#
+ vin_p w_4660_n6791# vin_p vin_p w_4660_n6791# w_4660_n6791# vin_p vin_p voe1 vin_p
+ voe1 vin_p vin_p voe1 w_4660_n6791# voe1 vin_p vin_p w_4660_n6791# w_4660_n6791#
+ w_4660_n6791# w_4660_n6791# voe1 vin_p voe1 vin_p vin_p w_4660_n6791# voe1 voe1
+ w_4660_n6791# voe1 w_4660_n6791# w_4660_n6791# vin_p w_4660_n6791# vin_p w_4660_n6791#
+ w_4660_n6791# vin_p vin_p vin_p voe1 voe1 w_4660_n6791# vin_p vin_p voe1 voe1 voe1
+ w_4660_n6791# voe1 vin_p vin_p vin_p voe1 vin_p vin_p vin_p voe1 voe1 vin_p w_4660_n6791#
+ vin_p voe1 vin_p vin_p w_4660_n6791# voe1 vin_p voe1 voe1 vin_p vin_p vin_p w_4660_n6791#
+ w_4660_n6791# vin_p vin_p vin_p voe1 vin_p w_4660_n6791# w_4660_n6791# vin_p vin_p
+ vin_p voe1 w_4660_n6791# vin_p w_4660_n6791# voe1 vin_p w_4660_n6791# vin_p vin_p
+ vin_p voe1 w_4660_n6791# vin_p voe1 voe1 vin_p w_4660_n6791# w_4660_n6791# vin_p
+ vin_p vin_p w_4660_n6791# w_4660_n6791# w_4660_n6791# vin_p vin_p w_4660_n6791#
+ w_4660_n6791# vin_p vin_p w_4660_n6791# voe1 vin_p voe1 w_4660_n6791# vin_p vin_p
+ w_4660_n6791# vin_p vin_p vin_p voe1 vin_p vin_p vin_p voe1 vin_p voe1 voe1 vin_p
+ vin_p w_4660_n6791# vin_p vin_p vin_p voe1 voe1 voe1 w_4660_n6791# vin_p w_4660_n6791#
+ vin_p w_4660_n6791# voe1 w_4660_n6791# vin_p voe1 w_4660_n6791# vin_p w_4660_n6791#
+ vin_p vin_p w_4660_n6791# vin_p vin_p vin_p vin_p vin_p w_4660_n6791# w_4660_n6791#
+ vin_p vin_p voe1 voe1 voe1 vin_p sky130_fd_pr__pfet_01v8_YCMRKB
Xsky130_fd_pr__pfet_01v8_YCMRKB_1 vin_n w_4660_n6791# vin_n vbn vbn vin_n vin_n vin_n
+ vbn vin_n vin_n vin_n vbn vbn vin_n w_4660_n6791# vin_n vin_n vin_n vin_n vin_n
+ w_4660_n6791# vbn vin_n w_4660_n6791# w_4660_n6791# vbn vin_n vbn w_4660_n6791#
+ vin_n w_4660_n6791# vin_n vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vbn vin_n
+ vbn vin_n vin_n vbn w_4660_n6791# vbn vin_n vin_n w_4660_n6791# w_4660_n6791# w_4660_n6791#
+ w_4660_n6791# vbn vin_n vbn vin_n vin_n w_4660_n6791# vbn vbn w_4660_n6791# vbn
+ w_4660_n6791# w_4660_n6791# vin_n w_4660_n6791# vin_n w_4660_n6791# w_4660_n6791#
+ vin_n vin_n vin_n vbn vbn w_4660_n6791# vin_n vin_n vbn vbn vbn w_4660_n6791# vbn
+ vin_n vin_n vin_n vbn vin_n vin_n vin_n vbn vbn vin_n w_4660_n6791# vin_n vbn vin_n
+ vin_n w_4660_n6791# vbn vin_n vbn vbn vin_n vin_n vin_n w_4660_n6791# w_4660_n6791#
+ vin_n vin_n vin_n vbn vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vin_n vbn w_4660_n6791#
+ vin_n w_4660_n6791# vbn vin_n w_4660_n6791# vin_n vin_n vin_n vbn w_4660_n6791#
+ vin_n vbn vbn vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vin_n w_4660_n6791#
+ w_4660_n6791# w_4660_n6791# vin_n vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n
+ w_4660_n6791# vbn vin_n vbn w_4660_n6791# vin_n vin_n w_4660_n6791# vin_n vin_n
+ vin_n vbn vin_n vin_n vin_n vbn vin_n vbn vbn vin_n vin_n w_4660_n6791# vin_n vin_n
+ vin_n vbn vbn vbn w_4660_n6791# vin_n w_4660_n6791# vin_n w_4660_n6791# vbn w_4660_n6791#
+ vin_n vbn w_4660_n6791# vin_n w_4660_n6791# vin_n vin_n w_4660_n6791# vin_n vin_n
+ vin_n vin_n vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vbn vbn vbn vin_n sky130_fd_pr__pfet_01v8_YCMRKB
Xsky130_fd_pr__pfet_01v8_YCMRKB_2 vin_n w_4660_n6791# vin_n vbn vbn vin_n vin_n vin_n
+ vbn vin_n vin_n vin_n vbn vbn vin_n w_4660_n6791# vin_n vin_n vin_n vin_n vin_n
+ w_4660_n6791# vbn vin_n w_4660_n6791# w_4660_n6791# vbn vin_n vbn w_4660_n6791#
+ vin_n w_4660_n6791# vin_n vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vbn vin_n
+ vbn vin_n vin_n vbn w_4660_n6791# vbn vin_n vin_n w_4660_n6791# w_4660_n6791# w_4660_n6791#
+ w_4660_n6791# vbn vin_n vbn vin_n vin_n w_4660_n6791# vbn vbn w_4660_n6791# vbn
+ w_4660_n6791# w_4660_n6791# vin_n w_4660_n6791# vin_n w_4660_n6791# w_4660_n6791#
+ vin_n vin_n vin_n vbn vbn w_4660_n6791# vin_n vin_n vbn vbn vbn w_4660_n6791# vbn
+ vin_n vin_n vin_n vbn vin_n vin_n vin_n vbn vbn vin_n w_4660_n6791# vin_n vbn vin_n
+ vin_n w_4660_n6791# vbn vin_n vbn vbn vin_n vin_n vin_n w_4660_n6791# w_4660_n6791#
+ vin_n vin_n vin_n vbn vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vin_n vbn w_4660_n6791#
+ vin_n w_4660_n6791# vbn vin_n w_4660_n6791# vin_n vin_n vin_n vbn w_4660_n6791#
+ vin_n vbn vbn vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vin_n w_4660_n6791#
+ w_4660_n6791# w_4660_n6791# vin_n vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n
+ w_4660_n6791# vbn vin_n vbn w_4660_n6791# vin_n vin_n w_4660_n6791# vin_n vin_n
+ vin_n vbn vin_n vin_n vin_n vbn vin_n vbn vbn vin_n vin_n w_4660_n6791# vin_n vin_n
+ vin_n vbn vbn vbn w_4660_n6791# vin_n w_4660_n6791# vin_n w_4660_n6791# vbn w_4660_n6791#
+ vin_n vbn w_4660_n6791# vin_n w_4660_n6791# vin_n vin_n w_4660_n6791# vin_n vin_n
+ vin_n vin_n vin_n w_4660_n6791# w_4660_n6791# vin_n vin_n vbn vbn vbn vin_n sky130_fd_pr__pfet_01v8_YCMRKB
Xsky130_fd_pr__nfet_01v8_8JUMX6_0 vss vout voe1 vout vss voe1 voe1 vout vout voe1
+ vss voe1 voe1 vss vout voe1 vss vss voe1 voe1 vout voe1 vout vss voe1 voe1 vss voe1
+ vss voe1 vout voe1 voe1 vss voe1 voe1 vout voe1 vout voe1 vout voe1 vss voe1 voe1
+ voe1 voe1 voe1 vout voe1 vss vss voe1 voe1 voe1 vout vout vout vout voe1 voe1 voe1
+ vss voe1 voe1 voe1 voe1 vss vout vout voe1 voe1 vout vss vout vout vout vss voe1
+ vss vout vss voe1 vss vout vss voe1 vout vss vout vout voe1 voe1 vss vss vss voe1
+ vout voe1 voe1 vout vss voe1 vss vss voe1 vout vss vss voe1 vout vout voe1 voe1
+ vss voe1 voe1 vss vout vout vss voe1 vout voe1 vss vout voe1 vss voe1 voe1 voe1
+ vss vout voe1 vout vss vout vout vout voe1 voe1 vss voe1 vss voe1 voe1 voe1 voe1
+ vss vout voe1 voe1 voe1 vout voe1 voe1 voe1 voe1 voe1 vss vss vss voe1 voe1 voe1
+ voe1 voe1 voe1 vss voe1 vout voe1 vss voe1 voe1 voe1 voe1 voe1 vout voe1 voe1 voe1
+ vss voe1 vout voe1 voe1 vout vss vout voe1 vout vss vss vss voe1 voe1 voe1 vout
+ vout voe1 voe1 vout vss voe1 vss vout voe1 voe1 vss vss vout vss vout voe1 vss vout
+ vss vss voe1 voe1 voe1 vss vout vss voe1 voe1 vss vss voe1 voe1 voe1 vout voe1 vout
+ voe1 vout voe1 vss vss voe1 voe1 voe1 voe1 voe1 vout vout voe1 voe1 vss vss vout
+ vss vss voe1 voe1 vss voe1 voe1 vss vout voe1 vout vout vss voe1 vss vss voe1 voe1
+ voe1 vout vout voe1 vss vout voe1 voe1 voe1 vout vout voe1 voe1 vss voe1 vout voe1
+ voe1 vout vout voe1 voe1 voe1 vout vss vout voe1 vss voe1 voe1 voe1 voe1 voe1 sky130_fd_pr__nfet_01v8_8JUMX6
Xsky130_fd_pr__pfet_01v8_YCMRKB_3 vin_p w_4660_n6791# vin_p voe1 voe1 vin_p vin_p
+ vin_p voe1 vin_p vin_p vin_p voe1 voe1 vin_p w_4660_n6791# vin_p vin_p vin_p vin_p
+ vin_p w_4660_n6791# voe1 vin_p w_4660_n6791# w_4660_n6791# voe1 vin_p voe1 w_4660_n6791#
+ vin_p w_4660_n6791# vin_p vin_p w_4660_n6791# w_4660_n6791# vin_p vin_p voe1 vin_p
+ voe1 vin_p vin_p voe1 w_4660_n6791# voe1 vin_p vin_p w_4660_n6791# w_4660_n6791#
+ w_4660_n6791# w_4660_n6791# voe1 vin_p voe1 vin_p vin_p w_4660_n6791# voe1 voe1
+ w_4660_n6791# voe1 w_4660_n6791# w_4660_n6791# vin_p w_4660_n6791# vin_p w_4660_n6791#
+ w_4660_n6791# vin_p vin_p vin_p voe1 voe1 w_4660_n6791# vin_p vin_p voe1 voe1 voe1
+ w_4660_n6791# voe1 vin_p vin_p vin_p voe1 vin_p vin_p vin_p voe1 voe1 vin_p w_4660_n6791#
+ vin_p voe1 vin_p vin_p w_4660_n6791# voe1 vin_p voe1 voe1 vin_p vin_p vin_p w_4660_n6791#
+ w_4660_n6791# vin_p vin_p vin_p voe1 vin_p w_4660_n6791# w_4660_n6791# vin_p vin_p
+ vin_p voe1 w_4660_n6791# vin_p w_4660_n6791# voe1 vin_p w_4660_n6791# vin_p vin_p
+ vin_p voe1 w_4660_n6791# vin_p voe1 voe1 vin_p w_4660_n6791# w_4660_n6791# vin_p
+ vin_p vin_p w_4660_n6791# w_4660_n6791# w_4660_n6791# vin_p vin_p w_4660_n6791#
+ w_4660_n6791# vin_p vin_p w_4660_n6791# voe1 vin_p voe1 w_4660_n6791# vin_p vin_p
+ w_4660_n6791# vin_p vin_p vin_p voe1 vin_p vin_p vin_p voe1 vin_p voe1 voe1 vin_p
+ vin_p w_4660_n6791# vin_p vin_p vin_p voe1 voe1 voe1 w_4660_n6791# vin_p w_4660_n6791#
+ vin_p w_4660_n6791# voe1 w_4660_n6791# vin_p voe1 w_4660_n6791# vin_p w_4660_n6791#
+ vin_p vin_p w_4660_n6791# vin_p vin_p vin_p vin_p vin_p w_4660_n6791# w_4660_n6791#
+ vin_p vin_p voe1 voe1 voe1 vin_p sky130_fd_pr__pfet_01v8_YCMRKB
.ends

.subckt TIA vin1 vin2 vout1 vout2 vdd vss
Xsky130_fd_pr__res_high_po_2p85_RN83L8_0 vout2 opamp_v1_1/vin_n vss sky130_fd_pr__res_high_po_2p85_RN83L8
Xsky130_fd_pr__nfet_01v8_UPGCN9_0 sky130_fd_pr__nfet_01v8_UPGCN9_0/G sky130_fd_pr__nfet_01v8_UPGCN9_0/G
+ vss vss sky130_fd_pr__nfet_01v8_UPGCN9
Xsky130_fd_pr__res_high_po_2p85_BNWAAK_0 vout1 opamp_v1_0/vin_n vss sky130_fd_pr__res_high_po_2p85_BNWAAK
Xsky130_fd_pr__nfet_01v8_LNQ4EK_0 iref vss sky130_fd_pr__nfet_01v8_UPGCN9_0/G vss
+ sky130_fd_pr__nfet_01v8_LNQ4EK
Xsky130_fd_pr__res_high_po_2p85_ZJW47V_0 vdd sky130_fd_pr__nfet_01v8_UPGCN9_0/G vss
+ sky130_fd_pr__res_high_po_2p85_ZJW47V
Xsky130_fd_pr__res_high_po_2p85_6SZAMJ_0 opamp_v1_0/vin_n vin2 vss sky130_fd_pr__res_high_po_2p85_6SZAMJ
Xsky130_fd_pr__res_high_po_2p85_6SZAMJ_1 vin1 opamp_v1_1/vin_n vss sky130_fd_pr__res_high_po_2p85_6SZAMJ
Xopamp_v1_0 vdd iref opamp_v1_0/vin_n vin1 vout1 vss vss opamp_v1
Xopamp_v1_1 vdd iref opamp_v1_1/vin_n vin2 vout2 vss vss opamp_v1
.ends


magic
tech sky130A
magscale 1 2
timestamp 1702074941
<< pwell >>
rect -285 -1679 285 1679
<< nmos >>
rect -89 -1531 -29 1469
rect 29 -1531 89 1469
<< ndiff >>
rect -147 1457 -89 1469
rect -147 -1519 -135 1457
rect -101 -1519 -89 1457
rect -147 -1531 -89 -1519
rect -29 1457 29 1469
rect -29 -1519 -17 1457
rect 17 -1519 29 1457
rect -29 -1531 29 -1519
rect 89 1457 147 1469
rect 89 -1519 101 1457
rect 135 -1519 147 1457
rect 89 -1531 147 -1519
<< ndiffc >>
rect -135 -1519 -101 1457
rect -17 -1519 17 1457
rect 101 -1519 135 1457
<< psubdiff >>
rect -249 1609 249 1643
rect -249 -1609 -215 1609
rect 215 -1609 249 1609
rect -249 -1643 -153 -1609
rect 153 -1643 249 -1609
<< psubdiffcont >>
rect -153 -1643 153 -1609
<< poly >>
rect -92 1541 -26 1557
rect -92 1507 -76 1541
rect -42 1507 -26 1541
rect -92 1491 -26 1507
rect 26 1541 92 1557
rect 26 1507 42 1541
rect 76 1507 92 1541
rect 26 1491 92 1507
rect -89 1469 -29 1491
rect 29 1469 89 1491
rect -89 -1557 -29 -1531
rect 29 -1557 89 -1531
<< polycont >>
rect -76 1507 -42 1541
rect 42 1507 76 1541
<< locali >>
rect -92 1507 -76 1541
rect -42 1507 -26 1541
rect 26 1507 42 1541
rect 76 1507 92 1541
rect -135 1457 -101 1473
rect -135 -1535 -101 -1519
rect -17 1457 17 1473
rect -17 -1535 17 -1519
rect 101 1457 135 1473
rect 101 -1535 135 -1519
rect -169 -1643 -153 -1609
rect 153 -1643 169 -1609
<< viali >>
rect -76 1507 -42 1541
rect 42 1507 76 1541
rect -135 -1519 -101 1457
rect -17 -1073 17 1011
rect 101 -1519 135 1457
<< metal1 >>
rect -88 1541 88 1547
rect -88 1507 -76 1541
rect -42 1507 42 1541
rect 76 1507 88 1541
rect -88 1501 88 1507
rect -141 1457 -95 1469
rect -141 -1519 -135 1457
rect -101 1405 -95 1457
rect 95 1457 141 1469
rect 95 1405 101 1457
rect -101 1366 101 1405
rect -101 -1519 -95 1366
rect -23 1011 23 1023
rect -23 -1073 -17 1011
rect 17 -1073 23 1011
rect -23 -1085 23 -1073
rect -141 -1531 -95 -1519
rect 95 -1519 101 1366
rect 135 -1519 141 1457
rect 95 -1531 141 -1519
<< labels >>
rlabel metal1 -101 1366 101 1405 1 D
port 1 n
rlabel metal1 -23 -1085 -17 1023 1 S
port 2 n
rlabel metal1 -42 1501 42 1547 1 G
port 3 n
rlabel locali -169 -1643 -153 -1609 1 B
port 4 n
<< properties >>
string FIXED_BBOX -232 -1626 232 1626
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 15 l 0.3 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 70 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

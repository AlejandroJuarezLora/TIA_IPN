magic
tech sky130A
magscale 1 2
timestamp 1702073221
<< error_p >>
rect -206 1372 -148 1378
rect -88 1372 -30 1378
rect 30 1372 88 1378
rect 148 1372 206 1378
rect -206 1338 -194 1372
rect -88 1338 -76 1372
rect 30 1338 42 1372
rect 148 1338 160 1372
rect -206 1332 -148 1338
rect -88 1332 -30 1338
rect 30 1332 88 1338
rect 148 1332 206 1338
rect -206 -1338 -148 -1332
rect -88 -1338 -30 -1332
rect 30 -1338 88 -1332
rect 148 -1338 206 -1332
rect -206 -1372 -194 -1338
rect -88 -1372 -76 -1338
rect 30 -1372 42 -1338
rect 148 -1372 160 -1338
rect -206 -1378 -148 -1372
rect -88 -1378 -30 -1372
rect 30 -1378 88 -1372
rect 148 -1378 206 -1372
<< pwell >>
rect -403 -1510 403 1510
<< nmos >>
rect -207 -1300 -147 1300
rect -89 -1300 -29 1300
rect 29 -1300 89 1300
rect 147 -1300 207 1300
<< ndiff >>
rect -265 1288 -207 1300
rect -265 -1288 -253 1288
rect -219 -1288 -207 1288
rect -265 -1300 -207 -1288
rect -147 1288 -89 1300
rect -147 -1288 -135 1288
rect -101 -1288 -89 1288
rect -147 -1300 -89 -1288
rect -29 1288 29 1300
rect -29 -1288 -17 1288
rect 17 -1288 29 1288
rect -29 -1300 29 -1288
rect 89 1288 147 1300
rect 89 -1288 101 1288
rect 135 -1288 147 1288
rect 89 -1300 147 -1288
rect 207 1288 265 1300
rect 207 -1288 219 1288
rect 253 -1288 265 1288
rect 207 -1300 265 -1288
<< ndiffc >>
rect -253 -1288 -219 1288
rect -135 -1288 -101 1288
rect -17 -1288 17 1288
rect 101 -1288 135 1288
rect 219 -1288 253 1288
<< psubdiff >>
rect -367 1440 -271 1474
rect 271 1440 367 1474
rect -367 1378 -333 1440
rect 333 1378 367 1440
rect -367 -1440 -333 -1378
rect 333 -1440 367 -1378
rect -367 -1474 -271 -1440
rect 271 -1474 367 -1440
<< psubdiffcont >>
rect -271 1440 271 1474
rect -367 -1378 -333 1378
rect 333 -1378 367 1378
rect -271 -1474 271 -1440
<< poly >>
rect -210 1372 -144 1388
rect -210 1338 -194 1372
rect -160 1338 -144 1372
rect -210 1322 -144 1338
rect -92 1372 -26 1388
rect -92 1338 -76 1372
rect -42 1338 -26 1372
rect -92 1322 -26 1338
rect 26 1372 92 1388
rect 26 1338 42 1372
rect 76 1338 92 1372
rect 26 1322 92 1338
rect 144 1372 210 1388
rect 144 1338 160 1372
rect 194 1338 210 1372
rect 144 1322 210 1338
rect -207 1300 -147 1322
rect -89 1300 -29 1322
rect 29 1300 89 1322
rect 147 1300 207 1322
rect -207 -1322 -147 -1300
rect -89 -1322 -29 -1300
rect 29 -1322 89 -1300
rect 147 -1322 207 -1300
rect -210 -1338 -144 -1322
rect -210 -1372 -194 -1338
rect -160 -1372 -144 -1338
rect -210 -1388 -144 -1372
rect -92 -1338 -26 -1322
rect -92 -1372 -76 -1338
rect -42 -1372 -26 -1338
rect -92 -1388 -26 -1372
rect 26 -1338 92 -1322
rect 26 -1372 42 -1338
rect 76 -1372 92 -1338
rect 26 -1388 92 -1372
rect 144 -1338 210 -1322
rect 144 -1372 160 -1338
rect 194 -1372 210 -1338
rect 144 -1388 210 -1372
<< polycont >>
rect -194 1338 -160 1372
rect -76 1338 -42 1372
rect 42 1338 76 1372
rect 160 1338 194 1372
rect -194 -1372 -160 -1338
rect -76 -1372 -42 -1338
rect 42 -1372 76 -1338
rect 160 -1372 194 -1338
<< locali >>
rect -367 1440 -271 1474
rect 271 1440 367 1474
rect -367 1378 -333 1440
rect 333 1378 367 1440
rect -210 1338 -194 1372
rect -160 1338 -144 1372
rect -92 1338 -76 1372
rect -42 1338 -26 1372
rect 26 1338 42 1372
rect 76 1338 92 1372
rect 144 1338 160 1372
rect 194 1338 210 1372
rect -253 1288 -219 1304
rect -253 -1304 -219 -1288
rect -135 1288 -101 1304
rect -135 -1304 -101 -1288
rect -17 1288 17 1304
rect -17 -1304 17 -1288
rect 101 1288 135 1304
rect 101 -1304 135 -1288
rect 219 1288 253 1304
rect 219 -1304 253 -1288
rect -210 -1372 -194 -1338
rect -160 -1372 -144 -1338
rect -92 -1372 -76 -1338
rect -42 -1372 -26 -1338
rect 26 -1372 42 -1338
rect 76 -1372 92 -1338
rect 144 -1372 160 -1338
rect 194 -1372 210 -1338
rect -367 -1440 -333 -1378
rect 333 -1440 367 -1378
rect -367 -1474 -271 -1440
rect 271 -1474 367 -1440
<< viali >>
rect -194 1338 -160 1372
rect -76 1338 -42 1372
rect 42 1338 76 1372
rect 160 1338 194 1372
rect -253 -1288 -219 1288
rect -135 -1288 -101 1288
rect -17 -1288 17 1288
rect 101 -1288 135 1288
rect 219 -1288 253 1288
rect -194 -1372 -160 -1338
rect -76 -1372 -42 -1338
rect 42 -1372 76 -1338
rect 160 -1372 194 -1338
<< metal1 >>
rect -206 1372 -148 1378
rect -206 1338 -194 1372
rect -160 1338 -148 1372
rect -206 1332 -148 1338
rect -88 1372 -30 1378
rect -88 1338 -76 1372
rect -42 1338 -30 1372
rect -88 1332 -30 1338
rect 30 1372 88 1378
rect 30 1338 42 1372
rect 76 1338 88 1372
rect 30 1332 88 1338
rect 148 1372 206 1378
rect 148 1338 160 1372
rect 194 1338 206 1372
rect 148 1332 206 1338
rect -259 1288 -213 1300
rect -259 -1288 -253 1288
rect -219 -1288 -213 1288
rect -259 -1300 -213 -1288
rect -141 1288 -95 1300
rect -141 -1288 -135 1288
rect -101 -1288 -95 1288
rect -141 -1300 -95 -1288
rect -23 1288 23 1300
rect -23 -1288 -17 1288
rect 17 -1288 23 1288
rect -23 -1300 23 -1288
rect 95 1288 141 1300
rect 95 -1288 101 1288
rect 135 -1288 141 1288
rect 95 -1300 141 -1288
rect 213 1288 259 1300
rect 213 -1288 219 1288
rect 253 -1288 259 1288
rect 213 -1300 259 -1288
rect -206 -1338 -148 -1332
rect -206 -1372 -194 -1338
rect -160 -1372 -148 -1338
rect -206 -1378 -148 -1372
rect -88 -1338 -30 -1332
rect -88 -1372 -76 -1338
rect -42 -1372 -30 -1338
rect -88 -1378 -30 -1372
rect 30 -1338 88 -1332
rect 30 -1372 42 -1338
rect 76 -1372 88 -1338
rect 30 -1378 88 -1372
rect 148 -1338 206 -1332
rect 148 -1372 160 -1338
rect 194 -1372 206 -1338
rect 148 -1378 206 -1372
<< properties >>
string FIXED_BBOX -350 -1457 350 1457
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 13 l 0.3 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

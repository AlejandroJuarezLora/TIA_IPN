magic
tech sky130A
magscale 1 2
timestamp 1702940054
<< locali >>
rect 1600 26431 1991 26465
rect 1600 25133 1634 26431
rect -818 25099 1634 25133
rect -818 17636 -784 25099
rect -818 17602 -570 17636
rect -814 17526 -780 17602
rect -814 17492 -606 17526
rect -812 15597 -778 17492
rect -1360 15563 -778 15597
rect -1360 12191 -1326 15563
rect -891 12191 -857 12276
rect -1360 12157 -857 12191
rect -891 11967 -857 12157
rect -891 11933 -464 11967
rect -337 11958 -302 12051
rect -794 11796 -760 11933
rect 443 11796 477 12058
rect -794 11762 477 11796
rect -794 11590 -760 11762
rect -794 11556 -630 11590
rect -794 941 -760 11556
rect -794 907 1667 941
rect 1633 275 1667 907
rect 1633 241 2017 275
<< metal1 >>
rect -610 26887 -604 27287
rect -204 26887 -198 27287
rect -604 24679 -204 26887
rect -472 17858 477 18031
rect 296 17405 477 17858
rect 296 17258 1045 17405
rect -488 17232 1045 17258
rect 1218 17232 1224 17405
rect -488 17085 469 17232
rect -2642 16018 -2394 16024
rect -2394 15770 -108 16018
rect -2642 15764 -2394 15770
rect -1011 15079 773 15123
rect -1011 15077 -782 15079
rect -720 15077 773 15079
rect -1011 14902 -965 15077
rect -824 14946 -782 14948
rect -824 14902 -730 14946
rect -778 14804 -732 14902
rect 727 14323 773 15077
rect -218 13504 -8 13689
rect 177 13504 190 13689
rect 1499 12461 1684 13109
rect 8989 12941 9629 13848
rect 860 12276 1684 12461
rect -1994 11218 -1988 11466
rect -1740 11218 -346 11466
rect -570 9882 562 10051
rect 376 9564 562 9882
rect 376 9395 1056 9564
rect 1225 9395 1231 9564
rect 376 9306 545 9395
rect -400 9137 545 9306
rect -586 -15 -186 1399
rect -592 -415 -586 -15
rect -186 -415 -180 -15
<< via1 >>
rect -604 26887 -204 27287
rect 1045 17232 1218 17405
rect -2642 15770 -2394 16018
rect -8 13504 177 13689
rect -1988 11218 -1740 11466
rect 1056 9395 1225 9564
rect -586 -415 -186 -15
<< metal2 >>
rect -604 27287 -204 27293
rect -608 26892 -604 27282
rect -204 26892 -200 27282
rect -604 26881 -204 26887
rect -4056 21291 1242 21539
rect -2648 15770 -2642 16018
rect -2394 15770 -2388 16018
rect -2642 5499 -2394 15770
rect -1988 11466 -1740 21291
rect 1045 17405 1218 17411
rect 1045 17226 1218 17232
rect -8 13689 190 14875
rect 177 13504 190 13689
rect -8 11903 190 13504
rect -1988 11212 -1740 11218
rect 1056 9564 1225 9570
rect 1056 9389 1225 9395
rect -3910 5251 1211 5499
rect -586 -15 -186 -9
rect -590 -410 -586 -20
rect -186 -410 -182 -20
rect -586 -421 -186 -415
<< via2 >>
rect -599 26892 -209 27282
rect -581 -410 -191 -20
<< metal3 >>
rect -604 27286 -204 27287
rect -609 26888 -603 27286
rect -205 26888 -199 27286
rect -604 26887 -204 26888
rect -585 -15 -187 -10
rect -586 -16 -186 -15
rect -586 -414 -585 -16
rect -187 -414 -186 -16
rect -586 -415 -186 -414
rect -585 -420 -187 -415
<< via3 >>
rect -603 27282 -205 27286
rect -603 26892 -599 27282
rect -599 26892 -209 27282
rect -209 26892 -205 27282
rect -603 26888 -205 26892
rect -585 -20 -187 -16
rect -585 -410 -581 -20
rect -581 -410 -191 -20
rect -191 -410 -187 -20
rect -585 -414 -187 -410
<< metal4 >>
rect -642 27286 24899 27287
rect -642 26888 -603 27286
rect -205 26888 24899 27286
rect -642 26887 24899 26888
rect 24499 20003 24899 26887
rect 24455 -15 24855 5488
rect -586 -16 -180 -15
rect -586 -414 -585 -16
rect -187 -32 -180 -16
rect 24454 -32 24855 -15
rect -187 -414 24855 -32
rect -586 -415 24855 -414
use opamp_v1  opamp_v1_0 ../mag
timestamp 1701460012
transform 1 0 -2072 0 -1 16762
box 2069 -10028 26971 3199
use opamp_v1  opamp_v1_1
timestamp 1701460012
transform 1 0 -2069 0 1 10028
box 2069 -10028 26971 3199
use sky130_fd_pr__nfet_01v8_LNQ4EK  sky130_fd_pr__nfet_01v8_LNQ4EK_0
timestamp 1702074941
transform 1 0 -319 0 1 13575
box -285 -1679 285 1679
use sky130_fd_pr__nfet_01v8_UPGCN9  sky130_fd_pr__nfet_01v8_UPGCN9_0
timestamp 1702073639
transform 1 0 -992 0 1 13601
box -403 -1479 403 1479
use sky130_fd_pr__res_high_po_2p85_6SZAMJ  sky130_fd_pr__res_high_po_2p85_6SZAMJ_0
timestamp 1701914711
transform 1 0 -402 0 1 16547
box -451 -1017 451 1017
use sky130_fd_pr__res_high_po_2p85_6SZAMJ  sky130_fd_pr__res_high_po_2p85_6SZAMJ_1
timestamp 1701914711
transform 1 0 -381 0 1 10612
box -451 -1017 451 1017
use sky130_fd_pr__res_high_po_2p85_BNWAAK  sky130_fd_pr__res_high_po_2p85_BNWAAK_0
timestamp 1701914995
transform -1 0 -403 0 1 21367
box -451 -3802 451 3802
use sky130_fd_pr__res_high_po_2p85_RN83L8  sky130_fd_pr__res_high_po_2p85_RN83L8_0
timestamp 1701914995
transform 1 0 -381 0 1 5233
box -451 -4360 451 4360
use sky130_fd_pr__res_high_po_2p85_ZJW47V  sky130_fd_pr__res_high_po_2p85_ZJW47V_0
timestamp 1702074941
transform 1 0 752 0 1 13342
box -451 -1352 451 1352
<< labels >>
rlabel metal2 -8 11903 190 14875 1 iref
rlabel metal4 24455 -415 24855 5488 0 vout2
port 3 nsew
flabel metal4 24499 20003 24899 27287 0 FreeSans 1600 0 0 0 vout1
port 2 nsew
flabel metal1 8989 12941 9629 13848 0 FreeSans 1600 0 0 0 vdd
port 4 nsew
flabel locali -794 907 1667 941 0 FreeSans 1600 0 0 0 vss
port 5 nsew
flabel metal2 s -4340 20896 -3476 21848 0 FreeSans 800 0 0 0 vin1
port 0 nsew
flabel metal2 s -4008 5032 -3566 5654 0 FreeSans 800 0 0 0 vin2
port 1 nsew
<< end >>

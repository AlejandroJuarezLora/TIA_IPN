** sch_path: /home/alex/Desktop/EDA/TIA_IPN/sch/TIA.sch
.subckt TIA vin1 vin2 vdd vss vout2 vout1
*.PININFO vin1:I vin2:I vdd:B vss:B vout2:O vout1:O
x1 vdd net1 net2 vin1 vout1 vss opamp_sky130
x2 vdd net1 net3 vin2 vout2 vss opamp_sky130
XR6 vout1 net2 vss sky130_fd_pr__res_high_po_2p85 L=31.85 mult=1 m=1
XR7 net3 vout2 vss sky130_fd_pr__res_high_po_2p85 L=37.354 mult=1 m=1
XR1 net2 vin2 vss sky130_fd_pr__res_high_po_2p85 L=4.348 mult=1 m=1
XR3 net3 vin1 vss sky130_fd_pr__res_high_po_2p85 L=4.348 mult=1 m=1
XM1 net1 net4 vss vss sky130_fd_pr__nfet_01v8 L=0.3 W=30 nf=1 m=1
XM2 net4 net4 vss vss sky130_fd_pr__nfet_01v8 L=0.3 W=54 nf=1 m=1
XR2 net4 vdd vss sky130_fd_pr__res_high_po_2p85 L=7.65 mult=1 m=1
.ends

* expanding   symbol:  /media/psf/EDA/TIA_IPN/sch/opamp_sky130.sym # of pins=6
** sym_path: /media/psf/EDA/TIA_IPN/sch/opamp_sky130.sym
** sch_path: /media/psf/EDA/TIA_IPN/sch/opamp_sky130.sch
.subckt opamp_sky130 vdd iref vin_n vin_p vout vss
*.PININFO vdd:B vss:B vin_n:I vin_p:I iref:I vout:O
XM1 vbn vin_n vp vp sky130_fd_pr__pfet_01v8 L=0.3 W=3 nf=1 m=200
XM2 voe1 vin_p vp vp sky130_fd_pr__pfet_01v8 L=0.3 W=3 nf=1 m=200
XM3 vbn vbn vss vss sky130_fd_pr__nfet_01v8 L=0.3 W=3 nf=1 m=30
XM4 voe1 vbn vss vss sky130_fd_pr__nfet_01v8 L=0.3 W=3 nf=1 m=30
XM5 vp iref vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=3 nf=1 m=30
XM7 vout iref vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=3 nf=1 m=150
XM8 iref iref vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=3 nf=1 m=15
XM9 net1 vdd voe1 vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.75 nf=1 m=6
XC1 net1 vout sky130_fd_pr__cap_mim_m3_1 W=17.55 L=15 m=6
XM6 vout voe1 vss vss sky130_fd_pr__nfet_01v8 L=0.45 W=4.5 nf=1 m=150
.ends

.end
